module fake_netlist_6_1198_n_5447 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_644, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_648, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_633, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_110, n_151, n_412, n_640, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_649, n_283, n_5447);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_648;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_633;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5447;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_677;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_3664;
wire n_1421;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_686;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_687;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_925;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_2767;
wire n_963;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_3299;
wire n_1419;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_858;
wire n_5182;
wire n_956;
wire n_663;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_664;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_662;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_3292;
wire n_1496;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_695;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_4027;
wire n_763;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_668;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_2356;
wire n_1511;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_666;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_659;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_3691;
wire n_1012;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_851;
wire n_682;
wire n_4991;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4866;
wire n_4889;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_688;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_936;
wire n_3821;
wire n_885;
wire n_2970;
wire n_2342;
wire n_2167;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_671;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_676;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_653;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5410;
wire n_2215;
wire n_1884;
wire n_665;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_681;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_5382;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_658;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_5374;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_689;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_692;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_690;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_696;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_3326;
wire n_2036;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_678;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_3252;
wire n_1634;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_656;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_684;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5442;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_651;
wire n_3407;
wire n_5313;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_2289;
wire n_1390;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_4754;
wire n_2993;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3501;
wire n_3475;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_2376;
wire n_1405;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5387;
wire n_654;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_1545;
wire n_4145;
wire n_4821;
wire n_3121;
wire n_4901;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_652;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_655;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_680;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_679;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_670;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_3910;
wire n_3812;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_821;
wire n_4372;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1014;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_4478;
wire n_1662;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_674;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_675;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_697;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_673;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_2316;
wire n_1771;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_657;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_2403;
wire n_1070;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1475;
wire n_716;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_4573;
wire n_5398;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_667;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5425;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_672;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_661;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_669;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_4243;
wire n_2205;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_5369;
wire n_975;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

BUFx3_ASAP7_75t_L g650 ( 
.A(n_560),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_610),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_446),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_412),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_303),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_31),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_314),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_421),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_452),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_450),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_20),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_544),
.Y(n_661)
);

BUFx8_ASAP7_75t_SL g662 ( 
.A(n_99),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_121),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_136),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_256),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_256),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_173),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_324),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_648),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_385),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_240),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_259),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_366),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_362),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_633),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_11),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_113),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_363),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_641),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_310),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_515),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_521),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_283),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_143),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_52),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_630),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_143),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_184),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_124),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_245),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_332),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_141),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_453),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_337),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_296),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_8),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_27),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_198),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_218),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_643),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_586),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_405),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_636),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_607),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_429),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_612),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_528),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_82),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_466),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_553),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_360),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_284),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_100),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_445),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_48),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_245),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_117),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_632),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_98),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_82),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_243),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_360),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_427),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_599),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_341),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_564),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_448),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_48),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_485),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_252),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_407),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_198),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_497),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_222),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_159),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_559),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_75),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_342),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_433),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_464),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_158),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_451),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_417),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_292),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_576),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_176),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_179),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_247),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_425),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_531),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_72),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_12),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_327),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_6),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_490),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_426),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_18),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_155),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_276),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_480),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_473),
.Y(n_761)
);

INVxp33_ASAP7_75t_R g762 ( 
.A(n_327),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_25),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_107),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_281),
.Y(n_765)
);

BUFx2_ASAP7_75t_SL g766 ( 
.A(n_21),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_126),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_308),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_443),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_121),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_40),
.Y(n_771)
);

BUFx5_ASAP7_75t_L g772 ( 
.A(n_260),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_46),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_217),
.Y(n_774)
);

BUFx10_ASAP7_75t_L g775 ( 
.A(n_101),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_296),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_210),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_625),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_371),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_66),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_104),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_30),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_20),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_73),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_547),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_179),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_628),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_223),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_112),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_441),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_167),
.Y(n_791)
);

CKINVDCx16_ASAP7_75t_R g792 ( 
.A(n_392),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_386),
.Y(n_793)
);

CKINVDCx14_ASAP7_75t_R g794 ( 
.A(n_116),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_605),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_259),
.Y(n_796)
);

CKINVDCx14_ASAP7_75t_R g797 ( 
.A(n_386),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_317),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_263),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_281),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_380),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_196),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_368),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_233),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_105),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_163),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_10),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_504),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_470),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_441),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_105),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_260),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_43),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_467),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_208),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_170),
.Y(n_816)
);

BUFx8_ASAP7_75t_SL g817 ( 
.A(n_9),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_215),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_159),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_417),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_230),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_66),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_563),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_313),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_123),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_347),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_378),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_596),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_543),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_399),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_475),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_156),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_68),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_394),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_646),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_585),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_295),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_156),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_93),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_626),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_21),
.Y(n_841)
);

BUFx10_ASAP7_75t_L g842 ( 
.A(n_570),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_318),
.Y(n_843)
);

CKINVDCx14_ASAP7_75t_R g844 ( 
.A(n_396),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_229),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_639),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_47),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_435),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_345),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_286),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_272),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_271),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_462),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_621),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_389),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_119),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_340),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_482),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_536),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_17),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_332),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_335),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_277),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_302),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_100),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_321),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_363),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_325),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_307),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_22),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_232),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_195),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_136),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_208),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_365),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_262),
.Y(n_876)
);

BUFx5_ASAP7_75t_L g877 ( 
.A(n_237),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_150),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_58),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_389),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_51),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_589),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_511),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_638),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_249),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_222),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_341),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_303),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_106),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_315),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_530),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_28),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_224),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_228),
.Y(n_894)
);

BUFx10_ASAP7_75t_L g895 ( 
.A(n_534),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_70),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_406),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_629),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_557),
.Y(n_899)
);

CKINVDCx14_ASAP7_75t_R g900 ( 
.A(n_225),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_345),
.Y(n_901)
);

BUFx10_ASAP7_75t_L g902 ( 
.A(n_141),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_187),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_365),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_336),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_359),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_217),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_135),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_170),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_115),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_435),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_181),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_421),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_371),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_405),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_387),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_197),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_5),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_193),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_177),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_297),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_284),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_74),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_119),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_457),
.Y(n_925)
);

BUFx8_ASAP7_75t_SL g926 ( 
.A(n_282),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_590),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_3),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_181),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_580),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_237),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_126),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_266),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_232),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_263),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_12),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_372),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_503),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_114),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_574),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_598),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_550),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_527),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_624),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_205),
.Y(n_945)
);

BUFx10_ASAP7_75t_L g946 ( 
.A(n_2),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_40),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_400),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_183),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_317),
.Y(n_950)
);

CKINVDCx6p67_ASAP7_75t_R g951 ( 
.A(n_392),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_418),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_380),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_68),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_50),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_305),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_301),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_9),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_406),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_1),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_571),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_106),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_115),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_197),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_353),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_368),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_533),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_430),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_300),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_191),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_62),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_216),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_350),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_622),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_58),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_523),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_465),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_619),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_310),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_253),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_396),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_608),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_276),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_416),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_125),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_93),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_597),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_282),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_385),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_461),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_420),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_236),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_577),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_410),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_50),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_70),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_460),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_304),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_313),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_193),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_38),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_39),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_316),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_471),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_63),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_418),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_551),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_315),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_278),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_176),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_173),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_397),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_647),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_344),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_267),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_357),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_125),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_274),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_535),
.Y(n_1019)
);

CKINVDCx16_ASAP7_75t_R g1020 ( 
.A(n_248),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_108),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_42),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_285),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_273),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_395),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_382),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_81),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_251),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_419),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_379),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_362),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_224),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_34),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_426),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_381),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_53),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_226),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_409),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_185),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_17),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_469),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_383),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_558),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_59),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_168),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_351),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_429),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_412),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_148),
.Y(n_1050)
);

BUFx10_ASAP7_75t_L g1051 ( 
.A(n_92),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_261),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_383),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_62),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_76),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_283),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_202),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_295),
.Y(n_1058)
);

CKINVDCx14_ASAP7_75t_R g1059 ( 
.A(n_507),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_288),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_488),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_230),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_153),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_407),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_110),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_378),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_147),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_290),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_272),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_422),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_67),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_101),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_513),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_45),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_253),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_273),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_400),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_279),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_235),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_7),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_134),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_336),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_449),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_81),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_518),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_487),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_107),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_593),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_644),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_520),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_279),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_250),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_424),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_339),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_145),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_280),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_448),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_36),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_347),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_246),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_573),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_415),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_302),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_172),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_582),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_255),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_328),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_203),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_142),
.Y(n_1109)
);

BUFx10_ASAP7_75t_L g1110 ( 
.A(n_123),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_63),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_330),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_205),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_356),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_387),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_157),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_157),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_269),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_234),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_377),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_352),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_481),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_10),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_290),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_286),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_565),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_903),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_772),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_772),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_772),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_772),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_903),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_772),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_772),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_986),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_772),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_986),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_772),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_877),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_877),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_877),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_877),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_1034),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_877),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_877),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_877),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_662),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_877),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_676),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_651),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_651),
.Y(n_1151)
);

INVxp33_ASAP7_75t_L g1152 ( 
.A(n_719),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_669),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_669),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_817),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_679),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_659),
.B(n_0),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_679),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_693),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_926),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_693),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1034),
.Y(n_1162)
);

INVxp67_ASAP7_75t_SL g1163 ( 
.A(n_1044),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_711),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_794),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_700),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_700),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_703),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_703),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_797),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_724),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_828),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_724),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_726),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_671),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_726),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_676),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_844),
.Y(n_1178)
);

CKINVDCx16_ASAP7_75t_R g1179 ( 
.A(n_764),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1060),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_742),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_900),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_792),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_742),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_810),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_787),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_787),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_650),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_702),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_722),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_859),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1020),
.Y(n_1192)
);

INVxp67_ASAP7_75t_SL g1193 ( 
.A(n_828),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_859),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_883),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1030),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1060),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_883),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_899),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_676),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_899),
.Y(n_1201)
);

INVxp33_ASAP7_75t_SL g1202 ( 
.A(n_721),
.Y(n_1202)
);

CKINVDCx14_ASAP7_75t_R g1203 ( 
.A(n_1059),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1091),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_927),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_927),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_977),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_977),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1057),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1091),
.Y(n_1210)
);

CKINVDCx16_ASAP7_75t_R g1211 ( 
.A(n_718),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_951),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_978),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_978),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_951),
.Y(n_1215)
);

XNOR2xp5_ASAP7_75t_L g1216 ( 
.A(n_753),
.B(n_0),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1050),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_990),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_990),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1013),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1013),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_822),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1042),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1042),
.Y(n_1224)
);

INVxp33_ASAP7_75t_SL g1225 ( 
.A(n_766),
.Y(n_1225)
);

INVxp33_ASAP7_75t_L g1226 ( 
.A(n_659),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_745),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1073),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1073),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_854),
.Y(n_1230)
);

INVxp33_ASAP7_75t_SL g1231 ( 
.A(n_766),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_676),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_745),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1085),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_652),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_653),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_654),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_676),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1085),
.Y(n_1239)
);

INVxp33_ASAP7_75t_SL g1240 ( 
.A(n_655),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1089),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_656),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_657),
.Y(n_1243)
);

CKINVDCx14_ASAP7_75t_R g1244 ( 
.A(n_854),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1089),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_824),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1090),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1090),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_832),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_870),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_722),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_811),
.Y(n_1252)
);

INVxp33_ASAP7_75t_L g1253 ( 
.A(n_663),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_811),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_996),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_650),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1004),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_661),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_996),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1022),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1022),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1065),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1065),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_695),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_745),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_878),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_695),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_695),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_695),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_695),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_735),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_735),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_1004),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_661),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_735),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_735),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_735),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1019),
.Y(n_1278)
);

CKINVDCx14_ASAP7_75t_R g1279 ( 
.A(n_1019),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_660),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_664),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_748),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_660),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_748),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_748),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_666),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_673),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_748),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_660),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_683),
.Y(n_1290)
);

INVxp33_ASAP7_75t_SL g1291 ( 
.A(n_684),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_748),
.Y(n_1292)
);

INVxp67_ASAP7_75t_SL g1293 ( 
.A(n_997),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_687),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_881),
.Y(n_1295)
);

CKINVDCx16_ASAP7_75t_R g1296 ( 
.A(n_667),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_780),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_780),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_780),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_997),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_688),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_780),
.Y(n_1302)
);

CKINVDCx14_ASAP7_75t_R g1303 ( 
.A(n_733),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_780),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_843),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_689),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_843),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_843),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_831),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_843),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_843),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_874),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_874),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_874),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_667),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_874),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_874),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_909),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_745),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_713),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_872),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_690),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_876),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_691),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_663),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_920),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_668),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_713),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_668),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_667),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_745),
.Y(n_1331)
);

INVxp33_ASAP7_75t_SL g1332 ( 
.A(n_692),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_670),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_733),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_670),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_672),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_672),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_674),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_674),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_744),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_677),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_677),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_678),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_678),
.Y(n_1344)
);

INVxp67_ASAP7_75t_SL g1345 ( 
.A(n_785),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_680),
.Y(n_1346)
);

INVxp33_ASAP7_75t_SL g1347 ( 
.A(n_694),
.Y(n_1347)
);

INVxp33_ASAP7_75t_L g1348 ( 
.A(n_680),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_696),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_729),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_697),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_697),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_698),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_698),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_714),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_714),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_728),
.Y(n_1357)
);

CKINVDCx14_ASAP7_75t_R g1358 ( 
.A(n_733),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_728),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_729),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_739),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_699),
.Y(n_1362)
);

CKINVDCx16_ASAP7_75t_R g1363 ( 
.A(n_685),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_739),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_741),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_741),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_685),
.Y(n_1367)
);

INVxp33_ASAP7_75t_SL g1368 ( 
.A(n_705),
.Y(n_1368)
);

INVxp33_ASAP7_75t_L g1369 ( 
.A(n_743),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_743),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_749),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_749),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_752),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_808),
.Y(n_1374)
);

INVxp33_ASAP7_75t_L g1375 ( 
.A(n_752),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_708),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1126),
.B(n_2),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_712),
.Y(n_1378)
);

INVxp33_ASAP7_75t_L g1379 ( 
.A(n_756),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_756),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_757),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_685),
.Y(n_1382)
);

INVxp33_ASAP7_75t_L g1383 ( 
.A(n_757),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_775),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_776),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_776),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_750),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_775),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_932),
.Y(n_1389)
);

INVxp33_ASAP7_75t_L g1390 ( 
.A(n_777),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_777),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_744),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_781),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_781),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_808),
.Y(n_1395)
);

INVxp33_ASAP7_75t_L g1396 ( 
.A(n_786),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_786),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_791),
.B(n_3),
.Y(n_1398)
);

INVxp33_ASAP7_75t_SL g1399 ( 
.A(n_715),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_814),
.B(n_4),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_791),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_799),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_799),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_800),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_800),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_804),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_804),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_806),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_814),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_806),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_759),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_818),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_759),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_818),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_826),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_716),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_943),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_826),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_827),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_827),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_833),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_833),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_768),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_834),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_834),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_823),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_847),
.Y(n_1427)
);

INVxp33_ASAP7_75t_SL g1428 ( 
.A(n_717),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_847),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_823),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_775),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_849),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_943),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_768),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_849),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_851),
.Y(n_1436)
);

CKINVDCx14_ASAP7_75t_R g1437 ( 
.A(n_750),
.Y(n_1437)
);

INVxp67_ASAP7_75t_SL g1438 ( 
.A(n_898),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_851),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_860),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_720),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_725),
.Y(n_1442)
);

INVxp67_ASAP7_75t_SL g1443 ( 
.A(n_898),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_860),
.Y(n_1444)
);

INVxp33_ASAP7_75t_L g1445 ( 
.A(n_862),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_862),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_871),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_964),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_871),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_886),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_886),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_727),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1122),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_888),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_790),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_790),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_779),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_888),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_892),
.Y(n_1459)
);

CKINVDCx16_ASAP7_75t_R g1460 ( 
.A(n_779),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_892),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1006),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_894),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1122),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_894),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1008),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_905),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_905),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_907),
.Y(n_1469)
);

INVxp33_ASAP7_75t_SL g1470 ( 
.A(n_730),
.Y(n_1470)
);

INVxp33_ASAP7_75t_L g1471 ( 
.A(n_907),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_731),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1126),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1024),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_910),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_910),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1029),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_916),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_916),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_918),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_918),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_919),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_665),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_943),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1033),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_919),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_779),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_921),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_921),
.Y(n_1489)
);

INVxp33_ASAP7_75t_SL g1490 ( 
.A(n_732),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_923),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_820),
.Y(n_1492)
);

INVxp33_ASAP7_75t_L g1493 ( 
.A(n_923),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_924),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_734),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_924),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_820),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_737),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_929),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_767),
.B(n_4),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_738),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_929),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_746),
.Y(n_1503)
);

INVxp33_ASAP7_75t_SL g1504 ( 
.A(n_747),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_852),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_958),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_958),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_960),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_943),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_943),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_960),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_852),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_911),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_962),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_962),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_751),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_754),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_975),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_975),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_911),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1055),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_758),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_913),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_981),
.Y(n_1524)
);

INVxp33_ASAP7_75t_L g1525 ( 
.A(n_981),
.Y(n_1525)
);

NOR2xp67_ASAP7_75t_L g1526 ( 
.A(n_767),
.B(n_5),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_984),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_984),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_998),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_998),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_999),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_750),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_999),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_913),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_789),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_763),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1000),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_914),
.Y(n_1538)
);

BUFx5_ASAP7_75t_L g1539 ( 
.A(n_842),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1000),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1005),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_765),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1177),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1312),
.Y(n_1544)
);

AND2x6_ASAP7_75t_L g1545 ( 
.A(n_1134),
.B(n_675),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1264),
.Y(n_1546)
);

INVx4_ASAP7_75t_L g1547 ( 
.A(n_1233),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1484),
.B(n_930),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1267),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1134),
.A2(n_1121),
.B(n_928),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1269),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1539),
.B(n_1293),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1227),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1244),
.B(n_830),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1227),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1539),
.B(n_658),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1270),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1203),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1203),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1175),
.Y(n_1560)
);

NOR2x1_ASAP7_75t_L g1561 ( 
.A(n_1334),
.B(n_1387),
.Y(n_1561)
);

BUFx12f_ASAP7_75t_L g1562 ( 
.A(n_1165),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1539),
.B(n_681),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1177),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1200),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1227),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1244),
.B(n_842),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1200),
.Y(n_1568)
);

AND2x6_ASAP7_75t_L g1569 ( 
.A(n_1233),
.B(n_914),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1331),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1377),
.A2(n_1011),
.B(n_1005),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1509),
.B(n_928),
.Y(n_1572)
);

BUFx12f_ASAP7_75t_L g1573 ( 
.A(n_1165),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1510),
.B(n_931),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1128),
.A2(n_1015),
.B(n_1011),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1232),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1331),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1539),
.B(n_682),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1331),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1129),
.A2(n_1131),
.B(n_1130),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1202),
.A2(n_701),
.B1(n_891),
.B2(n_778),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1188),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1183),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1331),
.Y(n_1584)
);

AND2x2_ASAP7_75t_SL g1585 ( 
.A(n_1157),
.B(n_1121),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1334),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1387),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1532),
.B(n_1007),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1417),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1417),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1149),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1232),
.Y(n_1592)
);

BUFx8_ASAP7_75t_SL g1593 ( 
.A(n_1147),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1271),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1233),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1238),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1233),
.Y(n_1597)
);

BUFx8_ASAP7_75t_L g1598 ( 
.A(n_1539),
.Y(n_1598)
);

OAI22x1_ASAP7_75t_SL g1599 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_1093),
.B2(n_1094),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1265),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1532),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1279),
.B(n_842),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1272),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1133),
.A2(n_945),
.B(n_931),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1211),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1265),
.Y(n_1606)
);

OAI22x1_ASAP7_75t_R g1607 ( 
.A1(n_1189),
.A2(n_1075),
.B1(n_762),
.B2(n_798),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1265),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1238),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1275),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1345),
.B(n_1350),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1265),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1276),
.Y(n_1613)
);

AND2x6_ASAP7_75t_L g1614 ( 
.A(n_1265),
.B(n_945),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1162),
.Y(n_1615)
);

BUFx12f_ASAP7_75t_L g1616 ( 
.A(n_1170),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1180),
.Y(n_1617)
);

AOI22x1_ASAP7_75t_SL g1618 ( 
.A1(n_1189),
.A2(n_1249),
.B1(n_1250),
.B2(n_1246),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1136),
.A2(n_1017),
.B(n_1015),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1149),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1279),
.A2(n_769),
.B1(n_771),
.B2(n_770),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1277),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1303),
.B(n_895),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1319),
.Y(n_1624)
);

CKINVDCx6p67_ASAP7_75t_R g1625 ( 
.A(n_1164),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1190),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1282),
.Y(n_1627)
);

OAI22x1_ASAP7_75t_SL g1628 ( 
.A1(n_1246),
.A2(n_1120),
.B1(n_1123),
.B2(n_1119),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1268),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1284),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1190),
.Y(n_1631)
);

BUFx12f_ASAP7_75t_L g1632 ( 
.A(n_1170),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1319),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1319),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1319),
.Y(n_1635)
);

OA21x2_ASAP7_75t_L g1636 ( 
.A1(n_1138),
.A2(n_1023),
.B(n_1017),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1286),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1539),
.B(n_686),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1319),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1188),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1285),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_R g1642 ( 
.A1(n_1202),
.A2(n_1124),
.B1(n_1049),
.B2(n_1071),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1288),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1360),
.B(n_950),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1268),
.Y(n_1645)
);

OAI22x1_ASAP7_75t_L g1646 ( 
.A1(n_1216),
.A2(n_830),
.B1(n_991),
.B2(n_906),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1305),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1433),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1433),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1294),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1305),
.Y(n_1651)
);

AOI22x1_ASAP7_75t_SL g1652 ( 
.A1(n_1249),
.A2(n_774),
.B1(n_782),
.B2(n_773),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1433),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1149),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1256),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1292),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1324),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1539),
.B(n_704),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1374),
.B(n_950),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1303),
.B(n_895),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1297),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1433),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1298),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1287),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1172),
.B(n_906),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1433),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1183),
.A2(n_1086),
.B1(n_783),
.B2(n_788),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1139),
.A2(n_966),
.B(n_957),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1358),
.B(n_895),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1395),
.B(n_1409),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1299),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1256),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1210),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1309),
.B(n_706),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1302),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1304),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1185),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1185),
.Y(n_1678)
);

BUFx12f_ASAP7_75t_L g1679 ( 
.A(n_1178),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1307),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1308),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1500),
.Y(n_1682)
);

INVx5_ASAP7_75t_L g1683 ( 
.A(n_1426),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1310),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1192),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1311),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1178),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1313),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1140),
.A2(n_966),
.B(n_957),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1258),
.Y(n_1690)
);

AND2x6_ASAP7_75t_L g1691 ( 
.A(n_1141),
.B(n_1010),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1258),
.B(n_707),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1314),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1316),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1274),
.Y(n_1695)
);

BUFx8_ASAP7_75t_SL g1696 ( 
.A(n_1147),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1317),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1274),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1534),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1150),
.Y(n_1700)
);

BUFx8_ASAP7_75t_SL g1701 ( 
.A(n_1155),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1300),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1193),
.A2(n_784),
.B1(n_796),
.B2(n_793),
.Y(n_1703)
);

CKINVDCx16_ASAP7_75t_R g1704 ( 
.A(n_1179),
.Y(n_1704)
);

BUFx8_ASAP7_75t_L g1705 ( 
.A(n_1442),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1426),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1358),
.B(n_789),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1142),
.Y(n_1708)
);

BUFx12f_ASAP7_75t_L g1709 ( 
.A(n_1182),
.Y(n_1709)
);

INVx6_ASAP7_75t_L g1710 ( 
.A(n_1300),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1526),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1151),
.Y(n_1712)
);

INVxp33_ASAP7_75t_SL g1713 ( 
.A(n_1182),
.Y(n_1713)
);

BUFx12f_ASAP7_75t_L g1714 ( 
.A(n_1155),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1153),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1144),
.A2(n_1026),
.B(n_1023),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1192),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1320),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1154),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1320),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1196),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1328),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1430),
.B(n_1010),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1328),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1156),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1158),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1340),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1145),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1340),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1392),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1159),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1161),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1392),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1146),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_1426),
.Y(n_1735)
);

BUFx12f_ASAP7_75t_L g1736 ( 
.A(n_1160),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1148),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1166),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1167),
.Y(n_1739)
);

AOI22x1_ASAP7_75t_SL g1740 ( 
.A1(n_1250),
.A2(n_801),
.B1(n_803),
.B2(n_802),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1437),
.B(n_789),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1411),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1411),
.Y(n_1743)
);

INVx4_ASAP7_75t_L g1744 ( 
.A(n_1413),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1413),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1196),
.Y(n_1746)
);

BUFx12f_ASAP7_75t_L g1747 ( 
.A(n_1160),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1423),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1209),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1423),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1434),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1437),
.B(n_902),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1212),
.B(n_902),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1163),
.B(n_709),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1434),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1168),
.Y(n_1756)
);

INVx5_ASAP7_75t_L g1757 ( 
.A(n_1455),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1438),
.B(n_1037),
.Y(n_1758)
);

BUFx8_ASAP7_75t_SL g1759 ( 
.A(n_1266),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1455),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1483),
.B(n_710),
.Y(n_1761)
);

INVx5_ASAP7_75t_L g1762 ( 
.A(n_1456),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1456),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1492),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1443),
.B(n_1037),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1542),
.Y(n_1766)
);

CKINVDCx8_ASAP7_75t_R g1767 ( 
.A(n_1283),
.Y(n_1767)
);

BUFx12f_ASAP7_75t_L g1768 ( 
.A(n_1209),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1453),
.B(n_1069),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1492),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1497),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1497),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1505),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1230),
.B(n_902),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1257),
.A2(n_805),
.B1(n_812),
.B2(n_807),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1464),
.B(n_1069),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1273),
.B(n_946),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1473),
.B(n_1092),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1169),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1278),
.B(n_736),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1171),
.B(n_1173),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1505),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1174),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1176),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1181),
.B(n_1092),
.Y(n_1785)
);

INVx5_ASAP7_75t_L g1786 ( 
.A(n_1512),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1184),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1222),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1186),
.A2(n_1102),
.B(n_1028),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1512),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1235),
.Y(n_1791)
);

BUFx6f_ASAP7_75t_L g1792 ( 
.A(n_1513),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1513),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1520),
.Y(n_1794)
);

AND2x6_ASAP7_75t_L g1795 ( 
.A(n_1400),
.B(n_1187),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1520),
.Y(n_1796)
);

BUFx8_ASAP7_75t_SL g1797 ( 
.A(n_1266),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1127),
.A2(n_813),
.B1(n_816),
.B2(n_815),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1235),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1236),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1236),
.Y(n_1801)
);

BUFx12f_ASAP7_75t_L g1802 ( 
.A(n_1212),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1191),
.B(n_1102),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1523),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1132),
.A2(n_819),
.B1(n_825),
.B2(n_821),
.Y(n_1805)
);

INVxp33_ASAP7_75t_L g1806 ( 
.A(n_1152),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1251),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1237),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1523),
.Y(n_1809)
);

BUFx8_ASAP7_75t_SL g1810 ( 
.A(n_1295),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1538),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1237),
.Y(n_1812)
);

BUFx12f_ASAP7_75t_L g1813 ( 
.A(n_1215),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1194),
.A2(n_1028),
.B(n_1026),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1538),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1325),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1327),
.Y(n_1817)
);

BUFx12f_ASAP7_75t_L g1818 ( 
.A(n_1215),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1329),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1252),
.B(n_740),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1333),
.Y(n_1821)
);

BUFx12f_ASAP7_75t_L g1822 ( 
.A(n_1242),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1195),
.B(n_991),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1335),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1198),
.B(n_1066),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1199),
.B(n_1066),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1336),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1242),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1243),
.B(n_946),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1243),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1201),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1205),
.A2(n_1039),
.B(n_1035),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1337),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1225),
.B(n_946),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1206),
.B(n_1113),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1281),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1281),
.B(n_955),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1290),
.B(n_955),
.Y(n_1838)
);

BUFx12f_ASAP7_75t_L g1839 ( 
.A(n_1290),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1254),
.B(n_755),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1338),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1339),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1341),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1255),
.B(n_760),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1207),
.Y(n_1845)
);

OA21x2_ASAP7_75t_L g1846 ( 
.A1(n_1208),
.A2(n_1039),
.B(n_1035),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1259),
.B(n_761),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1213),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1214),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1218),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1219),
.A2(n_1045),
.B(n_1040),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1220),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1221),
.Y(n_1853)
);

AOI22x1_ASAP7_75t_SL g1854 ( 
.A1(n_1295),
.A2(n_837),
.B1(n_839),
.B2(n_838),
.Y(n_1854)
);

XNOR2xp5_ASAP7_75t_L g1855 ( 
.A(n_1326),
.B(n_723),
.Y(n_1855)
);

AOI22x1_ASAP7_75t_SL g1856 ( 
.A1(n_1326),
.A2(n_841),
.B1(n_850),
.B2(n_845),
.Y(n_1856)
);

BUFx8_ASAP7_75t_L g1857 ( 
.A(n_1157),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1342),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1260),
.B(n_795),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1223),
.B(n_1113),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1240),
.A2(n_1332),
.B1(n_1347),
.B2(n_1291),
.Y(n_1861)
);

OAI22x1_ASAP7_75t_R g1862 ( 
.A1(n_1389),
.A2(n_868),
.B1(n_885),
.B2(n_857),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1301),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1240),
.A2(n_855),
.B1(n_861),
.B2(n_856),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1224),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1228),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1291),
.A2(n_1347),
.B1(n_1368),
.B2(n_1332),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1301),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1261),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1368),
.A2(n_863),
.B1(n_865),
.B2(n_864),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1229),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1343),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1234),
.B(n_1040),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1306),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1306),
.Y(n_1875)
);

OAI22x1_ASAP7_75t_SL g1876 ( 
.A1(n_1389),
.A2(n_1112),
.B1(n_1111),
.B2(n_866),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1239),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1241),
.B(n_1045),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1245),
.Y(n_1879)
);

AOI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1399),
.A2(n_867),
.B1(n_873),
.B2(n_869),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1262),
.B(n_809),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1344),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1322),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1346),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1351),
.Y(n_1885)
);

OAI21x1_ASAP7_75t_L g1886 ( 
.A1(n_1247),
.A2(n_1047),
.B(n_1046),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1248),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1322),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1349),
.B(n_955),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1318),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1352),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1321),
.Y(n_1892)
);

OAI21x1_ASAP7_75t_L g1893 ( 
.A1(n_1398),
.A2(n_1047),
.B(n_1046),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1892),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1710),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1893),
.B(n_1572),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1595),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1893),
.B(n_1353),
.Y(n_1898)
);

OAI21x1_ASAP7_75t_L g1899 ( 
.A1(n_1580),
.A2(n_1398),
.B(n_1263),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1572),
.B(n_1354),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1615),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1595),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1806),
.B(n_1349),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1700),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1553),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1712),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1715),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1806),
.B(n_1362),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1543),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1719),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1725),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1726),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1731),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1732),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1795),
.B(n_1362),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1615),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1738),
.Y(n_1917)
);

INVx3_ASAP7_75t_L g1918 ( 
.A(n_1595),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1739),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1756),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1553),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1572),
.B(n_1355),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1795),
.B(n_1376),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1552),
.B(n_1376),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1779),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1543),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1783),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1574),
.B(n_1356),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1784),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1787),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1795),
.B(n_1670),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1564),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1831),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1617),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1564),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1574),
.B(n_1357),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1574),
.B(n_1359),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1850),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1565),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1582),
.B(n_1323),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1565),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1814),
.B(n_1361),
.Y(n_1942)
);

INVx4_ASAP7_75t_L g1943 ( 
.A(n_1706),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1595),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1553),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1852),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1626),
.B(n_1378),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1795),
.B(n_1378),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1853),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1865),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1871),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1626),
.B(n_1226),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1795),
.B(n_1416),
.Y(n_1953)
);

BUFx8_ASAP7_75t_L g1954 ( 
.A(n_1562),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1670),
.B(n_1416),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1568),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1879),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1887),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1670),
.B(n_1441),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1548),
.B(n_1611),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1553),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1789),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1814),
.B(n_1364),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1631),
.B(n_1226),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1560),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1611),
.B(n_1441),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1789),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1617),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1548),
.B(n_1452),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1597),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1611),
.B(n_1452),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1597),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1568),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1708),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1759),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1832),
.B(n_1365),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1708),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1832),
.B(n_1886),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1728),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1555),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1728),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1548),
.B(n_1472),
.Y(n_1982)
);

AND2x6_ASAP7_75t_L g1983 ( 
.A(n_1623),
.B(n_1049),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1734),
.Y(n_1984)
);

INVx5_ASAP7_75t_L g1985 ( 
.A(n_1569),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1597),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1886),
.B(n_1366),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1734),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1576),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1737),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1737),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1834),
.A2(n_1428),
.B1(n_1470),
.B2(n_1399),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1807),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1788),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1555),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1807),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1576),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1869),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1869),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1710),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1597),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1631),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1592),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1592),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1591),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1585),
.B(n_1472),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1596),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1544),
.B(n_1699),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1673),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1600),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1596),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1567),
.B(n_1495),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1555),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1591),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1609),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1609),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1545),
.B(n_1495),
.Y(n_2017)
);

BUFx6f_ASAP7_75t_L g2018 ( 
.A(n_1555),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1545),
.B(n_1498),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1620),
.Y(n_2020)
);

CKINVDCx6p67_ASAP7_75t_R g2021 ( 
.A(n_1802),
.Y(n_2021)
);

XNOR2xp5_ASAP7_75t_L g2022 ( 
.A(n_1618),
.B(n_1448),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1620),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1873),
.B(n_1370),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1629),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1873),
.B(n_1371),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1629),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1645),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1645),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1781),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1781),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1873),
.B(n_1372),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1781),
.Y(n_2033)
);

NAND2xp33_ASAP7_75t_L g2034 ( 
.A(n_1545),
.B(n_1691),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1816),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1566),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1816),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1816),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1647),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1816),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1600),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1566),
.Y(n_2042)
);

AND2x6_ASAP7_75t_L g2043 ( 
.A(n_1660),
.B(n_1058),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1647),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1585),
.B(n_1253),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1545),
.B(n_1498),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1817),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1817),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_1890),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_1710),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1817),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_1682),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1545),
.B(n_1501),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1817),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1651),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_1878),
.B(n_1373),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1651),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1656),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1566),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1819),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1656),
.Y(n_2061)
);

INVx6_ASAP7_75t_L g2062 ( 
.A(n_1582),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1602),
.B(n_1501),
.Y(n_2063)
);

OAI21x1_ASAP7_75t_L g2064 ( 
.A1(n_1580),
.A2(n_1540),
.B(n_1537),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1682),
.B(n_1503),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1819),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1819),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1819),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1878),
.B(n_1380),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1566),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1820),
.B(n_1225),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1759),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1600),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1570),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1644),
.B(n_1503),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1821),
.Y(n_2076)
);

BUFx6f_ASAP7_75t_L g2077 ( 
.A(n_1570),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1821),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1821),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1663),
.Y(n_2080)
);

BUFx2_ASAP7_75t_L g2081 ( 
.A(n_1855),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1821),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1570),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1644),
.B(n_1253),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1663),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1676),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1570),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1676),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_1717),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1878),
.B(n_1381),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1680),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_SL g2092 ( 
.A1(n_1581),
.A2(n_1448),
.B1(n_1474),
.B2(n_1466),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_1600),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1824),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_1717),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1711),
.B(n_1516),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_L g2097 ( 
.A(n_1691),
.B(n_1516),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1680),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_SL g2099 ( 
.A1(n_1667),
.A2(n_1474),
.B1(n_1477),
.B2(n_1466),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1686),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1824),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1824),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1711),
.B(n_1517),
.Y(n_2103)
);

CKINVDCx11_ASAP7_75t_R g2104 ( 
.A(n_1767),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1686),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1824),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1654),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1644),
.B(n_1348),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1833),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1654),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1833),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1833),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1659),
.B(n_1348),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1833),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1577),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1672),
.B(n_1385),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1577),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1659),
.B(n_1369),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_1608),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_1583),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1842),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_1797),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1718),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1718),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1842),
.Y(n_2125)
);

AND2x2_ASAP7_75t_SL g2126 ( 
.A(n_1571),
.B(n_1058),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1842),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1842),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1718),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_L g2130 ( 
.A1(n_1550),
.A2(n_1668),
.B(n_1604),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1659),
.B(n_1369),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1843),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1843),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1718),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1692),
.B(n_1517),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1843),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1843),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1608),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1672),
.B(n_1522),
.Y(n_2139)
);

INVxp67_ASAP7_75t_L g2140 ( 
.A(n_1554),
.Y(n_2140)
);

XNOR2x2_ASAP7_75t_L g2141 ( 
.A(n_1646),
.B(n_1462),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1858),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1690),
.B(n_1522),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1858),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1858),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1858),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1872),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1872),
.Y(n_2148)
);

INVx4_ASAP7_75t_L g2149 ( 
.A(n_1706),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_1577),
.Y(n_2150)
);

AND3x2_ASAP7_75t_L g2151 ( 
.A(n_1753),
.B(n_1137),
.C(n_1135),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1872),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1872),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1720),
.Y(n_2154)
);

OAI22xp5_ASAP7_75t_SL g2155 ( 
.A1(n_1560),
.A2(n_1477),
.B1(n_1521),
.B2(n_1485),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_1690),
.B(n_1386),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1882),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1698),
.B(n_1536),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1882),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1720),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1882),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1882),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1720),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1640),
.Y(n_2164)
);

AND2x6_ASAP7_75t_L g2165 ( 
.A(n_1669),
.B(n_1064),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_SL g2166 ( 
.A(n_1830),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_1577),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1720),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1884),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1884),
.Y(n_2170)
);

AND2x6_ASAP7_75t_L g2171 ( 
.A(n_1707),
.B(n_1064),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1722),
.Y(n_2172)
);

BUFx6f_ASAP7_75t_L g2173 ( 
.A(n_1579),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1722),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1884),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_1554),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1722),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1884),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1723),
.B(n_1536),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_1698),
.B(n_1391),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1674),
.B(n_1556),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1885),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1885),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1722),
.Y(n_2184)
);

AND2x6_ASAP7_75t_L g2185 ( 
.A(n_1741),
.B(n_1067),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_1640),
.B(n_1393),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1885),
.Y(n_2187)
);

OAI21x1_ASAP7_75t_L g2188 ( 
.A1(n_1550),
.A2(n_1527),
.B(n_1524),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_1673),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1723),
.B(n_1375),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1885),
.Y(n_2191)
);

INVx5_ASAP7_75t_L g2192 ( 
.A(n_1569),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1827),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1723),
.B(n_1375),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1724),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1563),
.B(n_1428),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1724),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1827),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1841),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1841),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1845),
.Y(n_2201)
);

BUFx8_ASAP7_75t_L g2202 ( 
.A(n_1562),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_1840),
.B(n_1231),
.Y(n_2203)
);

NAND2xp33_ASAP7_75t_SL g2204 ( 
.A(n_1774),
.B(n_1152),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1579),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1724),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1724),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_1608),
.Y(n_2208)
);

INVx3_ASAP7_75t_L g2209 ( 
.A(n_1608),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1845),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1727),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1727),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1727),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1578),
.B(n_1470),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1777),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1638),
.B(n_1490),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1727),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1752),
.B(n_1296),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_1677),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1729),
.Y(n_2220)
);

INVx1_ASAP7_75t_SL g2221 ( 
.A(n_1797),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_1579),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1845),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1849),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1658),
.B(n_1490),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1849),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1849),
.Y(n_2227)
);

AND2x6_ASAP7_75t_L g2228 ( 
.A(n_1758),
.B(n_1067),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1729),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_1844),
.B(n_1231),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1655),
.B(n_1394),
.Y(n_2231)
);

AND2x4_ASAP7_75t_L g2232 ( 
.A(n_1655),
.B(n_1397),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1866),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1866),
.Y(n_2234)
);

BUFx8_ASAP7_75t_L g2235 ( 
.A(n_1573),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1729),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1729),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1706),
.B(n_1504),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1866),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_1590),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1546),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1549),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1551),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1735),
.B(n_1761),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1557),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1733),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1594),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1735),
.B(n_1504),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1735),
.B(n_829),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1603),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_1650),
.A2(n_1197),
.B1(n_1204),
.B2(n_1143),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1590),
.Y(n_2252)
);

INVx4_ASAP7_75t_L g2253 ( 
.A(n_1671),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1733),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1610),
.Y(n_2255)
);

OA21x2_ASAP7_75t_L g2256 ( 
.A1(n_1604),
.A2(n_1529),
.B(n_1528),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1590),
.Y(n_2257)
);

BUFx3_ASAP7_75t_L g2258 ( 
.A(n_1695),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_1590),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1733),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1613),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_1695),
.B(n_1401),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1758),
.B(n_1379),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1622),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1733),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1627),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1847),
.B(n_835),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_1864),
.A2(n_1217),
.B1(n_875),
.B2(n_880),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1758),
.B(n_1379),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1630),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1743),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_1612),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_1702),
.B(n_1402),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1765),
.B(n_1769),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1859),
.B(n_836),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_1881),
.B(n_1383),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1743),
.Y(n_2277)
);

INVx3_ASAP7_75t_L g2278 ( 
.A(n_1612),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1641),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1643),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1743),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1780),
.B(n_840),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1743),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1754),
.B(n_1586),
.Y(n_2284)
);

OR2x6_ASAP7_75t_L g2285 ( 
.A(n_1960),
.B(n_1822),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2188),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_2104),
.Y(n_2287)
);

INVx1_ASAP7_75t_SL g2288 ( 
.A(n_1994),
.Y(n_2288)
);

INVxp33_ASAP7_75t_L g2289 ( 
.A(n_1901),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1909),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2140),
.B(n_1830),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_1952),
.B(n_1586),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_1901),
.Y(n_2293)
);

NOR2x1p5_ASAP7_75t_L g2294 ( 
.A(n_2021),
.B(n_1625),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2188),
.Y(n_2295)
);

CKINVDCx11_ASAP7_75t_R g2296 ( 
.A(n_2104),
.Y(n_2296)
);

CKINVDCx20_ASAP7_75t_R g2297 ( 
.A(n_1965),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1904),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_L g2299 ( 
.A(n_1931),
.B(n_1569),
.Y(n_2299)
);

AND3x2_ASAP7_75t_L g2300 ( 
.A(n_2049),
.B(n_1685),
.C(n_1678),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1906),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1909),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_1896),
.Y(n_2303)
);

INVx3_ASAP7_75t_L g2304 ( 
.A(n_1896),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1926),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_2062),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_1896),
.B(n_2181),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_SL g2308 ( 
.A(n_1916),
.B(n_1767),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1926),
.Y(n_2309)
);

INVx3_ASAP7_75t_L g2310 ( 
.A(n_2256),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1898),
.B(n_1861),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_2256),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_2256),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1942),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2276),
.B(n_1571),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1907),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_1960),
.A2(n_1867),
.B1(n_1766),
.B2(n_1664),
.Y(n_2317)
);

INVx3_ASAP7_75t_L g2318 ( 
.A(n_1898),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1910),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_1952),
.B(n_1587),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1932),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1932),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2176),
.B(n_1791),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1935),
.Y(n_2324)
);

NAND2xp33_ASAP7_75t_L g2325 ( 
.A(n_2228),
.B(n_1569),
.Y(n_2325)
);

INVx5_ASAP7_75t_L g2326 ( 
.A(n_1978),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1911),
.Y(n_2327)
);

INVx2_ASAP7_75t_SL g2328 ( 
.A(n_2126),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_1935),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1939),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1939),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_R g2332 ( 
.A(n_2072),
.B(n_1558),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1941),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1912),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_1898),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1913),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1915),
.B(n_1598),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1914),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2276),
.B(n_1571),
.Y(n_2339)
);

HB1xp67_ASAP7_75t_L g2340 ( 
.A(n_1916),
.Y(n_2340)
);

BUFx10_ASAP7_75t_L g2341 ( 
.A(n_2166),
.Y(n_2341)
);

AO22x2_ASAP7_75t_L g2342 ( 
.A1(n_2006),
.A2(n_1740),
.B1(n_1854),
.B2(n_1652),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1917),
.Y(n_2343)
);

NAND2xp33_ASAP7_75t_L g2344 ( 
.A(n_2228),
.B(n_1569),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1941),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2126),
.A2(n_1665),
.B1(n_1619),
.B2(n_1636),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_1964),
.B(n_1587),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2084),
.Y(n_2348)
);

HB1xp67_ASAP7_75t_L g2349 ( 
.A(n_1934),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1919),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1920),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1956),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1925),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1956),
.Y(n_2354)
);

OR2x6_ASAP7_75t_L g2355 ( 
.A(n_2017),
.B(n_1822),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2071),
.B(n_1791),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2274),
.B(n_1601),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1927),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1929),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_1923),
.B(n_1598),
.Y(n_2360)
);

AOI22xp5_ASAP7_75t_L g2361 ( 
.A1(n_2071),
.A2(n_1863),
.B1(n_1874),
.B2(n_1808),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2203),
.B(n_1808),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_2130),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1930),
.Y(n_2364)
);

OR2x6_ASAP7_75t_L g2365 ( 
.A(n_2019),
.B(n_1839),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_L g2366 ( 
.A1(n_1942),
.A2(n_1665),
.B1(n_1619),
.B2(n_1636),
.Y(n_2366)
);

BUFx10_ASAP7_75t_L g2367 ( 
.A(n_2166),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1973),
.Y(n_2368)
);

INVx4_ASAP7_75t_L g2369 ( 
.A(n_1943),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1933),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1938),
.Y(n_2371)
);

NAND3xp33_ASAP7_75t_L g2372 ( 
.A(n_2006),
.B(n_1880),
.C(n_1870),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2274),
.B(n_1601),
.Y(n_2373)
);

OR2x2_ASAP7_75t_L g2374 ( 
.A(n_1934),
.B(n_1637),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2072),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_R g2376 ( 
.A(n_1965),
.B(n_1558),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1973),
.Y(n_2377)
);

INVx3_ASAP7_75t_L g2378 ( 
.A(n_2130),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2021),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1989),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1946),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1949),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_2166),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_1942),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1989),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1950),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_1948),
.B(n_1598),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_1963),
.Y(n_2388)
);

INVxp67_ASAP7_75t_SL g2389 ( 
.A(n_2272),
.Y(n_2389)
);

BUFx4f_ASAP7_75t_L g2390 ( 
.A(n_1983),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1997),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1951),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1957),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_1997),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2003),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1958),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_1953),
.B(n_1863),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2003),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_1964),
.B(n_2084),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2004),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_1963),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_1963),
.Y(n_2402)
);

NAND2xp33_ASAP7_75t_L g2403 ( 
.A(n_2228),
.B(n_1614),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2004),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2203),
.B(n_1889),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_1976),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2007),
.Y(n_2407)
);

CKINVDCx6p67_ASAP7_75t_R g2408 ( 
.A(n_1975),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2007),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2011),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_2230),
.B(n_1874),
.Y(n_2411)
);

NOR3xp33_ASAP7_75t_L g2412 ( 
.A(n_1969),
.B(n_1704),
.C(n_2155),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2230),
.B(n_1829),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2011),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2244),
.B(n_2284),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2015),
.Y(n_2416)
);

AOI22xp33_ASAP7_75t_L g2417 ( 
.A1(n_1976),
.A2(n_1619),
.B1(n_1636),
.B2(n_1575),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_R g2418 ( 
.A(n_2204),
.B(n_1559),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_1924),
.B(n_1713),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_1978),
.B(n_1976),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_1987),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_1987),
.Y(n_2422)
);

AOI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2045),
.A2(n_1924),
.B1(n_2043),
.B2(n_1983),
.Y(n_2423)
);

INVx5_ASAP7_75t_L g2424 ( 
.A(n_1978),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1894),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2015),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_1954),
.Y(n_2427)
);

OAI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_1982),
.A2(n_1637),
.B1(n_1657),
.B2(n_1799),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2030),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2016),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_L g2431 ( 
.A(n_1955),
.B(n_1713),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2031),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2016),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_1987),
.B(n_1588),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2108),
.B(n_1702),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2033),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2025),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2193),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2025),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2198),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_2045),
.B(n_1801),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2199),
.Y(n_2442)
);

INVxp33_ASAP7_75t_SL g2443 ( 
.A(n_1968),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_SL g2444 ( 
.A(n_2164),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2196),
.B(n_1828),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_1959),
.B(n_1799),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2200),
.Y(n_2447)
);

AO22x2_ASAP7_75t_L g2448 ( 
.A1(n_1969),
.A2(n_1856),
.B1(n_1642),
.B2(n_1621),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2064),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2064),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_1966),
.B(n_1800),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2108),
.B(n_2113),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2186),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2113),
.B(n_1837),
.Y(n_2454)
);

INVx3_ASAP7_75t_L g2455 ( 
.A(n_1962),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_1967),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2027),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2214),
.B(n_1868),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2027),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2186),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2028),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2118),
.B(n_1838),
.Y(n_2462)
);

NAND3xp33_ASAP7_75t_SL g2463 ( 
.A(n_1992),
.B(n_1521),
.C(n_1485),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2186),
.Y(n_2464)
);

AND3x2_ASAP7_75t_L g2465 ( 
.A(n_1968),
.B(n_1746),
.C(n_1721),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2028),
.Y(n_2466)
);

OAI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_2216),
.A2(n_2225),
.B1(n_1971),
.B2(n_2053),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2029),
.Y(n_2468)
);

AND2x2_ASAP7_75t_SL g2469 ( 
.A(n_2034),
.B(n_1575),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_1899),
.Y(n_2470)
);

NAND2xp33_ASAP7_75t_R g2471 ( 
.A(n_2089),
.B(n_1605),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2231),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2062),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2118),
.B(n_1800),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_2000),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2029),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2046),
.B(n_1875),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2039),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2039),
.Y(n_2479)
);

BUFx3_ASAP7_75t_L g2480 ( 
.A(n_2062),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2044),
.Y(n_2481)
);

OR2x6_ASAP7_75t_L g2482 ( 
.A(n_2131),
.B(n_1839),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2231),
.Y(n_2483)
);

INVx2_ASAP7_75t_SL g2484 ( 
.A(n_2131),
.Y(n_2484)
);

AND2x6_ASAP7_75t_L g2485 ( 
.A(n_2190),
.B(n_1561),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2044),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_1954),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2190),
.B(n_1883),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2055),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2231),
.Y(n_2490)
);

INVx4_ASAP7_75t_SL g2491 ( 
.A(n_2228),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2232),
.Y(n_2492)
);

INVx4_ASAP7_75t_L g2493 ( 
.A(n_1943),
.Y(n_2493)
);

NOR2x1p5_ASAP7_75t_L g2494 ( 
.A(n_2218),
.B(n_1625),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2000),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2232),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2050),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2055),
.Y(n_2498)
);

INVx1_ASAP7_75t_SL g2499 ( 
.A(n_1903),
.Y(n_2499)
);

INVx8_ASAP7_75t_L g2500 ( 
.A(n_2228),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2194),
.B(n_1575),
.Y(n_2501)
);

CKINVDCx20_ASAP7_75t_R g2502 ( 
.A(n_2092),
.Y(n_2502)
);

NAND3xp33_ASAP7_75t_L g2503 ( 
.A(n_2215),
.B(n_1857),
.C(n_1775),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_1954),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2232),
.Y(n_2505)
);

INVx2_ASAP7_75t_SL g2506 ( 
.A(n_2194),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2263),
.B(n_1716),
.Y(n_2507)
);

BUFx8_ASAP7_75t_SL g2508 ( 
.A(n_2081),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2057),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2262),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2057),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2058),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_SL g2513 ( 
.A(n_2164),
.Y(n_2513)
);

INVx4_ASAP7_75t_L g2514 ( 
.A(n_1943),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2263),
.B(n_1716),
.Y(n_2515)
);

AND2x6_ASAP7_75t_L g2516 ( 
.A(n_2269),
.B(n_1071),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2058),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2262),
.Y(n_2518)
);

XOR2x2_ASAP7_75t_L g2519 ( 
.A(n_2099),
.B(n_1607),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2269),
.B(n_1812),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2262),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_2050),
.Y(n_2522)
);

OAI22xp33_ASAP7_75t_SL g2523 ( 
.A1(n_2075),
.A2(n_1363),
.B1(n_1367),
.B2(n_1315),
.Y(n_2523)
);

INVx5_ASAP7_75t_L g2524 ( 
.A(n_1985),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_1899),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2061),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2273),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2061),
.Y(n_2528)
);

INVxp67_ASAP7_75t_L g2529 ( 
.A(n_1908),
.Y(n_2529)
);

BUFx10_ASAP7_75t_L g2530 ( 
.A(n_2151),
.Y(n_2530)
);

AO21x2_ASAP7_75t_L g2531 ( 
.A1(n_2034),
.A2(n_1689),
.B(n_1668),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2273),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2080),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2080),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2273),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2201),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2085),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_1905),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2085),
.Y(n_2539)
);

OR2x2_ASAP7_75t_L g2540 ( 
.A(n_2009),
.B(n_1657),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2210),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2223),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_L g2543 ( 
.A(n_2052),
.B(n_1812),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2086),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2086),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2224),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2088),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2088),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2238),
.B(n_1888),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_2248),
.B(n_1836),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2226),
.Y(n_2551)
);

NAND2xp33_ASAP7_75t_L g2552 ( 
.A(n_1983),
.B(n_1614),
.Y(n_2552)
);

NAND3xp33_ASAP7_75t_L g2553 ( 
.A(n_2215),
.B(n_1857),
.C(n_1703),
.Y(n_2553)
);

BUFx10_ASAP7_75t_L g2554 ( 
.A(n_2171),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2258),
.Y(n_2555)
);

BUFx4f_ASAP7_75t_L g2556 ( 
.A(n_1983),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2149),
.B(n_1836),
.Y(n_2557)
);

INVxp33_ASAP7_75t_L g2558 ( 
.A(n_2009),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2227),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_2149),
.B(n_1947),
.Y(n_2560)
);

INVx3_ASAP7_75t_L g2561 ( 
.A(n_2107),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2233),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2091),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2202),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2258),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2234),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2002),
.B(n_1749),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2239),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_2202),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2091),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_1900),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_1905),
.Y(n_2572)
);

BUFx3_ASAP7_75t_L g2573 ( 
.A(n_1895),
.Y(n_2573)
);

AOI22xp33_ASAP7_75t_L g2574 ( 
.A1(n_1900),
.A2(n_1716),
.B1(n_1691),
.B2(n_1765),
.Y(n_2574)
);

OR2x6_ASAP7_75t_L g2575 ( 
.A(n_1895),
.B(n_1768),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2149),
.B(n_1857),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2098),
.Y(n_2577)
);

BUFx10_ASAP7_75t_L g2578 ( 
.A(n_2171),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_1900),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_1922),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_1922),
.A2(n_1691),
.B1(n_1769),
.B2(n_1765),
.Y(n_2581)
);

OAI22xp33_ASAP7_75t_L g2582 ( 
.A1(n_2135),
.A2(n_1687),
.B1(n_1384),
.B2(n_1431),
.Y(n_2582)
);

INVx4_ASAP7_75t_L g2583 ( 
.A(n_1985),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_1922),
.A2(n_1691),
.B1(n_1776),
.B2(n_1769),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2098),
.Y(n_2585)
);

INVx4_ASAP7_75t_L g2586 ( 
.A(n_1985),
.Y(n_2586)
);

NAND2xp33_ASAP7_75t_L g2587 ( 
.A(n_1983),
.B(n_1614),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2139),
.B(n_1687),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2100),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2282),
.B(n_1776),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_1928),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2043),
.B(n_1776),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2100),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2143),
.B(n_2158),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2105),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_1928),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_1928),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2105),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2189),
.B(n_2002),
.Y(n_2599)
);

BUFx4f_ASAP7_75t_L g2600 ( 
.A(n_2043),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2107),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2110),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2043),
.B(n_1778),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_1936),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2110),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2065),
.B(n_1388),
.Y(n_2606)
);

INVx3_ASAP7_75t_L g2607 ( 
.A(n_2123),
.Y(n_2607)
);

AOI21x1_ASAP7_75t_L g2608 ( 
.A1(n_2249),
.A2(n_1689),
.B(n_1675),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2043),
.B(n_1778),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_1974),
.Y(n_2610)
);

OR2x6_ASAP7_75t_L g2611 ( 
.A(n_1936),
.B(n_1768),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_1977),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2075),
.B(n_1605),
.Y(n_2613)
);

INVxp33_ASAP7_75t_L g2614 ( 
.A(n_2189),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2165),
.B(n_1778),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_1979),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_1936),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_1937),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_1981),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_1937),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_1937),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_1905),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_1984),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_1988),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_1985),
.B(n_1559),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2241),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_1990),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_2202),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2242),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_1991),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_1993),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2192),
.B(n_1683),
.Y(n_2632)
);

BUFx6f_ASAP7_75t_L g2633 ( 
.A(n_1905),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2243),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2245),
.Y(n_2635)
);

AND3x1_ASAP7_75t_L g2636 ( 
.A(n_2251),
.B(n_1076),
.C(n_1074),
.Y(n_2636)
);

BUFx8_ASAP7_75t_SL g2637 ( 
.A(n_2120),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2247),
.Y(n_2638)
);

INVxp33_ASAP7_75t_L g2639 ( 
.A(n_2096),
.Y(n_2639)
);

INVx3_ASAP7_75t_L g2640 ( 
.A(n_2123),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_2116),
.Y(n_2641)
);

BUFx2_ASAP7_75t_L g2642 ( 
.A(n_2095),
.Y(n_2642)
);

BUFx6f_ASAP7_75t_L g2643 ( 
.A(n_1921),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2124),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2103),
.B(n_1460),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2250),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2165),
.B(n_1846),
.Y(n_2647)
);

INVx3_ASAP7_75t_L g2648 ( 
.A(n_2124),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2005),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2255),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2261),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2014),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2020),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2023),
.Y(n_2654)
);

OAI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_2179),
.A2(n_2280),
.B1(n_2266),
.B2(n_2270),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2129),
.Y(n_2656)
);

BUFx10_ASAP7_75t_L g2657 ( 
.A(n_2171),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2024),
.A2(n_1851),
.B1(n_1846),
.B2(n_1825),
.Y(n_2658)
);

AND2x4_ASAP7_75t_L g2659 ( 
.A(n_2024),
.B(n_1823),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2264),
.Y(n_2660)
);

INVx6_ASAP7_75t_L g2661 ( 
.A(n_2116),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2279),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_1996),
.Y(n_2663)
);

NAND2xp33_ASAP7_75t_L g2664 ( 
.A(n_2165),
.B(n_1614),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_1998),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2179),
.B(n_1573),
.Y(n_2666)
);

NAND2xp33_ASAP7_75t_SL g2667 ( 
.A(n_2012),
.B(n_1074),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_1999),
.Y(n_2668)
);

NAND3xp33_ASAP7_75t_L g2669 ( 
.A(n_2204),
.B(n_1805),
.C(n_1798),
.Y(n_2669)
);

INVx1_ASAP7_75t_SL g2670 ( 
.A(n_2219),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2165),
.A2(n_853),
.B1(n_858),
.B2(n_846),
.Y(n_2671)
);

INVx2_ASAP7_75t_SL g2672 ( 
.A(n_2116),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2024),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2268),
.B(n_1280),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2165),
.B(n_1846),
.Y(n_2675)
);

CKINVDCx5p33_ASAP7_75t_R g2676 ( 
.A(n_2235),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2129),
.Y(n_2677)
);

BUFx3_ASAP7_75t_L g2678 ( 
.A(n_2026),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2134),
.Y(n_2679)
);

OR2x2_ASAP7_75t_L g2680 ( 
.A(n_2063),
.B(n_1289),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_2008),
.B(n_1616),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2026),
.Y(n_2682)
);

INVx1_ASAP7_75t_SL g2683 ( 
.A(n_2122),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2026),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2134),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2032),
.Y(n_2686)
);

BUFx10_ASAP7_75t_L g2687 ( 
.A(n_2171),
.Y(n_2687)
);

OAI21xp33_ASAP7_75t_SL g2688 ( 
.A1(n_2008),
.A2(n_1077),
.B(n_1076),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2032),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2495),
.B(n_2032),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2512),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2512),
.Y(n_2692)
);

AND2x2_ASAP7_75t_SL g2693 ( 
.A(n_2356),
.B(n_2097),
.Y(n_2693)
);

INVx5_ASAP7_75t_L g2694 ( 
.A(n_2611),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2495),
.B(n_2056),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2415),
.B(n_2171),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2517),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2304),
.Y(n_2698)
);

BUFx2_ASAP7_75t_L g2699 ( 
.A(n_2642),
.Y(n_2699)
);

AND2x4_ASAP7_75t_L g2700 ( 
.A(n_2497),
.B(n_2056),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_2599),
.Y(n_2701)
);

INVx2_ASAP7_75t_SL g2702 ( 
.A(n_2288),
.Y(n_2702)
);

AND2x6_ASAP7_75t_L g2703 ( 
.A(n_2423),
.B(n_2304),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2517),
.Y(n_2704)
);

INVx1_ASAP7_75t_SL g2705 ( 
.A(n_2670),
.Y(n_2705)
);

BUFx6f_ASAP7_75t_L g2706 ( 
.A(n_2303),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2526),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2526),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2474),
.B(n_2156),
.Y(n_2709)
);

INVx4_ASAP7_75t_L g2710 ( 
.A(n_2303),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_2297),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2528),
.Y(n_2712)
);

INVxp67_ASAP7_75t_L g2713 ( 
.A(n_2567),
.Y(n_2713)
);

INVx3_ASAP7_75t_L g2714 ( 
.A(n_2303),
.Y(n_2714)
);

OR2x6_ASAP7_75t_L g2715 ( 
.A(n_2611),
.B(n_1714),
.Y(n_2715)
);

INVx4_ASAP7_75t_L g2716 ( 
.A(n_2303),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_L g2717 ( 
.A(n_2362),
.B(n_1616),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2528),
.Y(n_2718)
);

NAND3xp33_ASAP7_75t_L g2719 ( 
.A(n_2411),
.B(n_1705),
.C(n_2097),
.Y(n_2719)
);

INVx8_ASAP7_75t_L g2720 ( 
.A(n_2611),
.Y(n_2720)
);

BUFx4f_ASAP7_75t_L g2721 ( 
.A(n_2611),
.Y(n_2721)
);

INVx1_ASAP7_75t_SL g2722 ( 
.A(n_2443),
.Y(n_2722)
);

AND2x4_ASAP7_75t_SL g2723 ( 
.A(n_2341),
.B(n_2156),
.Y(n_2723)
);

OR2x2_ASAP7_75t_L g2724 ( 
.A(n_2374),
.B(n_2221),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2533),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2533),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2314),
.Y(n_2727)
);

INVx3_ASAP7_75t_L g2728 ( 
.A(n_2304),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_L g2729 ( 
.A1(n_2328),
.A2(n_2185),
.B1(n_2069),
.B2(n_2090),
.Y(n_2729)
);

NAND3x1_ASAP7_75t_L g2730 ( 
.A(n_2412),
.B(n_1599),
.C(n_2022),
.Y(n_2730)
);

AND2x4_ASAP7_75t_L g2731 ( 
.A(n_2497),
.B(n_2056),
.Y(n_2731)
);

INVx1_ASAP7_75t_SL g2732 ( 
.A(n_2443),
.Y(n_2732)
);

NOR2x1p5_ASAP7_75t_L g2733 ( 
.A(n_2379),
.B(n_1802),
.Y(n_2733)
);

NOR2xp33_ASAP7_75t_L g2734 ( 
.A(n_2405),
.B(n_1632),
.Y(n_2734)
);

CKINVDCx20_ASAP7_75t_R g2735 ( 
.A(n_2297),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2429),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2314),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2432),
.Y(n_2738)
);

HB1xp67_ASAP7_75t_L g2739 ( 
.A(n_2293),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2522),
.B(n_2069),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2436),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_L g2742 ( 
.A1(n_2328),
.A2(n_2185),
.B1(n_2090),
.B2(n_2069),
.Y(n_2742)
);

AND2x4_ASAP7_75t_L g2743 ( 
.A(n_2522),
.B(n_2090),
.Y(n_2743)
);

AND2x4_ASAP7_75t_L g2744 ( 
.A(n_2555),
.B(n_2156),
.Y(n_2744)
);

OR2x2_ASAP7_75t_SL g2745 ( 
.A(n_2463),
.B(n_1862),
.Y(n_2745)
);

AND2x4_ASAP7_75t_L g2746 ( 
.A(n_2555),
.B(n_2180),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2565),
.B(n_2180),
.Y(n_2747)
);

AOI22xp33_ASAP7_75t_L g2748 ( 
.A1(n_2516),
.A2(n_2185),
.B1(n_2180),
.B2(n_2035),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2467),
.B(n_2267),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2384),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2594),
.B(n_2185),
.Y(n_2751)
);

NAND2x1p5_ASAP7_75t_L g2752 ( 
.A(n_2306),
.B(n_1940),
.Y(n_2752)
);

INVx8_ASAP7_75t_L g2753 ( 
.A(n_2482),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2340),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_L g2755 ( 
.A(n_2413),
.B(n_1632),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2534),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2534),
.Y(n_2757)
);

INVx1_ASAP7_75t_SL g2758 ( 
.A(n_2349),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2565),
.B(n_2185),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2537),
.Y(n_2760)
);

INVxp67_ASAP7_75t_L g2761 ( 
.A(n_2680),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2537),
.Y(n_2762)
);

AND2x4_ASAP7_75t_L g2763 ( 
.A(n_2306),
.B(n_1823),
.Y(n_2763)
);

BUFx6f_ASAP7_75t_L g2764 ( 
.A(n_2314),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2540),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2539),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2384),
.Y(n_2767)
);

AOI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2452),
.A2(n_2311),
.B1(n_2399),
.B2(n_2307),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2520),
.B(n_1330),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2292),
.B(n_1382),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2539),
.Y(n_2771)
);

HB1xp67_ASAP7_75t_L g2772 ( 
.A(n_2529),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_2291),
.B(n_1679),
.Y(n_2773)
);

AND2x6_ASAP7_75t_L g2774 ( 
.A(n_2318),
.B(n_2154),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2384),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2452),
.B(n_2275),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2388),
.Y(n_2777)
);

BUFx2_ASAP7_75t_L g2778 ( 
.A(n_2637),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2323),
.B(n_2446),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2314),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2311),
.A2(n_2038),
.B1(n_2040),
.B2(n_2037),
.Y(n_2781)
);

AOI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2307),
.A2(n_2048),
.B1(n_2051),
.B2(n_2047),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_L g2783 ( 
.A1(n_2516),
.A2(n_2054),
.B1(n_2066),
.B2(n_2060),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2348),
.B(n_2067),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2544),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2451),
.B(n_1679),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2348),
.B(n_1705),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2499),
.B(n_1709),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2320),
.B(n_2347),
.Y(n_2789)
);

INVxp33_ASAP7_75t_L g2790 ( 
.A(n_2376),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2544),
.Y(n_2791)
);

OR2x2_ASAP7_75t_SL g2792 ( 
.A(n_2372),
.B(n_1810),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2388),
.Y(n_2793)
);

BUFx6f_ASAP7_75t_L g2794 ( 
.A(n_2401),
.Y(n_2794)
);

BUFx10_ASAP7_75t_L g2795 ( 
.A(n_2681),
.Y(n_2795)
);

AND2x4_ASAP7_75t_L g2796 ( 
.A(n_2473),
.B(n_2480),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2545),
.Y(n_2797)
);

INVxp67_ASAP7_75t_L g2798 ( 
.A(n_2543),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_SL g2799 ( 
.A(n_2484),
.B(n_1705),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2401),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2401),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2545),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2547),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2401),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2547),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2484),
.B(n_2192),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2548),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2548),
.Y(n_2808)
);

BUFx6f_ASAP7_75t_L g2809 ( 
.A(n_2402),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2506),
.B(n_2192),
.Y(n_2810)
);

INVx1_ASAP7_75t_SL g2811 ( 
.A(n_2289),
.Y(n_2811)
);

INVx3_ASAP7_75t_L g2812 ( 
.A(n_2402),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2402),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2506),
.B(n_2068),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2454),
.B(n_2192),
.Y(n_2815)
);

CKINVDCx5p33_ASAP7_75t_R g2816 ( 
.A(n_2332),
.Y(n_2816)
);

BUFx6f_ASAP7_75t_L g2817 ( 
.A(n_2402),
.Y(n_2817)
);

AND2x6_ASAP7_75t_L g2818 ( 
.A(n_2318),
.B(n_2154),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2563),
.Y(n_2819)
);

NAND2xp33_ASAP7_75t_L g2820 ( 
.A(n_2406),
.B(n_2076),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2590),
.B(n_2078),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2473),
.B(n_1823),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2563),
.Y(n_2823)
);

BUFx2_ASAP7_75t_L g2824 ( 
.A(n_2637),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2462),
.B(n_2079),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2406),
.Y(n_2826)
);

HB1xp67_ASAP7_75t_L g2827 ( 
.A(n_2435),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2570),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2406),
.Y(n_2829)
);

INVxp67_ASAP7_75t_L g2830 ( 
.A(n_2308),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2570),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2577),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2639),
.B(n_1709),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2577),
.Y(n_2834)
);

AND2x6_ASAP7_75t_L g2835 ( 
.A(n_2318),
.B(n_2160),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2357),
.B(n_2082),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2516),
.A2(n_2101),
.B1(n_2102),
.B2(n_2094),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2388),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2289),
.B(n_1457),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2585),
.Y(n_2840)
);

BUFx3_ASAP7_75t_L g2841 ( 
.A(n_2508),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_SL g2842 ( 
.A(n_2641),
.B(n_1813),
.Y(n_2842)
);

NAND2x1p5_ASAP7_75t_L g2843 ( 
.A(n_2480),
.B(n_2253),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2435),
.B(n_1487),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2585),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2589),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2589),
.Y(n_2847)
);

AOI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2516),
.A2(n_2109),
.B1(n_2111),
.B2(n_2106),
.Y(n_2848)
);

AND2x4_ASAP7_75t_L g2849 ( 
.A(n_2678),
.B(n_1825),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2421),
.Y(n_2850)
);

OR2x6_ASAP7_75t_L g2851 ( 
.A(n_2482),
.B(n_1714),
.Y(n_2851)
);

OAI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2574),
.A2(n_2114),
.B1(n_2121),
.B2(n_2112),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2406),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2593),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2593),
.Y(n_2855)
);

BUFx6f_ASAP7_75t_L g2856 ( 
.A(n_2475),
.Y(n_2856)
);

NAND2x1p5_ASAP7_75t_L g2857 ( 
.A(n_2689),
.B(n_2678),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2595),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2595),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2373),
.B(n_2125),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2475),
.Y(n_2861)
);

BUFx6f_ASAP7_75t_L g2862 ( 
.A(n_2475),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2598),
.Y(n_2863)
);

BUFx3_ASAP7_75t_L g2864 ( 
.A(n_2508),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2639),
.B(n_1810),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_2471),
.Y(n_2866)
);

NAND2x1p5_ASAP7_75t_L g2867 ( 
.A(n_2689),
.B(n_2253),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2598),
.Y(n_2868)
);

BUFx3_ASAP7_75t_L g2869 ( 
.A(n_2408),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2571),
.Y(n_2870)
);

INVx4_ASAP7_75t_L g2871 ( 
.A(n_2475),
.Y(n_2871)
);

INVx4_ASAP7_75t_L g2872 ( 
.A(n_2661),
.Y(n_2872)
);

INVx4_ASAP7_75t_SL g2873 ( 
.A(n_2444),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2421),
.Y(n_2874)
);

AND2x6_ASAP7_75t_L g2875 ( 
.A(n_2335),
.B(n_2421),
.Y(n_2875)
);

INVx8_ASAP7_75t_L g2876 ( 
.A(n_2482),
.Y(n_2876)
);

BUFx3_ASAP7_75t_L g2877 ( 
.A(n_2408),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2641),
.B(n_1813),
.Y(n_2878)
);

AOI22xp33_ASAP7_75t_SL g2879 ( 
.A1(n_2419),
.A2(n_2141),
.B1(n_1818),
.B2(n_2235),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_2558),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2579),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2422),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2558),
.B(n_1535),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2431),
.B(n_1818),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2315),
.A2(n_2128),
.B1(n_2132),
.B2(n_2127),
.Y(n_2885)
);

CKINVDCx20_ASAP7_75t_R g2886 ( 
.A(n_2296),
.Y(n_2886)
);

NAND2x1p5_ASAP7_75t_L g2887 ( 
.A(n_2672),
.B(n_2253),
.Y(n_2887)
);

OR2x2_ASAP7_75t_L g2888 ( 
.A(n_2441),
.B(n_2141),
.Y(n_2888)
);

HB1xp67_ASAP7_75t_L g2889 ( 
.A(n_2659),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2614),
.B(n_1736),
.Y(n_2890)
);

CKINVDCx20_ASAP7_75t_R g2891 ( 
.A(n_2296),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2672),
.B(n_2673),
.Y(n_2892)
);

INVx3_ASAP7_75t_L g2893 ( 
.A(n_2335),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2580),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2422),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2614),
.B(n_1383),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2591),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2422),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2596),
.Y(n_2899)
);

OAI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2339),
.A2(n_2136),
.B1(n_2137),
.B2(n_2133),
.Y(n_2900)
);

CKINVDCx20_ASAP7_75t_R g2901 ( 
.A(n_2287),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2597),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2560),
.B(n_2142),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2604),
.Y(n_2904)
);

BUFx6f_ASAP7_75t_L g2905 ( 
.A(n_2538),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2516),
.A2(n_2145),
.B1(n_2146),
.B2(n_2144),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2560),
.B(n_2147),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2290),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2290),
.Y(n_2909)
);

BUFx2_ASAP7_75t_L g2910 ( 
.A(n_2659),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2302),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2550),
.B(n_2588),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2302),
.Y(n_2913)
);

INVx2_ASAP7_75t_SL g2914 ( 
.A(n_2606),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2661),
.Y(n_2915)
);

BUFx6f_ASAP7_75t_L g2916 ( 
.A(n_2538),
.Y(n_2916)
);

OAI21xp33_ASAP7_75t_L g2917 ( 
.A1(n_2613),
.A2(n_1396),
.B(n_1390),
.Y(n_2917)
);

INVx4_ASAP7_75t_L g2918 ( 
.A(n_2661),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2645),
.B(n_1390),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2335),
.Y(n_2920)
);

INVx4_ASAP7_75t_L g2921 ( 
.A(n_2538),
.Y(n_2921)
);

OR2x2_ASAP7_75t_L g2922 ( 
.A(n_2441),
.B(n_1825),
.Y(n_2922)
);

INVx4_ASAP7_75t_L g2923 ( 
.A(n_2538),
.Y(n_2923)
);

INVx4_ASAP7_75t_L g2924 ( 
.A(n_2572),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2305),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2305),
.Y(n_2926)
);

HB1xp67_ASAP7_75t_L g2927 ( 
.A(n_2659),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2682),
.B(n_1826),
.Y(n_2928)
);

BUFx6f_ASAP7_75t_L g2929 ( 
.A(n_2572),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2550),
.B(n_1736),
.Y(n_2930)
);

OAI22xp33_ASAP7_75t_L g2931 ( 
.A1(n_2669),
.A2(n_2152),
.B1(n_2153),
.B2(n_2148),
.Y(n_2931)
);

AND2x4_ASAP7_75t_L g2932 ( 
.A(n_2684),
.B(n_1826),
.Y(n_2932)
);

INVx6_ASAP7_75t_L g2933 ( 
.A(n_2294),
.Y(n_2933)
);

NAND2x1p5_ASAP7_75t_L g2934 ( 
.A(n_2369),
.B(n_2157),
.Y(n_2934)
);

NOR2x1p5_ASAP7_75t_L g2935 ( 
.A(n_2379),
.B(n_1747),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2309),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2655),
.B(n_2159),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2309),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2321),
.Y(n_2939)
);

INVx4_ASAP7_75t_L g2940 ( 
.A(n_2572),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2321),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2488),
.B(n_1396),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2322),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2322),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2324),
.Y(n_2945)
);

INVx4_ASAP7_75t_L g2946 ( 
.A(n_2572),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2324),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2346),
.B(n_2161),
.Y(n_2948)
);

BUFx6f_ASAP7_75t_L g2949 ( 
.A(n_2622),
.Y(n_2949)
);

AND2x4_ASAP7_75t_L g2950 ( 
.A(n_2686),
.B(n_1826),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2329),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2329),
.Y(n_2952)
);

INVx2_ASAP7_75t_SL g2953 ( 
.A(n_2663),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_L g2954 ( 
.A(n_2622),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2330),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2445),
.B(n_1747),
.Y(n_2956)
);

INVx6_ASAP7_75t_L g2957 ( 
.A(n_2341),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2488),
.B(n_1445),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2581),
.B(n_2162),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2330),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_2557),
.B(n_2169),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_2622),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2331),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2331),
.Y(n_2964)
);

OR2x2_ASAP7_75t_SL g2965 ( 
.A(n_2674),
.B(n_1628),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_SL g2966 ( 
.A(n_2557),
.B(n_2170),
.Y(n_2966)
);

AND2x6_ASAP7_75t_L g2967 ( 
.A(n_2310),
.B(n_2160),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2333),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2333),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2361),
.B(n_1445),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2445),
.B(n_1471),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2345),
.Y(n_2972)
);

CKINVDCx5p33_ASAP7_75t_R g2973 ( 
.A(n_2375),
.Y(n_2973)
);

OA22x2_ASAP7_75t_L g2974 ( 
.A1(n_2317),
.A2(n_972),
.B1(n_995),
.B2(n_848),
.Y(n_2974)
);

BUFx3_ASAP7_75t_L g2975 ( 
.A(n_2482),
.Y(n_2975)
);

INVx4_ASAP7_75t_SL g2976 ( 
.A(n_2444),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_SL g2977 ( 
.A(n_2375),
.B(n_2235),
.Y(n_2977)
);

AO21x2_ASAP7_75t_L g2978 ( 
.A1(n_2647),
.A2(n_2178),
.B(n_2175),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2345),
.Y(n_2979)
);

AND2x6_ASAP7_75t_L g2980 ( 
.A(n_2310),
.B(n_2163),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2607),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2352),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_L g2983 ( 
.A(n_2458),
.B(n_1593),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2584),
.B(n_2182),
.Y(n_2984)
);

OR2x2_ASAP7_75t_L g2985 ( 
.A(n_2458),
.B(n_1835),
.Y(n_2985)
);

NAND2x1p5_ASAP7_75t_L g2986 ( 
.A(n_2369),
.B(n_2183),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2352),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2354),
.Y(n_2988)
);

CKINVDCx5p33_ASAP7_75t_R g2989 ( 
.A(n_2287),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2617),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2618),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2620),
.Y(n_2992)
);

BUFx6f_ASAP7_75t_L g2993 ( 
.A(n_2622),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2354),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2549),
.B(n_1593),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2549),
.B(n_1471),
.Y(n_2996)
);

BUFx6f_ASAP7_75t_L g2997 ( 
.A(n_2633),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2397),
.B(n_2187),
.Y(n_2998)
);

INVx4_ASAP7_75t_L g2999 ( 
.A(n_2633),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2621),
.Y(n_3000)
);

BUFx3_ASAP7_75t_L g3001 ( 
.A(n_2575),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2610),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2368),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2610),
.Y(n_3004)
);

INVx4_ASAP7_75t_L g3005 ( 
.A(n_2633),
.Y(n_3005)
);

AO22x2_ASAP7_75t_L g3006 ( 
.A1(n_2503),
.A2(n_2553),
.B1(n_2576),
.B2(n_2477),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2368),
.Y(n_3007)
);

INVxp33_ASAP7_75t_L g3008 ( 
.A(n_2666),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2377),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2377),
.Y(n_3010)
);

INVx3_ASAP7_75t_L g3011 ( 
.A(n_2607),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2380),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2380),
.Y(n_3013)
);

AND2x4_ASAP7_75t_L g3014 ( 
.A(n_2573),
.B(n_1835),
.Y(n_3014)
);

BUFx6f_ASAP7_75t_L g3015 ( 
.A(n_2633),
.Y(n_3015)
);

INVx3_ASAP7_75t_L g3016 ( 
.A(n_2607),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2658),
.B(n_2191),
.Y(n_3017)
);

INVx3_ASAP7_75t_L g3018 ( 
.A(n_2640),
.Y(n_3018)
);

AND2x4_ASAP7_75t_L g3019 ( 
.A(n_2573),
.B(n_1835),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2298),
.B(n_2163),
.Y(n_3020)
);

INVx5_ASAP7_75t_L g3021 ( 
.A(n_2341),
.Y(n_3021)
);

AOI21x1_ASAP7_75t_L g3022 ( 
.A1(n_2501),
.A2(n_2172),
.B(n_2168),
.Y(n_3022)
);

AND2x4_ASAP7_75t_SL g3023 ( 
.A(n_2367),
.B(n_2168),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2385),
.Y(n_3024)
);

BUFx6f_ASAP7_75t_L g3025 ( 
.A(n_2643),
.Y(n_3025)
);

OR2x2_ASAP7_75t_L g3026 ( 
.A(n_2683),
.B(n_1860),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2385),
.Y(n_3027)
);

HB1xp67_ASAP7_75t_L g3028 ( 
.A(n_2453),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2391),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_SL g3030 ( 
.A(n_2397),
.B(n_2172),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2631),
.B(n_1493),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2301),
.B(n_2316),
.Y(n_3032)
);

NAND2x1p5_ASAP7_75t_L g3033 ( 
.A(n_2369),
.B(n_2493),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_SL g3034 ( 
.A(n_2631),
.B(n_2174),
.Y(n_3034)
);

BUFx6f_ASAP7_75t_L g3035 ( 
.A(n_2643),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2643),
.Y(n_3036)
);

BUFx3_ASAP7_75t_L g3037 ( 
.A(n_2575),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2319),
.B(n_2327),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_2460),
.B(n_1860),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2530),
.B(n_2174),
.Y(n_3040)
);

AOI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2516),
.A2(n_2184),
.B1(n_2195),
.B2(n_2177),
.Y(n_3041)
);

AND2x4_ASAP7_75t_L g3042 ( 
.A(n_2464),
.B(n_1860),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2612),
.Y(n_3043)
);

BUFx6f_ASAP7_75t_L g3044 ( 
.A(n_2643),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2612),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2391),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2616),
.Y(n_3047)
);

NAND2x1p5_ASAP7_75t_L g3048 ( 
.A(n_2493),
.B(n_2277),
.Y(n_3048)
);

AND2x4_ASAP7_75t_L g3049 ( 
.A(n_2472),
.B(n_1891),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2394),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2483),
.B(n_1493),
.Y(n_3051)
);

BUFx6f_ASAP7_75t_L g3052 ( 
.A(n_2367),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2490),
.B(n_1525),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_2434),
.A2(n_2184),
.B1(n_2195),
.B2(n_2177),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_2477),
.B(n_2428),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2492),
.B(n_1525),
.Y(n_3056)
);

INVx4_ASAP7_75t_L g3057 ( 
.A(n_2500),
.Y(n_3057)
);

AO22x2_ASAP7_75t_L g3058 ( 
.A1(n_2576),
.A2(n_1077),
.B1(n_1082),
.B2(n_1080),
.Y(n_3058)
);

BUFx10_ASAP7_75t_L g3059 ( 
.A(n_2300),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2394),
.Y(n_3060)
);

INVx3_ASAP7_75t_L g3061 ( 
.A(n_2640),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2395),
.Y(n_3062)
);

BUFx6f_ASAP7_75t_L g3063 ( 
.A(n_2367),
.Y(n_3063)
);

INVx4_ASAP7_75t_L g3064 ( 
.A(n_2500),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2395),
.Y(n_3065)
);

AND2x4_ASAP7_75t_L g3066 ( 
.A(n_2496),
.B(n_1891),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2398),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2398),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_2582),
.B(n_1696),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2400),
.Y(n_3070)
);

AND2x6_ASAP7_75t_L g3071 ( 
.A(n_2310),
.B(n_2197),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2400),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2404),
.Y(n_3073)
);

INVx8_ASAP7_75t_L g3074 ( 
.A(n_2444),
.Y(n_3074)
);

INVx4_ASAP7_75t_SL g3075 ( 
.A(n_2513),
.Y(n_3075)
);

NAND3x1_ASAP7_75t_L g3076 ( 
.A(n_2519),
.B(n_1082),
.C(n_1080),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_2912),
.B(n_2530),
.Y(n_3077)
);

CKINVDCx11_ASAP7_75t_R g3078 ( 
.A(n_2886),
.Y(n_3078)
);

AOI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2779),
.A2(n_2485),
.B1(n_2434),
.B2(n_2667),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_2798),
.B(n_2523),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_SL g3081 ( 
.A(n_2709),
.B(n_2530),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2776),
.B(n_2507),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_SL g3083 ( 
.A(n_2744),
.B(n_2418),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2691),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2691),
.Y(n_3085)
);

NOR2xp33_ASAP7_75t_L g3086 ( 
.A(n_3008),
.B(n_2285),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2768),
.B(n_2515),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2692),
.Y(n_3088)
);

OR2x2_ASAP7_75t_L g3089 ( 
.A(n_2705),
.B(n_2667),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2789),
.B(n_2366),
.Y(n_3090)
);

AOI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_3055),
.A2(n_2485),
.B1(n_2285),
.B2(n_2505),
.Y(n_3091)
);

BUFx3_ASAP7_75t_L g3092 ( 
.A(n_2699),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2693),
.B(n_2312),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2825),
.B(n_2312),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2827),
.B(n_2312),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2905),
.Y(n_3096)
);

INVx2_ASAP7_75t_SL g3097 ( 
.A(n_2702),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2692),
.Y(n_3098)
);

OR2x2_ASAP7_75t_L g3099 ( 
.A(n_2811),
.B(n_2285),
.Y(n_3099)
);

NOR2xp33_ASAP7_75t_L g3100 ( 
.A(n_2786),
.B(n_2285),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2703),
.B(n_2313),
.Y(n_3101)
);

AOI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2734),
.A2(n_2755),
.B1(n_2485),
.B2(n_2914),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2761),
.B(n_2383),
.Y(n_3103)
);

OAI22xp5_ASAP7_75t_SL g3104 ( 
.A1(n_2879),
.A2(n_2502),
.B1(n_2636),
.B2(n_2519),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2697),
.Y(n_3105)
);

INVxp67_ASAP7_75t_L g3106 ( 
.A(n_2739),
.Y(n_3106)
);

AOI22xp33_ASAP7_75t_L g3107 ( 
.A1(n_2888),
.A2(n_2485),
.B1(n_2518),
.B2(n_2510),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2703),
.B(n_2313),
.Y(n_3108)
);

OAI22xp5_ASAP7_75t_L g3109 ( 
.A1(n_2751),
.A2(n_2556),
.B1(n_2600),
.B2(n_2390),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2696),
.A2(n_2424),
.B(n_2326),
.Y(n_3110)
);

BUFx6f_ASAP7_75t_SL g3111 ( 
.A(n_2841),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2703),
.B(n_2313),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2703),
.B(n_2485),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2892),
.A2(n_2485),
.B1(n_2527),
.B2(n_2521),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2717),
.B(n_2884),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2744),
.B(n_2383),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2821),
.B(n_2536),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2697),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2704),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2704),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2880),
.B(n_2502),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2707),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_3031),
.B(n_2334),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_SL g3124 ( 
.A(n_2746),
.B(n_2493),
.Y(n_3124)
);

NOR2xp33_ASAP7_75t_L g3125 ( 
.A(n_2758),
.B(n_2665),
.Y(n_3125)
);

NOR2x1p5_ASAP7_75t_L g3126 ( 
.A(n_2864),
.B(n_2427),
.Y(n_3126)
);

NAND3xp33_ASAP7_75t_SL g3127 ( 
.A(n_2773),
.B(n_2487),
.C(n_2427),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_SL g3128 ( 
.A(n_2746),
.B(n_2514),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2707),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_L g3130 ( 
.A(n_2713),
.B(n_2668),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2708),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2770),
.B(n_2336),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2919),
.B(n_2532),
.Y(n_3133)
);

AOI22xp5_ASAP7_75t_L g3134 ( 
.A1(n_2910),
.A2(n_2535),
.B1(n_2603),
.B2(n_2592),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2708),
.Y(n_3135)
);

OAI21xp5_ASAP7_75t_L g3136 ( 
.A1(n_2948),
.A2(n_2420),
.B(n_2469),
.Y(n_3136)
);

NOR2xp33_ASAP7_75t_L g3137 ( 
.A(n_2722),
.B(n_2338),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2712),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2747),
.B(n_2514),
.Y(n_3139)
);

BUFx8_ASAP7_75t_L g3140 ( 
.A(n_2778),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_L g3141 ( 
.A(n_2732),
.B(n_2343),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_2747),
.B(n_2514),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2942),
.B(n_2660),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2958),
.B(n_2662),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2917),
.B(n_2350),
.Y(n_3145)
);

O2A1O1Ixp5_ASAP7_75t_L g3146 ( 
.A1(n_2749),
.A2(n_2360),
.B(n_2387),
.C(n_2337),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_2892),
.A2(n_2351),
.B1(n_2358),
.B2(n_2353),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2712),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_3014),
.B(n_2359),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_2724),
.B(n_2364),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_3014),
.B(n_2370),
.Y(n_3151)
);

AOI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_3017),
.A2(n_2424),
.B(n_2326),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2718),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_2701),
.B(n_2371),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2844),
.B(n_2971),
.Y(n_3155)
);

OR2x2_ASAP7_75t_L g3156 ( 
.A(n_2765),
.B(n_2381),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2996),
.B(n_2382),
.Y(n_3157)
);

A2O1A1Ixp33_ASAP7_75t_L g3158 ( 
.A1(n_2736),
.A2(n_2390),
.B(n_2600),
.C(n_2556),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2718),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2836),
.B(n_2541),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2725),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2725),
.Y(n_3162)
);

NAND2x1p5_ASAP7_75t_L g3163 ( 
.A(n_2727),
.B(n_2390),
.Y(n_3163)
);

INVxp67_ASAP7_75t_L g3164 ( 
.A(n_2754),
.Y(n_3164)
);

AND2x4_ASAP7_75t_L g3165 ( 
.A(n_2796),
.B(n_2386),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2860),
.B(n_2542),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_3019),
.B(n_2392),
.Y(n_3167)
);

AND2x6_ASAP7_75t_SL g3168 ( 
.A(n_3069),
.B(n_2575),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_2830),
.B(n_2393),
.Y(n_3169)
);

O2A1O1Ixp33_ASAP7_75t_L g3170 ( 
.A1(n_2970),
.A2(n_2688),
.B(n_2425),
.C(n_2626),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2726),
.B(n_2546),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2726),
.Y(n_3172)
);

NOR2x1p5_ASAP7_75t_L g3173 ( 
.A(n_2869),
.B(n_2487),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2797),
.Y(n_3174)
);

INVx4_ASAP7_75t_L g3175 ( 
.A(n_2856),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_2737),
.Y(n_3176)
);

AOI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_3019),
.A2(n_2609),
.B1(n_2615),
.B2(n_2396),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2738),
.B(n_2629),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2797),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2769),
.B(n_2448),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2741),
.B(n_2634),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2802),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_3032),
.B(n_2635),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2802),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_3038),
.B(n_2650),
.Y(n_3185)
);

AOI22xp33_ASAP7_75t_L g3186 ( 
.A1(n_2974),
.A2(n_2646),
.B1(n_2651),
.B2(n_2638),
.Y(n_3186)
);

OAI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_2729),
.A2(n_2600),
.B1(n_2556),
.B2(n_2420),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2803),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_3051),
.B(n_2438),
.Y(n_3189)
);

A2O1A1Ixp33_ASAP7_75t_L g3190 ( 
.A1(n_2937),
.A2(n_2675),
.B(n_2559),
.C(n_2562),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_3053),
.B(n_2440),
.Y(n_3191)
);

INVxp67_ASAP7_75t_L g3192 ( 
.A(n_2839),
.Y(n_3192)
);

OAI22xp33_ASAP7_75t_L g3193 ( 
.A1(n_2985),
.A2(n_2365),
.B1(n_2355),
.B2(n_2575),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_3056),
.B(n_2442),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2896),
.B(n_2447),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2803),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2690),
.B(n_2326),
.Y(n_3197)
);

NOR3xp33_ASAP7_75t_L g3198 ( 
.A(n_2788),
.B(n_2625),
.C(n_2360),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_SL g3199 ( 
.A(n_2690),
.B(n_2326),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2870),
.B(n_2649),
.Y(n_3200)
);

BUFx6f_ASAP7_75t_L g3201 ( 
.A(n_2905),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2805),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2805),
.Y(n_3203)
);

A2O1A1Ixp33_ASAP7_75t_L g3204 ( 
.A1(n_2881),
.A2(n_2551),
.B(n_2568),
.C(n_2566),
.Y(n_3204)
);

OAI22xp33_ASAP7_75t_L g3205 ( 
.A1(n_2922),
.A2(n_2365),
.B1(n_2355),
.B2(n_2500),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_L g3206 ( 
.A1(n_2894),
.A2(n_2899),
.B1(n_2902),
.B2(n_2897),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2904),
.B(n_2649),
.Y(n_3207)
);

O2A1O1Ixp5_ASAP7_75t_L g3208 ( 
.A1(n_2885),
.A2(n_2387),
.B(n_2337),
.C(n_2608),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2807),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_2772),
.B(n_2866),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2990),
.B(n_2652),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_SL g3212 ( 
.A(n_2695),
.B(n_2326),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2807),
.B(n_2616),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2808),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_L g3215 ( 
.A(n_2883),
.B(n_2355),
.Y(n_3215)
);

AOI22xp33_ASAP7_75t_L g3216 ( 
.A1(n_2991),
.A2(n_2448),
.B1(n_2653),
.B2(n_2652),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_L g3217 ( 
.A(n_2795),
.B(n_2355),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2808),
.B(n_2619),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_2795),
.B(n_2365),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2908),
.B(n_2619),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2908),
.B(n_2623),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2909),
.B(n_2623),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2909),
.B(n_2624),
.Y(n_3223)
);

A2O1A1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_2992),
.A2(n_2654),
.B(n_2653),
.C(n_2627),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_2790),
.B(n_2365),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2911),
.B(n_2624),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2911),
.B(n_2627),
.Y(n_3227)
);

AOI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_2889),
.A2(n_2448),
.B1(n_2342),
.B2(n_2671),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2913),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_2973),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2913),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2925),
.Y(n_3232)
);

OAI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_2959),
.A2(n_2469),
.B(n_2417),
.Y(n_3233)
);

OR2x2_ASAP7_75t_L g3234 ( 
.A(n_3026),
.B(n_2654),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_SL g3235 ( 
.A(n_2695),
.B(n_2424),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_2700),
.B(n_2424),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2925),
.Y(n_3237)
);

INVxp33_ASAP7_75t_L g3238 ( 
.A(n_2890),
.Y(n_3238)
);

A2O1A1Ixp33_ASAP7_75t_L g3239 ( 
.A1(n_3000),
.A2(n_2630),
.B(n_2500),
.C(n_2299),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2938),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2938),
.Y(n_3241)
);

AND2x4_ASAP7_75t_SL g3242 ( 
.A(n_2872),
.B(n_2630),
.Y(n_3242)
);

AND2x2_ASAP7_75t_SL g3243 ( 
.A(n_2721),
.B(n_2552),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_SL g3244 ( 
.A(n_2700),
.B(n_2424),
.Y(n_3244)
);

NOR2xp33_ASAP7_75t_SL g3245 ( 
.A(n_2989),
.B(n_2676),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2939),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2939),
.Y(n_3247)
);

NOR2xp33_ASAP7_75t_L g3248 ( 
.A(n_2930),
.B(n_2513),
.Y(n_3248)
);

OAI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_2953),
.A2(n_2564),
.B1(n_2628),
.B2(n_2504),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_2731),
.B(n_2491),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2941),
.B(n_2404),
.Y(n_3251)
);

BUFx6f_ASAP7_75t_L g3252 ( 
.A(n_2905),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2941),
.Y(n_3253)
);

OR2x6_ASAP7_75t_L g3254 ( 
.A(n_2720),
.B(n_3074),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_2731),
.B(n_2491),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2956),
.B(n_2513),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2944),
.B(n_2407),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2740),
.B(n_2494),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_SL g3259 ( 
.A(n_2740),
.B(n_2743),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_2944),
.B(n_2407),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2945),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2743),
.B(n_2849),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_SL g3263 ( 
.A(n_2849),
.B(n_2491),
.Y(n_3263)
);

O2A1O1Ixp5_ASAP7_75t_L g3264 ( 
.A1(n_2900),
.A2(n_2295),
.B(n_2286),
.C(n_2656),
.Y(n_3264)
);

AOI22xp33_ASAP7_75t_L g3265 ( 
.A1(n_3039),
.A2(n_2342),
.B1(n_2625),
.B2(n_2656),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2945),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2947),
.B(n_2409),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_2737),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2947),
.B(n_2409),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2951),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2951),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_2833),
.B(n_2465),
.Y(n_3272)
);

O2A1O1Ixp5_ASAP7_75t_L g3273 ( 
.A1(n_2815),
.A2(n_2679),
.B(n_2685),
.C(n_2677),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2952),
.B(n_2410),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_2952),
.B(n_2410),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2955),
.B(n_2414),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_2737),
.Y(n_3277)
);

AOI22xp33_ASAP7_75t_L g3278 ( 
.A1(n_3039),
.A2(n_2342),
.B1(n_2679),
.B2(n_2677),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2955),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3002),
.B(n_2414),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3004),
.B(n_2416),
.Y(n_3281)
);

BUFx2_ASAP7_75t_L g3282 ( 
.A(n_2711),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2960),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_2960),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_3043),
.B(n_2416),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3045),
.B(n_3047),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_3042),
.A2(n_2685),
.B1(n_2299),
.B2(n_2561),
.Y(n_3287)
);

NOR3xp33_ASAP7_75t_L g3288 ( 
.A(n_2842),
.B(n_2564),
.C(n_2504),
.Y(n_3288)
);

NOR3xp33_ASAP7_75t_L g3289 ( 
.A(n_2878),
.B(n_2628),
.C(n_2569),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_2865),
.B(n_1696),
.Y(n_3290)
);

BUFx6f_ASAP7_75t_L g3291 ( 
.A(n_2916),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2964),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2964),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3042),
.A2(n_2561),
.B1(n_2602),
.B2(n_2601),
.Y(n_3294)
);

AOI22xp33_ASAP7_75t_L g3295 ( 
.A1(n_3049),
.A2(n_2561),
.B1(n_2602),
.B2(n_2601),
.Y(n_3295)
);

BUFx3_ASAP7_75t_L g3296 ( 
.A(n_3074),
.Y(n_3296)
);

NOR3xp33_ASAP7_75t_L g3297 ( 
.A(n_2787),
.B(n_2569),
.C(n_2676),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_L g3298 ( 
.A(n_2927),
.B(n_1701),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3049),
.B(n_2426),
.Y(n_3299)
);

AO22x1_ASAP7_75t_L g3300 ( 
.A1(n_2983),
.A2(n_887),
.B1(n_889),
.B2(n_879),
.Y(n_3300)
);

NAND2x1p5_ASAP7_75t_L g3301 ( 
.A(n_2727),
.B(n_2640),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2968),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_2872),
.B(n_2657),
.Y(n_3303)
);

CKINVDCx5p33_ASAP7_75t_R g3304 ( 
.A(n_2816),
.Y(n_3304)
);

AOI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_3066),
.A2(n_2605),
.B1(n_2430),
.B2(n_2433),
.Y(n_3305)
);

AND2x4_ASAP7_75t_L g3306 ( 
.A(n_2796),
.B(n_2644),
.Y(n_3306)
);

INVx2_ASAP7_75t_SL g3307 ( 
.A(n_2763),
.Y(n_3307)
);

AND2x4_ASAP7_75t_L g3308 ( 
.A(n_2763),
.B(n_2644),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_SL g3309 ( 
.A(n_2915),
.B(n_2657),
.Y(n_3309)
);

BUFx6f_ASAP7_75t_SL g3310 ( 
.A(n_2877),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3066),
.B(n_2426),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_2968),
.Y(n_3312)
);

AOI22xp33_ASAP7_75t_L g3313 ( 
.A1(n_2928),
.A2(n_2605),
.B1(n_2433),
.B2(n_2437),
.Y(n_3313)
);

NOR2xp33_ASAP7_75t_R g3314 ( 
.A(n_2735),
.B(n_2644),
.Y(n_3314)
);

INVx4_ASAP7_75t_L g3315 ( 
.A(n_2856),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_SL g3316 ( 
.A(n_2977),
.B(n_1701),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2969),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3028),
.B(n_2784),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2969),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_2928),
.A2(n_2437),
.B1(n_2439),
.B2(n_2430),
.Y(n_3320)
);

AOI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3006),
.A2(n_2325),
.B1(n_2403),
.B2(n_2344),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2982),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2814),
.B(n_2714),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2714),
.B(n_2439),
.Y(n_3324)
);

INVx3_ASAP7_75t_L g3325 ( 
.A(n_2764),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_L g3326 ( 
.A(n_2995),
.B(n_1876),
.Y(n_3326)
);

INVxp67_ASAP7_75t_L g3327 ( 
.A(n_2822),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2982),
.B(n_2457),
.Y(n_3328)
);

NOR2xp67_ASAP7_75t_L g3329 ( 
.A(n_2719),
.B(n_2648),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_2915),
.B(n_2554),
.Y(n_3330)
);

BUFx6f_ASAP7_75t_L g3331 ( 
.A(n_2916),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3010),
.Y(n_3332)
);

INVx2_ASAP7_75t_SL g3333 ( 
.A(n_2822),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3010),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3013),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3013),
.Y(n_3336)
);

INVx4_ASAP7_75t_L g3337 ( 
.A(n_2856),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2801),
.B(n_2457),
.Y(n_3338)
);

HB1xp67_ASAP7_75t_L g3339 ( 
.A(n_2932),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_2965),
.B(n_2648),
.Y(n_3340)
);

AND2x4_ASAP7_75t_L g3341 ( 
.A(n_2873),
.B(n_2648),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3024),
.Y(n_3342)
);

AOI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_3006),
.A2(n_2759),
.B1(n_2950),
.B2(n_2932),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_2801),
.B(n_2459),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3024),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_2812),
.B(n_2459),
.Y(n_3346)
);

BUFx6f_ASAP7_75t_L g3347 ( 
.A(n_2916),
.Y(n_3347)
);

NAND3xp33_ASAP7_75t_SL g3348 ( 
.A(n_2799),
.B(n_893),
.C(n_890),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2812),
.B(n_2461),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2829),
.B(n_2461),
.Y(n_3350)
);

CKINVDCx20_ASAP7_75t_R g3351 ( 
.A(n_2901),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3029),
.Y(n_3352)
);

A2O1A1Ixp33_ASAP7_75t_L g3353 ( 
.A1(n_2742),
.A2(n_2587),
.B(n_2664),
.C(n_2552),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2829),
.B(n_2466),
.Y(n_3354)
);

OAI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_2748),
.A2(n_2456),
.B1(n_2455),
.B2(n_2378),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2950),
.B(n_2466),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3029),
.Y(n_3357)
);

AOI22xp33_ASAP7_75t_L g3358 ( 
.A1(n_2759),
.A2(n_2476),
.B1(n_2478),
.B2(n_2468),
.Y(n_3358)
);

NOR3xp33_ASAP7_75t_L g3359 ( 
.A(n_3040),
.B(n_2824),
.C(n_2918),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3062),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3062),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3068),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_2723),
.B(n_1785),
.Y(n_3363)
);

OAI22xp5_ASAP7_75t_L g3364 ( 
.A1(n_2984),
.A2(n_2728),
.B1(n_2893),
.B2(n_2783),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_2745),
.B(n_2918),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2728),
.B(n_2468),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_L g3367 ( 
.A(n_2893),
.B(n_2476),
.Y(n_3367)
);

INVx3_ASAP7_75t_L g3368 ( 
.A(n_2764),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3068),
.B(n_2478),
.Y(n_3369)
);

INVx8_ASAP7_75t_L g3370 ( 
.A(n_2720),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3070),
.Y(n_3371)
);

OAI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_2750),
.A2(n_2456),
.B1(n_2455),
.B2(n_2378),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3070),
.B(n_2479),
.Y(n_3373)
);

OAI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_2694),
.A2(n_2481),
.B1(n_2486),
.B2(n_2479),
.Y(n_3374)
);

NAND2x1_ASAP7_75t_L g3375 ( 
.A(n_3057),
.B(n_2583),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3072),
.B(n_2481),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3072),
.B(n_2486),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2926),
.B(n_2489),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3058),
.A2(n_2498),
.B1(n_2511),
.B2(n_2509),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_2706),
.B(n_2554),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2936),
.B(n_2489),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_2943),
.B(n_2498),
.Y(n_3382)
);

INVx2_ASAP7_75t_SL g3383 ( 
.A(n_2957),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_2963),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_SL g3385 ( 
.A(n_2706),
.B(n_2554),
.Y(n_3385)
);

AOI22xp5_ASAP7_75t_L g3386 ( 
.A1(n_2998),
.A2(n_2344),
.B1(n_2403),
.B2(n_2325),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_L g3387 ( 
.A1(n_3058),
.A2(n_2511),
.B1(n_2509),
.B2(n_2531),
.Y(n_3387)
);

BUFx3_ASAP7_75t_L g3388 ( 
.A(n_3052),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_2972),
.B(n_2389),
.Y(n_3389)
);

INVx2_ASAP7_75t_SL g3390 ( 
.A(n_2957),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_3033),
.A2(n_2586),
.B(n_2583),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_2698),
.B(n_2455),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_L g3393 ( 
.A(n_2792),
.B(n_2767),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_SL g3394 ( 
.A(n_2891),
.B(n_2578),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2775),
.B(n_2456),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_2777),
.B(n_2363),
.Y(n_3396)
);

NAND2x1p5_ASAP7_75t_L g3397 ( 
.A(n_2710),
.B(n_2583),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2756),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2793),
.B(n_2363),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2838),
.B(n_2363),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_2757),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2850),
.B(n_2378),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2874),
.B(n_2197),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2760),
.Y(n_3404)
);

NOR3xp33_ASAP7_75t_SL g3405 ( 
.A(n_3030),
.B(n_897),
.C(n_896),
.Y(n_3405)
);

AOI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_2882),
.A2(n_2531),
.B1(n_2206),
.B2(n_2211),
.Y(n_3406)
);

NOR2xp67_ASAP7_75t_L g3407 ( 
.A(n_3021),
.B(n_2206),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_2895),
.B(n_2207),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2898),
.B(n_2207),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2762),
.Y(n_3410)
);

INVx8_ASAP7_75t_L g3411 ( 
.A(n_2753),
.Y(n_3411)
);

BUFx3_ASAP7_75t_L g3412 ( 
.A(n_3052),
.Y(n_3412)
);

BUFx4_ASAP7_75t_L g3413 ( 
.A(n_2873),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_2979),
.Y(n_3414)
);

AOI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_2903),
.A2(n_2586),
.B(n_2524),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2920),
.B(n_2211),
.Y(n_3416)
);

INVxp67_ASAP7_75t_L g3417 ( 
.A(n_3001),
.Y(n_3417)
);

INVxp67_ASAP7_75t_L g3418 ( 
.A(n_3037),
.Y(n_3418)
);

AOI22xp5_ASAP7_75t_L g3419 ( 
.A1(n_2961),
.A2(n_2664),
.B1(n_2587),
.B2(n_884),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2766),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_2976),
.B(n_1785),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_2706),
.B(n_2578),
.Y(n_3422)
);

AND2x4_ASAP7_75t_L g3423 ( 
.A(n_2976),
.B(n_2531),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2771),
.B(n_2212),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2785),
.B(n_2212),
.Y(n_3425)
);

INVxp67_ASAP7_75t_SL g3426 ( 
.A(n_2764),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_2987),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3075),
.B(n_1785),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2791),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_2819),
.B(n_2213),
.Y(n_3430)
);

NOR2x1p5_ASAP7_75t_L g3431 ( 
.A(n_2975),
.B(n_1403),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_2823),
.B(n_2213),
.Y(n_3432)
);

NAND2xp33_ASAP7_75t_L g3433 ( 
.A(n_2780),
.B(n_2524),
.Y(n_3433)
);

AOI22xp33_ASAP7_75t_L g3434 ( 
.A1(n_2966),
.A2(n_2217),
.B1(n_2229),
.B2(n_2220),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_SL g3435 ( 
.A(n_2721),
.B(n_2578),
.Y(n_3435)
);

INVxp33_ASAP7_75t_L g3436 ( 
.A(n_2733),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3075),
.B(n_2470),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2988),
.Y(n_3438)
);

O2A1O1Ixp33_ASAP7_75t_L g3439 ( 
.A1(n_3020),
.A2(n_2931),
.B(n_3034),
.C(n_2852),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_2780),
.B(n_2794),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3180),
.B(n_3133),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_L g3442 ( 
.A(n_3115),
.B(n_2694),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_L g3443 ( 
.A(n_3238),
.B(n_2694),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3398),
.Y(n_3444)
);

BUFx2_ASAP7_75t_L g3445 ( 
.A(n_3092),
.Y(n_3445)
);

INVxp67_ASAP7_75t_SL g3446 ( 
.A(n_3106),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3085),
.Y(n_3447)
);

BUFx8_ASAP7_75t_L g3448 ( 
.A(n_3111),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3401),
.Y(n_3449)
);

BUFx12f_ASAP7_75t_L g3450 ( 
.A(n_3078),
.Y(n_3450)
);

BUFx3_ASAP7_75t_L g3451 ( 
.A(n_3296),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3404),
.Y(n_3452)
);

INVx1_ASAP7_75t_SL g3453 ( 
.A(n_3150),
.Y(n_3453)
);

NOR2xp67_ASAP7_75t_L g3454 ( 
.A(n_3102),
.B(n_2871),
.Y(n_3454)
);

CKINVDCx6p67_ASAP7_75t_R g3455 ( 
.A(n_3111),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3410),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3098),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3096),
.Y(n_3458)
);

OR2x2_ASAP7_75t_L g3459 ( 
.A(n_3155),
.B(n_2752),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3420),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_3137),
.B(n_3021),
.Y(n_3461)
);

INVx3_ASAP7_75t_L g3462 ( 
.A(n_3437),
.Y(n_3462)
);

BUFx3_ASAP7_75t_L g3463 ( 
.A(n_3388),
.Y(n_3463)
);

INVxp67_ASAP7_75t_L g3464 ( 
.A(n_3125),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3429),
.Y(n_3465)
);

INVxp67_ASAP7_75t_SL g3466 ( 
.A(n_3164),
.Y(n_3466)
);

BUFx4f_ASAP7_75t_L g3467 ( 
.A(n_3370),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3082),
.B(n_2828),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3084),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_3314),
.Y(n_3470)
);

INVxp67_ASAP7_75t_L g3471 ( 
.A(n_3141),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3192),
.B(n_2857),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_3230),
.Y(n_3473)
);

BUFx6f_ASAP7_75t_L g3474 ( 
.A(n_3096),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3105),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3088),
.Y(n_3476)
);

CKINVDCx11_ASAP7_75t_R g3477 ( 
.A(n_3351),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3119),
.Y(n_3478)
);

CKINVDCx5p33_ASAP7_75t_R g3479 ( 
.A(n_3304),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_SL g3480 ( 
.A(n_3132),
.B(n_3021),
.Y(n_3480)
);

HB1xp67_ASAP7_75t_L g3481 ( 
.A(n_3097),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3118),
.Y(n_3482)
);

BUFx6f_ASAP7_75t_L g3483 ( 
.A(n_3096),
.Y(n_3483)
);

INVx6_ASAP7_75t_L g3484 ( 
.A(n_3140),
.Y(n_3484)
);

INVx2_ASAP7_75t_SL g3485 ( 
.A(n_3412),
.Y(n_3485)
);

INVx3_ASAP7_75t_L g3486 ( 
.A(n_3437),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3131),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3183),
.B(n_2710),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3185),
.B(n_2716),
.Y(n_3489)
);

NAND3xp33_ASAP7_75t_L g3490 ( 
.A(n_3100),
.B(n_2781),
.C(n_2782),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3120),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_3169),
.B(n_2780),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3122),
.Y(n_3493)
);

HB1xp67_ASAP7_75t_L g3494 ( 
.A(n_3156),
.Y(n_3494)
);

INVx1_ASAP7_75t_SL g3495 ( 
.A(n_3089),
.Y(n_3495)
);

AOI221xp5_ASAP7_75t_L g3496 ( 
.A1(n_3080),
.A2(n_904),
.B1(n_912),
.B2(n_908),
.C(n_901),
.Y(n_3496)
);

INVxp67_ASAP7_75t_SL g3497 ( 
.A(n_3095),
.Y(n_3497)
);

AND2x4_ASAP7_75t_SL g3498 ( 
.A(n_3254),
.B(n_2871),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3135),
.Y(n_3499)
);

INVx2_ASAP7_75t_SL g3500 ( 
.A(n_3383),
.Y(n_3500)
);

HB1xp67_ASAP7_75t_L g3501 ( 
.A(n_3234),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3129),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3138),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3148),
.Y(n_3504)
);

AOI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3079),
.A2(n_3076),
.B1(n_2730),
.B2(n_2876),
.Y(n_3505)
);

BUFx6f_ASAP7_75t_L g3506 ( 
.A(n_3201),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3153),
.Y(n_3507)
);

NOR2x1p5_ASAP7_75t_SL g3508 ( 
.A(n_3172),
.B(n_3022),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3179),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_3210),
.B(n_3052),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3159),
.Y(n_3511)
);

BUFx2_ASAP7_75t_L g3512 ( 
.A(n_3282),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3161),
.Y(n_3513)
);

CKINVDCx5p33_ASAP7_75t_R g3514 ( 
.A(n_3140),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3162),
.Y(n_3515)
);

BUFx2_ASAP7_75t_L g3516 ( 
.A(n_3165),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3182),
.Y(n_3517)
);

O2A1O1Ixp33_ASAP7_75t_L g3518 ( 
.A1(n_3077),
.A2(n_2820),
.B(n_1096),
.C(n_1100),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_3310),
.Y(n_3519)
);

INVx3_ASAP7_75t_L g3520 ( 
.A(n_3306),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3174),
.Y(n_3521)
);

BUFx3_ASAP7_75t_L g3522 ( 
.A(n_3390),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3209),
.Y(n_3523)
);

INVx2_ASAP7_75t_SL g3524 ( 
.A(n_3413),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3184),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3121),
.B(n_3063),
.Y(n_3526)
);

INVx3_ASAP7_75t_SL g3527 ( 
.A(n_3254),
.Y(n_3527)
);

INVx5_ASAP7_75t_L g3528 ( 
.A(n_3201),
.Y(n_3528)
);

BUFx6f_ASAP7_75t_L g3529 ( 
.A(n_3201),
.Y(n_3529)
);

BUFx3_ASAP7_75t_L g3530 ( 
.A(n_3370),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3082),
.B(n_2831),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3188),
.Y(n_3532)
);

AOI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3215),
.A2(n_2876),
.B1(n_2753),
.B2(n_2907),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3117),
.B(n_2832),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3117),
.B(n_2834),
.Y(n_3535)
);

AND2x4_ASAP7_75t_L g3536 ( 
.A(n_3262),
.B(n_3023),
.Y(n_3536)
);

AOI21x1_ASAP7_75t_L g3537 ( 
.A1(n_3329),
.A2(n_2450),
.B(n_2449),
.Y(n_3537)
);

INVx4_ASAP7_75t_L g3538 ( 
.A(n_3370),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3196),
.Y(n_3539)
);

OAI22xp33_ASAP7_75t_L g3540 ( 
.A1(n_3316),
.A2(n_2715),
.B1(n_2851),
.B2(n_3063),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3202),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3232),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3237),
.Y(n_3543)
);

NOR2xp67_ASAP7_75t_L g3544 ( 
.A(n_3091),
.B(n_2716),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3160),
.B(n_2994),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3203),
.Y(n_3546)
);

OAI22xp33_ASAP7_75t_L g3547 ( 
.A1(n_3228),
.A2(n_2715),
.B1(n_2851),
.B2(n_3063),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3214),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3160),
.B(n_2840),
.Y(n_3549)
);

BUFx2_ASAP7_75t_L g3550 ( 
.A(n_3165),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3123),
.B(n_1803),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3240),
.Y(n_3552)
);

OAI22xp5_ASAP7_75t_SL g3553 ( 
.A1(n_3104),
.A2(n_915),
.B1(n_922),
.B2(n_917),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3248),
.B(n_3318),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_3103),
.B(n_2794),
.Y(n_3555)
);

INVx2_ASAP7_75t_SL g3556 ( 
.A(n_3431),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3247),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3166),
.B(n_2845),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3229),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3231),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3241),
.Y(n_3561)
);

INVx2_ASAP7_75t_SL g3562 ( 
.A(n_3258),
.Y(n_3562)
);

INVxp33_ASAP7_75t_L g3563 ( 
.A(n_3393),
.Y(n_3563)
);

BUFx6f_ASAP7_75t_L g3564 ( 
.A(n_3252),
.Y(n_3564)
);

INVxp67_ASAP7_75t_L g3565 ( 
.A(n_3154),
.Y(n_3565)
);

BUFx3_ASAP7_75t_L g3566 ( 
.A(n_3411),
.Y(n_3566)
);

INVx3_ASAP7_75t_L g3567 ( 
.A(n_3306),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3246),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_SL g3569 ( 
.A(n_3256),
.B(n_2794),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3166),
.B(n_2846),
.Y(n_3570)
);

OAI22xp33_ASAP7_75t_L g3571 ( 
.A1(n_3245),
.A2(n_2848),
.B1(n_2906),
.B2(n_2837),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3270),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3095),
.B(n_2847),
.Y(n_3573)
);

BUFx6f_ASAP7_75t_L g3574 ( 
.A(n_3252),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3271),
.Y(n_3575)
);

HB1xp67_ASAP7_75t_L g3576 ( 
.A(n_3339),
.Y(n_3576)
);

NOR2xp33_ASAP7_75t_L g3577 ( 
.A(n_3157),
.B(n_3059),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_L g3578 ( 
.A(n_3143),
.B(n_3059),
.Y(n_3578)
);

NAND2xp33_ASAP7_75t_L g3579 ( 
.A(n_3198),
.B(n_2800),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_SL g3580 ( 
.A(n_3144),
.B(n_2800),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3090),
.B(n_3093),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3253),
.Y(n_3582)
);

INVx4_ASAP7_75t_L g3583 ( 
.A(n_3411),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3195),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3130),
.B(n_1803),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_SL g3586 ( 
.A(n_3189),
.B(n_2800),
.Y(n_3586)
);

NOR2xp33_ASAP7_75t_L g3587 ( 
.A(n_3086),
.B(n_2861),
.Y(n_3587)
);

INVxp67_ASAP7_75t_L g3588 ( 
.A(n_3099),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3261),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3365),
.A2(n_2854),
.B1(n_2858),
.B2(n_2855),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3266),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3279),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_3284),
.Y(n_3593)
);

INVx3_ASAP7_75t_SL g3594 ( 
.A(n_3254),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_SL g3595 ( 
.A(n_3191),
.B(n_2804),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3127),
.B(n_2861),
.Y(n_3596)
);

AOI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3343),
.A2(n_2859),
.B1(n_2868),
.B2(n_2863),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_SL g3598 ( 
.A(n_3194),
.B(n_2804),
.Y(n_3598)
);

INVx3_ASAP7_75t_L g3599 ( 
.A(n_3341),
.Y(n_3599)
);

CKINVDCx5p33_ASAP7_75t_R g3600 ( 
.A(n_3310),
.Y(n_3600)
);

INVx4_ASAP7_75t_L g3601 ( 
.A(n_3411),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3283),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_3147),
.B(n_3178),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3090),
.B(n_3060),
.Y(n_3604)
);

BUFx2_ASAP7_75t_L g3605 ( 
.A(n_3417),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3319),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3292),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3216),
.B(n_3003),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3293),
.Y(n_3609)
);

BUFx6f_ASAP7_75t_L g3610 ( 
.A(n_3252),
.Y(n_3610)
);

NOR2xp33_ASAP7_75t_L g3611 ( 
.A(n_3327),
.B(n_2861),
.Y(n_3611)
);

AND2x4_ASAP7_75t_L g3612 ( 
.A(n_3259),
.B(n_2862),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3332),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3181),
.B(n_3007),
.Y(n_3614)
);

INVx3_ASAP7_75t_L g3615 ( 
.A(n_3341),
.Y(n_3615)
);

CKINVDCx5p33_ASAP7_75t_R g3616 ( 
.A(n_3168),
.Y(n_3616)
);

INVxp67_ASAP7_75t_SL g3617 ( 
.A(n_3433),
.Y(n_3617)
);

INVx2_ASAP7_75t_SL g3618 ( 
.A(n_3173),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3302),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3312),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3317),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3322),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3334),
.Y(n_3623)
);

CKINVDCx5p33_ASAP7_75t_R g3624 ( 
.A(n_3126),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3249),
.B(n_2804),
.Y(n_3625)
);

INVx2_ASAP7_75t_SL g3626 ( 
.A(n_3421),
.Y(n_3626)
);

BUFx3_ASAP7_75t_L g3627 ( 
.A(n_3291),
.Y(n_3627)
);

BUFx6f_ASAP7_75t_L g3628 ( 
.A(n_3291),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3336),
.Y(n_3629)
);

CKINVDCx5p33_ASAP7_75t_R g3630 ( 
.A(n_3298),
.Y(n_3630)
);

CKINVDCx5p33_ASAP7_75t_R g3631 ( 
.A(n_3225),
.Y(n_3631)
);

INVx1_ASAP7_75t_SL g3632 ( 
.A(n_3101),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_3335),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3342),
.Y(n_3634)
);

AO22x1_ASAP7_75t_L g3635 ( 
.A1(n_3288),
.A2(n_3289),
.B1(n_3297),
.B2(n_3326),
.Y(n_3635)
);

BUFx4f_ASAP7_75t_L g3636 ( 
.A(n_3243),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_SL g3637 ( 
.A(n_3272),
.B(n_2809),
.Y(n_3637)
);

NAND2x1p5_ASAP7_75t_L g3638 ( 
.A(n_3175),
.B(n_2809),
.Y(n_3638)
);

AOI22xp5_ASAP7_75t_SL g3639 ( 
.A1(n_3300),
.A2(n_1099),
.B1(n_1100),
.B2(n_1096),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3093),
.B(n_3073),
.Y(n_3640)
);

AOI22xp33_ASAP7_75t_L g3641 ( 
.A1(n_3107),
.A2(n_2875),
.B1(n_2809),
.B2(n_2817),
.Y(n_3641)
);

INVx4_ASAP7_75t_L g3642 ( 
.A(n_3291),
.Y(n_3642)
);

INVxp67_ASAP7_75t_L g3643 ( 
.A(n_3340),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3345),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_3307),
.B(n_2862),
.Y(n_3645)
);

INVx2_ASAP7_75t_SL g3646 ( 
.A(n_3428),
.Y(n_3646)
);

NOR2xp33_ASAP7_75t_L g3647 ( 
.A(n_3149),
.B(n_2862),
.Y(n_3647)
);

INVx4_ASAP7_75t_L g3648 ( 
.A(n_3331),
.Y(n_3648)
);

AND2x4_ASAP7_75t_L g3649 ( 
.A(n_3333),
.B(n_2813),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_SL g3650 ( 
.A(n_3193),
.B(n_2813),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3360),
.Y(n_3651)
);

CKINVDCx5p33_ASAP7_75t_R g3652 ( 
.A(n_3217),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3145),
.B(n_3009),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3362),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3206),
.B(n_3012),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3087),
.B(n_3046),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3352),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3357),
.Y(n_3658)
);

AND2x4_ASAP7_75t_L g3659 ( 
.A(n_3083),
.B(n_2813),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_SL g3660 ( 
.A(n_3308),
.B(n_2817),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_SL g3661 ( 
.A(n_3308),
.B(n_2817),
.Y(n_3661)
);

AOI22xp5_ASAP7_75t_L g3662 ( 
.A1(n_3186),
.A2(n_2875),
.B1(n_3050),
.B2(n_3027),
.Y(n_3662)
);

NOR2xp67_ASAP7_75t_L g3663 ( 
.A(n_3299),
.B(n_3054),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3278),
.B(n_3065),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3361),
.Y(n_3665)
);

OR2x2_ASAP7_75t_L g3666 ( 
.A(n_3081),
.B(n_3067),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3363),
.B(n_1803),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3418),
.B(n_2935),
.Y(n_3668)
);

CKINVDCx5p33_ASAP7_75t_R g3669 ( 
.A(n_3219),
.Y(n_3669)
);

INVx1_ASAP7_75t_SL g3670 ( 
.A(n_3101),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3323),
.B(n_2826),
.Y(n_3671)
);

HB1xp67_ASAP7_75t_L g3672 ( 
.A(n_3331),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3200),
.B(n_3207),
.Y(n_3673)
);

AOI22xp33_ASAP7_75t_L g3674 ( 
.A1(n_3348),
.A2(n_2875),
.B1(n_2853),
.B2(n_2826),
.Y(n_3674)
);

INVxp67_ASAP7_75t_L g3675 ( 
.A(n_3116),
.Y(n_3675)
);

AND2x4_ASAP7_75t_L g3676 ( 
.A(n_3151),
.B(n_2826),
.Y(n_3676)
);

INVxp67_ASAP7_75t_SL g3677 ( 
.A(n_3367),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3371),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3286),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_SL g3680 ( 
.A(n_3359),
.B(n_2853),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3171),
.Y(n_3681)
);

BUFx6f_ASAP7_75t_L g3682 ( 
.A(n_3331),
.Y(n_3682)
);

NAND2x1p5_ASAP7_75t_L g3683 ( 
.A(n_3175),
.B(n_2853),
.Y(n_3683)
);

BUFx3_ASAP7_75t_L g3684 ( 
.A(n_3347),
.Y(n_3684)
);

AOI22xp5_ASAP7_75t_L g3685 ( 
.A1(n_3265),
.A2(n_2875),
.B1(n_1851),
.B2(n_925),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3384),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3414),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3171),
.Y(n_3688)
);

AND2x4_ASAP7_75t_L g3689 ( 
.A(n_3167),
.B(n_3057),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3290),
.B(n_2933),
.Y(n_3690)
);

BUFx2_ASAP7_75t_SL g3691 ( 
.A(n_3407),
.Y(n_3691)
);

INVx1_ASAP7_75t_SL g3692 ( 
.A(n_3108),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3211),
.B(n_3011),
.Y(n_3693)
);

INVx5_ASAP7_75t_L g3694 ( 
.A(n_3347),
.Y(n_3694)
);

AOI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3113),
.A2(n_1851),
.B1(n_938),
.B2(n_940),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3087),
.B(n_2981),
.Y(n_3696)
);

BUFx6f_ASAP7_75t_L g3697 ( 
.A(n_3347),
.Y(n_3697)
);

INVx3_ASAP7_75t_L g3698 ( 
.A(n_3462),
.Y(n_3698)
);

HB1xp67_ASAP7_75t_L g3699 ( 
.A(n_3453),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3657),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_SL g3701 ( 
.A(n_3554),
.B(n_3177),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3665),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3471),
.B(n_3170),
.Y(n_3703)
);

OAI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3464),
.A2(n_3113),
.B1(n_3321),
.B2(n_3114),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3469),
.Y(n_3705)
);

O2A1O1Ixp5_ASAP7_75t_SL g3706 ( 
.A1(n_3650),
.A2(n_3440),
.B(n_1099),
.C(n_1107),
.Y(n_3706)
);

O2A1O1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_3643),
.A2(n_3146),
.B(n_3205),
.C(n_3190),
.Y(n_3707)
);

O2A1O1Ixp33_ASAP7_75t_L g3708 ( 
.A1(n_3547),
.A2(n_3204),
.B(n_3405),
.C(n_3239),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3678),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_L g3710 ( 
.A(n_3453),
.Y(n_3710)
);

NOR2x1_ASAP7_75t_L g3711 ( 
.A(n_3461),
.B(n_3315),
.Y(n_3711)
);

NOR2xp33_ASAP7_75t_L g3712 ( 
.A(n_3563),
.B(n_3394),
.Y(n_3712)
);

AOI22xp33_ASAP7_75t_L g3713 ( 
.A1(n_3553),
.A2(n_3356),
.B1(n_3197),
.B2(n_3212),
.Y(n_3713)
);

BUFx2_ASAP7_75t_L g3714 ( 
.A(n_3445),
.Y(n_3714)
);

NOR2xp33_ASAP7_75t_L g3715 ( 
.A(n_3565),
.B(n_3436),
.Y(n_3715)
);

AOI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_3579),
.A2(n_3187),
.B(n_3109),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3441),
.B(n_3427),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3631),
.B(n_3438),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3468),
.A2(n_3158),
.B(n_3233),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3468),
.A2(n_3439),
.B(n_3208),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3476),
.Y(n_3721)
);

NOR2xp33_ASAP7_75t_L g3722 ( 
.A(n_3577),
.B(n_3199),
.Y(n_3722)
);

BUFx6f_ASAP7_75t_L g3723 ( 
.A(n_3467),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_SL g3724 ( 
.A(n_3442),
.B(n_3435),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3531),
.A2(n_3355),
.B(n_3152),
.Y(n_3725)
);

INVx4_ASAP7_75t_SL g3726 ( 
.A(n_3484),
.Y(n_3726)
);

AOI22xp33_ASAP7_75t_L g3727 ( 
.A1(n_3553),
.A2(n_3235),
.B1(n_3244),
.B2(n_3236),
.Y(n_3727)
);

OR2x6_ASAP7_75t_L g3728 ( 
.A(n_3484),
.B(n_2933),
.Y(n_3728)
);

BUFx6f_ASAP7_75t_L g3729 ( 
.A(n_3467),
.Y(n_3729)
);

BUFx2_ASAP7_75t_L g3730 ( 
.A(n_3516),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3584),
.B(n_3311),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3447),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3531),
.A2(n_3617),
.B(n_3673),
.Y(n_3733)
);

AOI22xp5_ASAP7_75t_L g3734 ( 
.A1(n_3578),
.A2(n_3505),
.B1(n_3533),
.B2(n_3526),
.Y(n_3734)
);

BUFx12f_ASAP7_75t_L g3735 ( 
.A(n_3477),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3501),
.B(n_3213),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3679),
.B(n_3213),
.Y(n_3737)
);

BUFx6f_ASAP7_75t_L g3738 ( 
.A(n_3528),
.Y(n_3738)
);

AOI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_3534),
.A2(n_3094),
.B(n_3110),
.Y(n_3739)
);

HB1xp67_ASAP7_75t_L g3740 ( 
.A(n_3494),
.Y(n_3740)
);

HB1xp67_ASAP7_75t_L g3741 ( 
.A(n_3481),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3478),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3681),
.B(n_3218),
.Y(n_3743)
);

NOR2xp67_ASAP7_75t_L g3744 ( 
.A(n_3473),
.B(n_3315),
.Y(n_3744)
);

AO21x1_ASAP7_75t_L g3745 ( 
.A1(n_3492),
.A2(n_3374),
.B(n_3364),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3457),
.Y(n_3746)
);

AOI22xp33_ASAP7_75t_L g3747 ( 
.A1(n_3496),
.A2(n_3134),
.B1(n_3128),
.B2(n_3124),
.Y(n_3747)
);

OAI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_3636),
.A2(n_3495),
.B1(n_3677),
.B2(n_3675),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3491),
.Y(n_3749)
);

NAND2x1p5_ASAP7_75t_L g3750 ( 
.A(n_3528),
.B(n_3337),
.Y(n_3750)
);

OR2x6_ASAP7_75t_SL g3751 ( 
.A(n_3616),
.B(n_933),
.Y(n_3751)
);

AND2x4_ASAP7_75t_L g3752 ( 
.A(n_3538),
.B(n_3250),
.Y(n_3752)
);

INVx5_ASAP7_75t_L g3753 ( 
.A(n_3528),
.Y(n_3753)
);

OAI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3636),
.A2(n_3353),
.B1(n_3386),
.B2(n_3419),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3688),
.B(n_3218),
.Y(n_3755)
);

BUFx6f_ASAP7_75t_L g3756 ( 
.A(n_3694),
.Y(n_3756)
);

AOI21xp5_ASAP7_75t_L g3757 ( 
.A1(n_3534),
.A2(n_3094),
.B(n_3136),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_SL g3758 ( 
.A(n_3459),
.B(n_3139),
.Y(n_3758)
);

AND2x2_ASAP7_75t_SL g3759 ( 
.A(n_3685),
.B(n_3423),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3495),
.B(n_3220),
.Y(n_3760)
);

HB1xp67_ASAP7_75t_L g3761 ( 
.A(n_3576),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_3475),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_L g3763 ( 
.A(n_3512),
.B(n_3176),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3493),
.Y(n_3764)
);

HB1xp67_ASAP7_75t_L g3765 ( 
.A(n_3466),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3585),
.B(n_3581),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3472),
.B(n_3176),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_3652),
.B(n_3669),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3502),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3535),
.A2(n_3391),
.B(n_3309),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3482),
.Y(n_3771)
);

NOR2xp33_ASAP7_75t_SL g3772 ( 
.A(n_3479),
.B(n_3337),
.Y(n_3772)
);

A2O1A1Ixp33_ASAP7_75t_L g3773 ( 
.A1(n_3490),
.A2(n_3224),
.B(n_3242),
.C(n_3142),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3487),
.Y(n_3774)
);

AOI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3505),
.A2(n_3263),
.B1(n_3255),
.B2(n_3423),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3581),
.B(n_3220),
.Y(n_3776)
);

AOI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_3535),
.A2(n_3330),
.B(n_3303),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3549),
.A2(n_3372),
.B(n_3380),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3549),
.A2(n_3422),
.B(n_3385),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3499),
.Y(n_3780)
);

AOI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3533),
.A2(n_3630),
.B1(n_3690),
.B2(n_3556),
.Y(n_3781)
);

AND2x4_ASAP7_75t_L g3782 ( 
.A(n_3538),
.B(n_3583),
.Y(n_3782)
);

AOI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3443),
.A2(n_3426),
.B1(n_3277),
.B2(n_3325),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_3558),
.A2(n_3570),
.B(n_3656),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3551),
.B(n_3221),
.Y(n_3785)
);

INVx3_ASAP7_75t_L g3786 ( 
.A(n_3462),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_3558),
.A2(n_3415),
.B(n_3112),
.Y(n_3787)
);

BUFx2_ASAP7_75t_L g3788 ( 
.A(n_3550),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_SL g3789 ( 
.A(n_3510),
.B(n_3221),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_3588),
.B(n_3268),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_SL g3791 ( 
.A(n_3488),
.B(n_3222),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3503),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3570),
.A2(n_3112),
.B(n_3108),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3497),
.B(n_3222),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3656),
.A2(n_3406),
.B(n_3226),
.Y(n_3795)
);

AOI22x1_ASAP7_75t_L g3796 ( 
.A1(n_3639),
.A2(n_3301),
.B1(n_3163),
.B2(n_3277),
.Y(n_3796)
);

INVx5_ASAP7_75t_L g3797 ( 
.A(n_3694),
.Y(n_3797)
);

INVxp67_ASAP7_75t_SL g3798 ( 
.A(n_3446),
.Y(n_3798)
);

AND2x2_ASAP7_75t_SL g3799 ( 
.A(n_3685),
.B(n_3064),
.Y(n_3799)
);

AOI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3490),
.A2(n_1110),
.B1(n_1051),
.B2(n_3287),
.Y(n_3800)
);

NOR2xp33_ASAP7_75t_L g3801 ( 
.A(n_3470),
.B(n_3268),
.Y(n_3801)
);

OA22x2_ASAP7_75t_L g3802 ( 
.A1(n_3605),
.A2(n_934),
.B1(n_936),
.B2(n_935),
.Y(n_3802)
);

BUFx2_ASAP7_75t_L g3803 ( 
.A(n_3463),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3562),
.B(n_3325),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3545),
.B(n_3223),
.Y(n_3805)
);

OAI22xp5_ASAP7_75t_L g3806 ( 
.A1(n_3641),
.A2(n_3590),
.B1(n_3489),
.B2(n_3544),
.Y(n_3806)
);

AOI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3696),
.A2(n_3226),
.B(n_3223),
.Y(n_3807)
);

BUFx2_ASAP7_75t_L g3808 ( 
.A(n_3672),
.Y(n_3808)
);

AOI21xp5_ASAP7_75t_L g3809 ( 
.A1(n_3696),
.A2(n_3227),
.B(n_3251),
.Y(n_3809)
);

BUFx6f_ASAP7_75t_L g3810 ( 
.A(n_3694),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3626),
.B(n_3368),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_SL g3812 ( 
.A(n_3587),
.B(n_3227),
.Y(n_3812)
);

A2O1A1Ixp33_ASAP7_75t_L g3813 ( 
.A1(n_3639),
.A2(n_3273),
.B(n_3264),
.C(n_3379),
.Y(n_3813)
);

A2O1A1Ixp33_ASAP7_75t_L g3814 ( 
.A1(n_3695),
.A2(n_3041),
.B(n_3368),
.C(n_3389),
.Y(n_3814)
);

O2A1O1Ixp33_ASAP7_75t_L g3815 ( 
.A1(n_3637),
.A2(n_1103),
.B(n_1108),
.C(n_1107),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3603),
.A2(n_3544),
.B(n_3454),
.Y(n_3816)
);

AOI22xp33_ASAP7_75t_L g3817 ( 
.A1(n_3667),
.A2(n_1051),
.B1(n_1110),
.B2(n_3313),
.Y(n_3817)
);

A2O1A1Ixp33_ASAP7_75t_L g3818 ( 
.A1(n_3695),
.A2(n_3294),
.B(n_3320),
.C(n_3358),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3509),
.Y(n_3819)
);

A2O1A1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_3518),
.A2(n_3281),
.B(n_3285),
.C(n_3280),
.Y(n_3820)
);

OAI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_3590),
.A2(n_3295),
.B1(n_3305),
.B2(n_3163),
.Y(n_3821)
);

INVx4_ASAP7_75t_L g3822 ( 
.A(n_3458),
.Y(n_3822)
);

BUFx2_ASAP7_75t_L g3823 ( 
.A(n_3627),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3520),
.B(n_1404),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3632),
.B(n_3251),
.Y(n_3825)
);

AOI21xp5_ASAP7_75t_L g3826 ( 
.A1(n_3454),
.A2(n_3260),
.B(n_3257),
.Y(n_3826)
);

AOI21xp5_ASAP7_75t_L g3827 ( 
.A1(n_3653),
.A2(n_3260),
.B(n_3257),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3646),
.A2(n_3064),
.B1(n_2867),
.B2(n_3387),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3573),
.A2(n_3269),
.B(n_3267),
.Y(n_3829)
);

NAND2x1p5_ASAP7_75t_L g3830 ( 
.A(n_3583),
.B(n_2946),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3632),
.B(n_3267),
.Y(n_3831)
);

AOI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_3573),
.A2(n_3274),
.B(n_3269),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3517),
.Y(n_3833)
);

A2O1A1Ixp33_ASAP7_75t_SL g3834 ( 
.A1(n_3596),
.A2(n_3011),
.B(n_3016),
.C(n_2981),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3523),
.Y(n_3835)
);

BUFx12f_ASAP7_75t_L g3836 ( 
.A(n_3448),
.Y(n_3836)
);

BUFx6f_ASAP7_75t_L g3837 ( 
.A(n_3458),
.Y(n_3837)
);

AND2x2_ASAP7_75t_L g3838 ( 
.A(n_3520),
.B(n_1405),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3670),
.B(n_3274),
.Y(n_3839)
);

BUFx6f_ASAP7_75t_L g3840 ( 
.A(n_3458),
.Y(n_3840)
);

BUFx6f_ASAP7_75t_L g3841 ( 
.A(n_3474),
.Y(n_3841)
);

BUFx6f_ASAP7_75t_L g3842 ( 
.A(n_3474),
.Y(n_3842)
);

AOI21xp5_ASAP7_75t_L g3843 ( 
.A1(n_3693),
.A2(n_3276),
.B(n_3275),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3670),
.B(n_3692),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3663),
.A2(n_3276),
.B(n_3275),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3692),
.B(n_3328),
.Y(n_3846)
);

BUFx6f_ASAP7_75t_L g3847 ( 
.A(n_3474),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_SL g3848 ( 
.A(n_3540),
.B(n_3328),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3663),
.A2(n_3399),
.B(n_3396),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3542),
.Y(n_3850)
);

A2O1A1Ixp33_ASAP7_75t_L g3851 ( 
.A1(n_3662),
.A2(n_3395),
.B(n_3392),
.C(n_3338),
.Y(n_3851)
);

BUFx3_ASAP7_75t_L g3852 ( 
.A(n_3451),
.Y(n_3852)
);

O2A1O1Ixp33_ASAP7_75t_L g3853 ( 
.A1(n_3480),
.A2(n_3625),
.B(n_3569),
.C(n_3555),
.Y(n_3853)
);

A2O1A1Ixp33_ASAP7_75t_L g3854 ( 
.A1(n_3662),
.A2(n_3395),
.B(n_3392),
.C(n_3344),
.Y(n_3854)
);

OAI22xp5_ASAP7_75t_L g3855 ( 
.A1(n_3674),
.A2(n_2887),
.B1(n_2843),
.B2(n_3301),
.Y(n_3855)
);

NOR2xp33_ASAP7_75t_R g3856 ( 
.A(n_3624),
.B(n_2929),
.Y(n_3856)
);

NOR2xp33_ASAP7_75t_L g3857 ( 
.A(n_3567),
.B(n_882),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3614),
.B(n_3369),
.Y(n_3858)
);

A2O1A1Ixp33_ASAP7_75t_L g3859 ( 
.A1(n_3647),
.A2(n_3346),
.B(n_3349),
.C(n_3324),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3543),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3640),
.B(n_3373),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_SL g3862 ( 
.A(n_3659),
.B(n_3366),
.Y(n_3862)
);

AOI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3580),
.A2(n_1110),
.B1(n_1051),
.B2(n_2774),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3504),
.Y(n_3864)
);

AOI21xp5_ASAP7_75t_L g3865 ( 
.A1(n_3604),
.A2(n_3399),
.B(n_3396),
.Y(n_3865)
);

INVx5_ASAP7_75t_L g3866 ( 
.A(n_3483),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3640),
.B(n_3376),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3604),
.A2(n_3402),
.B(n_3400),
.Y(n_3868)
);

NOR2xp33_ASAP7_75t_L g3869 ( 
.A(n_3567),
.B(n_3635),
.Y(n_3869)
);

NOR2xp33_ASAP7_75t_L g3870 ( 
.A(n_3536),
.B(n_941),
.Y(n_3870)
);

NOR2xp33_ASAP7_75t_L g3871 ( 
.A(n_3536),
.B(n_942),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3552),
.Y(n_3872)
);

O2A1O1Ixp33_ASAP7_75t_L g3873 ( 
.A1(n_3680),
.A2(n_3571),
.B(n_3595),
.C(n_3586),
.Y(n_3873)
);

OAI22xp5_ASAP7_75t_L g3874 ( 
.A1(n_3597),
.A2(n_3354),
.B1(n_3350),
.B2(n_2986),
.Y(n_3874)
);

OAI22xp5_ASAP7_75t_SL g3875 ( 
.A1(n_3524),
.A2(n_939),
.B1(n_947),
.B2(n_937),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3686),
.B(n_3377),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3687),
.B(n_3378),
.Y(n_3877)
);

OR2x2_ASAP7_75t_L g3878 ( 
.A(n_3557),
.B(n_3403),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3655),
.A2(n_3402),
.B(n_3400),
.Y(n_3879)
);

OAI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3597),
.A2(n_2934),
.B1(n_2923),
.B2(n_2924),
.Y(n_3880)
);

BUFx3_ASAP7_75t_L g3881 ( 
.A(n_3522),
.Y(n_3881)
);

NOR3xp33_ASAP7_75t_L g3882 ( 
.A(n_3668),
.B(n_1407),
.C(n_1406),
.Y(n_3882)
);

BUFx6f_ASAP7_75t_L g3883 ( 
.A(n_3483),
.Y(n_3883)
);

OAI21xp33_ASAP7_75t_SL g3884 ( 
.A1(n_3598),
.A2(n_2810),
.B(n_2806),
.Y(n_3884)
);

O2A1O1Ixp33_ASAP7_75t_L g3885 ( 
.A1(n_3664),
.A2(n_3608),
.B(n_3661),
.C(n_3660),
.Y(n_3885)
);

AOI21xp33_ASAP7_75t_L g3886 ( 
.A1(n_3666),
.A2(n_3408),
.B(n_3403),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3659),
.B(n_3381),
.Y(n_3887)
);

BUFx2_ASAP7_75t_L g3888 ( 
.A(n_3684),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3582),
.B(n_3382),
.Y(n_3889)
);

BUFx6f_ASAP7_75t_L g3890 ( 
.A(n_3483),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3676),
.B(n_2929),
.Y(n_3891)
);

AOI21xp5_ASAP7_75t_L g3892 ( 
.A1(n_3671),
.A2(n_2525),
.B(n_2470),
.Y(n_3892)
);

A2O1A1Ixp33_ASAP7_75t_L g3893 ( 
.A1(n_3611),
.A2(n_3425),
.B(n_3430),
.C(n_3424),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3689),
.A2(n_2525),
.B(n_2470),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3689),
.A2(n_2525),
.B(n_2586),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3507),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3511),
.A2(n_2978),
.B(n_3375),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3589),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_3599),
.B(n_944),
.Y(n_3899)
);

AOI22xp5_ASAP7_75t_L g3900 ( 
.A1(n_3618),
.A2(n_967),
.B1(n_974),
.B2(n_961),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3513),
.A2(n_2978),
.B(n_3424),
.Y(n_3901)
);

OAI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3444),
.A2(n_2923),
.B1(n_2924),
.B2(n_2921),
.Y(n_3902)
);

O2A1O1Ixp33_ASAP7_75t_L g3903 ( 
.A1(n_3449),
.A2(n_1108),
.B(n_1109),
.C(n_1103),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3515),
.A2(n_3430),
.B(n_3425),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3521),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3591),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3593),
.B(n_3408),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3606),
.B(n_1408),
.Y(n_3908)
);

A2O1A1Ixp33_ASAP7_75t_L g3909 ( 
.A1(n_3452),
.A2(n_3432),
.B(n_3416),
.C(n_3409),
.Y(n_3909)
);

NAND3xp33_ASAP7_75t_L g3910 ( 
.A(n_3448),
.B(n_949),
.C(n_948),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3613),
.Y(n_3911)
);

OAI21x1_ASAP7_75t_L g3912 ( 
.A1(n_3537),
.A2(n_3432),
.B(n_3416),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3525),
.A2(n_3048),
.B(n_2524),
.Y(n_3913)
);

AOI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3612),
.A2(n_982),
.B1(n_987),
.B2(n_976),
.Y(n_3914)
);

OAI21x1_ASAP7_75t_SL g3915 ( 
.A1(n_3532),
.A2(n_3409),
.B(n_2940),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3633),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3539),
.A2(n_2524),
.B(n_3397),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3634),
.B(n_3654),
.Y(n_3918)
);

CKINVDCx14_ASAP7_75t_R g3919 ( 
.A(n_3450),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3651),
.B(n_3599),
.Y(n_3920)
);

NOR3xp33_ASAP7_75t_L g3921 ( 
.A(n_3615),
.B(n_1412),
.C(n_1410),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3541),
.A2(n_2524),
.B(n_3397),
.Y(n_3922)
);

AND2x4_ASAP7_75t_L g3923 ( 
.A(n_3601),
.B(n_2929),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3546),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3456),
.B(n_3460),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3548),
.A2(n_2940),
.B(n_2921),
.Y(n_3926)
);

NOR3xp33_ASAP7_75t_SL g3927 ( 
.A(n_3519),
.B(n_953),
.C(n_952),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3465),
.B(n_1848),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3615),
.B(n_1414),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_3676),
.B(n_2949),
.Y(n_3930)
);

NAND3xp33_ASAP7_75t_SL g3931 ( 
.A(n_3600),
.B(n_956),
.C(n_954),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3559),
.B(n_1848),
.Y(n_3932)
);

AOI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3701),
.A2(n_3612),
.B1(n_3455),
.B2(n_3594),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3705),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3721),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3766),
.B(n_3644),
.Y(n_3936)
);

CKINVDCx20_ASAP7_75t_R g3937 ( 
.A(n_3919),
.Y(n_3937)
);

INVx4_ASAP7_75t_L g3938 ( 
.A(n_3738),
.Y(n_3938)
);

INVx2_ASAP7_75t_SL g3939 ( 
.A(n_3852),
.Y(n_3939)
);

CKINVDCx5p33_ASAP7_75t_R g3940 ( 
.A(n_3735),
.Y(n_3940)
);

AOI22xp33_ASAP7_75t_L g3941 ( 
.A1(n_3759),
.A2(n_3527),
.B1(n_3649),
.B2(n_3645),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3742),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3749),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3764),
.Y(n_3944)
);

BUFx6f_ASAP7_75t_L g3945 ( 
.A(n_3881),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3844),
.Y(n_3946)
);

INVxp67_ASAP7_75t_SL g3947 ( 
.A(n_3765),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3731),
.B(n_3658),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3700),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3769),
.Y(n_3950)
);

BUFx6f_ASAP7_75t_L g3951 ( 
.A(n_3738),
.Y(n_3951)
);

BUFx2_ASAP7_75t_L g3952 ( 
.A(n_3798),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3702),
.Y(n_3953)
);

INVx5_ASAP7_75t_L g3954 ( 
.A(n_3753),
.Y(n_3954)
);

INVx5_ASAP7_75t_L g3955 ( 
.A(n_3753),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3733),
.A2(n_3561),
.B(n_3560),
.Y(n_3956)
);

A2O1A1Ixp33_ASAP7_75t_L g3957 ( 
.A1(n_3708),
.A2(n_3498),
.B(n_3508),
.C(n_3568),
.Y(n_3957)
);

AND2x4_ASAP7_75t_L g3958 ( 
.A(n_3767),
.B(n_3601),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3709),
.Y(n_3959)
);

AOI221xp5_ASAP7_75t_L g3960 ( 
.A1(n_3903),
.A2(n_965),
.B1(n_968),
.B2(n_963),
.C(n_959),
.Y(n_3960)
);

AOI221xp5_ASAP7_75t_L g3961 ( 
.A1(n_3800),
.A2(n_3703),
.B1(n_3815),
.B2(n_3882),
.C(n_3720),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3864),
.Y(n_3962)
);

AOI22xp33_ASAP7_75t_L g3963 ( 
.A1(n_3869),
.A2(n_3649),
.B1(n_3645),
.B2(n_3486),
.Y(n_3963)
);

INVx1_ASAP7_75t_SL g3964 ( 
.A(n_3714),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3896),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3905),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3734),
.A2(n_3530),
.B1(n_3566),
.B2(n_3691),
.Y(n_3967)
);

HB1xp67_ASAP7_75t_L g3968 ( 
.A(n_3699),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3924),
.Y(n_3969)
);

BUFx4_ASAP7_75t_SL g3970 ( 
.A(n_3728),
.Y(n_3970)
);

INVxp67_ASAP7_75t_L g3971 ( 
.A(n_3710),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3732),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3925),
.Y(n_3973)
);

AOI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3848),
.A2(n_3486),
.B1(n_1114),
.B2(n_1115),
.Y(n_3974)
);

AOI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3784),
.A2(n_3575),
.B(n_3572),
.Y(n_3975)
);

INVx3_ASAP7_75t_L g3976 ( 
.A(n_3723),
.Y(n_3976)
);

A2O1A1Ixp33_ASAP7_75t_L g3977 ( 
.A1(n_3707),
.A2(n_3602),
.B(n_3607),
.C(n_3592),
.Y(n_3977)
);

INVx2_ASAP7_75t_SL g3978 ( 
.A(n_3803),
.Y(n_3978)
);

INVx3_ASAP7_75t_L g3979 ( 
.A(n_3723),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3760),
.B(n_3609),
.Y(n_3980)
);

A2O1A1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3716),
.A2(n_3620),
.B(n_3621),
.C(n_3619),
.Y(n_3981)
);

OR2x6_ASAP7_75t_L g3982 ( 
.A(n_3723),
.B(n_3638),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3746),
.Y(n_3983)
);

BUFx6f_ASAP7_75t_L g3984 ( 
.A(n_3729),
.Y(n_3984)
);

BUFx6f_ASAP7_75t_L g3985 ( 
.A(n_3729),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3762),
.Y(n_3986)
);

AOI221xp5_ASAP7_75t_L g3987 ( 
.A1(n_3875),
.A2(n_971),
.B1(n_973),
.B2(n_970),
.C(n_969),
.Y(n_3987)
);

OR2x6_ASAP7_75t_L g3988 ( 
.A(n_3729),
.B(n_3744),
.Y(n_3988)
);

BUFx2_ASAP7_75t_L g3989 ( 
.A(n_3740),
.Y(n_3989)
);

BUFx3_ASAP7_75t_L g3990 ( 
.A(n_3823),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3771),
.Y(n_3991)
);

BUFx6f_ASAP7_75t_L g3992 ( 
.A(n_3738),
.Y(n_3992)
);

BUFx12f_ASAP7_75t_L g3993 ( 
.A(n_3836),
.Y(n_3993)
);

INVx1_ASAP7_75t_SL g3994 ( 
.A(n_3718),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3736),
.B(n_3623),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3774),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3717),
.B(n_3622),
.Y(n_3997)
);

BUFx4f_ASAP7_75t_L g3998 ( 
.A(n_3756),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3737),
.B(n_3629),
.Y(n_3999)
);

BUFx3_ASAP7_75t_L g4000 ( 
.A(n_3888),
.Y(n_4000)
);

OR2x2_ASAP7_75t_SL g4001 ( 
.A(n_3931),
.B(n_1109),
.Y(n_4001)
);

BUFx3_ASAP7_75t_L g4002 ( 
.A(n_3728),
.Y(n_4002)
);

OR2x2_ASAP7_75t_L g4003 ( 
.A(n_3761),
.B(n_3485),
.Y(n_4003)
);

OR2x2_ASAP7_75t_L g4004 ( 
.A(n_3748),
.B(n_3500),
.Y(n_4004)
);

BUFx2_ASAP7_75t_L g4005 ( 
.A(n_3884),
.Y(n_4005)
);

BUFx2_ASAP7_75t_L g4006 ( 
.A(n_3808),
.Y(n_4006)
);

AOI21xp5_ASAP7_75t_L g4007 ( 
.A1(n_3816),
.A2(n_2999),
.B(n_2946),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3920),
.B(n_3506),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3780),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3789),
.B(n_3506),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3722),
.B(n_3506),
.Y(n_4011)
);

AOI22xp5_ASAP7_75t_L g4012 ( 
.A1(n_3712),
.A2(n_3514),
.B1(n_980),
.B2(n_983),
.Y(n_4012)
);

BUFx4f_ASAP7_75t_L g4013 ( 
.A(n_3756),
.Y(n_4013)
);

INVx1_ASAP7_75t_SL g4014 ( 
.A(n_3730),
.Y(n_4014)
);

NOR2x1_ASAP7_75t_SL g4015 ( 
.A(n_3753),
.B(n_3529),
.Y(n_4015)
);

BUFx6f_ASAP7_75t_L g4016 ( 
.A(n_3756),
.Y(n_4016)
);

BUFx6f_ASAP7_75t_L g4017 ( 
.A(n_3810),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3792),
.Y(n_4018)
);

O2A1O1Ixp33_ASAP7_75t_L g4019 ( 
.A1(n_3724),
.A2(n_1115),
.B(n_1116),
.C(n_1114),
.Y(n_4019)
);

INVx8_ASAP7_75t_L g4020 ( 
.A(n_3797),
.Y(n_4020)
);

OAI21x1_ASAP7_75t_SL g4021 ( 
.A1(n_3915),
.A2(n_3648),
.B(n_3642),
.Y(n_4021)
);

HB1xp67_ASAP7_75t_L g4022 ( 
.A(n_3741),
.Y(n_4022)
);

BUFx2_ASAP7_75t_L g4023 ( 
.A(n_3788),
.Y(n_4023)
);

AOI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3781),
.A2(n_985),
.B1(n_988),
.B2(n_979),
.Y(n_4024)
);

INVx3_ASAP7_75t_L g4025 ( 
.A(n_3822),
.Y(n_4025)
);

OR2x6_ASAP7_75t_L g4026 ( 
.A(n_3782),
.B(n_3638),
.Y(n_4026)
);

NOR2xp67_ASAP7_75t_L g4027 ( 
.A(n_3768),
.B(n_3642),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_SL g4028 ( 
.A(n_3711),
.B(n_3529),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3824),
.B(n_3529),
.Y(n_4029)
);

AOI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3715),
.A2(n_992),
.B1(n_994),
.B2(n_989),
.Y(n_4030)
);

AOI22xp33_ASAP7_75t_L g4031 ( 
.A1(n_3802),
.A2(n_1117),
.B1(n_1118),
.B2(n_1116),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3819),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3776),
.B(n_3564),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_L g4034 ( 
.A1(n_3921),
.A2(n_1118),
.B1(n_1124),
.B2(n_1117),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3833),
.Y(n_4035)
);

INVx3_ASAP7_75t_L g4036 ( 
.A(n_3822),
.Y(n_4036)
);

OAI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3773),
.A2(n_3434),
.B(n_3683),
.Y(n_4037)
);

AOI22xp5_ASAP7_75t_L g4038 ( 
.A1(n_3870),
.A2(n_1001),
.B1(n_1003),
.B2(n_1002),
.Y(n_4038)
);

CKINVDCx11_ASAP7_75t_R g4039 ( 
.A(n_3751),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_3835),
.Y(n_4040)
);

BUFx8_ASAP7_75t_L g4041 ( 
.A(n_3810),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3850),
.Y(n_4042)
);

BUFx4_ASAP7_75t_SL g4043 ( 
.A(n_3910),
.Y(n_4043)
);

AOI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_3826),
.A2(n_3005),
.B(n_2999),
.Y(n_4044)
);

BUFx6f_ASAP7_75t_L g4045 ( 
.A(n_3810),
.Y(n_4045)
);

OAI21x1_ASAP7_75t_L g4046 ( 
.A1(n_3912),
.A2(n_3018),
.B(n_3016),
.Y(n_4046)
);

AOI22xp5_ASAP7_75t_L g4047 ( 
.A1(n_3871),
.A2(n_1009),
.B1(n_1014),
.B2(n_1012),
.Y(n_4047)
);

HB1xp67_ASAP7_75t_L g4048 ( 
.A(n_3825),
.Y(n_4048)
);

CKINVDCx20_ASAP7_75t_R g4049 ( 
.A(n_3856),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_3838),
.B(n_3564),
.Y(n_4050)
);

AOI22xp33_ASAP7_75t_L g4051 ( 
.A1(n_3704),
.A2(n_1418),
.B1(n_1419),
.B2(n_1415),
.Y(n_4051)
);

BUFx2_ASAP7_75t_L g4052 ( 
.A(n_3831),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3860),
.Y(n_4053)
);

INVx2_ASAP7_75t_SL g4054 ( 
.A(n_3837),
.Y(n_4054)
);

BUFx12f_ASAP7_75t_L g4055 ( 
.A(n_3837),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3801),
.B(n_3564),
.Y(n_4056)
);

INVx3_ASAP7_75t_L g4057 ( 
.A(n_3782),
.Y(n_4057)
);

AOI22xp5_ASAP7_75t_L g4058 ( 
.A1(n_3772),
.A2(n_1016),
.B1(n_1021),
.B2(n_1018),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3812),
.B(n_3574),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_L g4060 ( 
.A(n_3763),
.B(n_3574),
.Y(n_4060)
);

CKINVDCx20_ASAP7_75t_R g4061 ( 
.A(n_3726),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3872),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_3752),
.B(n_3648),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3898),
.Y(n_4064)
);

A2O1A1Ixp33_ASAP7_75t_L g4065 ( 
.A1(n_3873),
.A2(n_1421),
.B(n_1422),
.C(n_1420),
.Y(n_4065)
);

OAI22xp33_ASAP7_75t_L g4066 ( 
.A1(n_3775),
.A2(n_3754),
.B1(n_3806),
.B2(n_3914),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3906),
.Y(n_4067)
);

CKINVDCx6p67_ASAP7_75t_R g4068 ( 
.A(n_3797),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_3747),
.A2(n_1025),
.B1(n_1031),
.B2(n_1027),
.Y(n_4069)
);

BUFx6f_ASAP7_75t_L g4070 ( 
.A(n_3837),
.Y(n_4070)
);

BUFx6f_ASAP7_75t_L g4071 ( 
.A(n_3840),
.Y(n_4071)
);

NAND2xp33_ASAP7_75t_L g4072 ( 
.A(n_3727),
.B(n_3574),
.Y(n_4072)
);

AOI22xp33_ASAP7_75t_L g4073 ( 
.A1(n_3713),
.A2(n_1425),
.B1(n_1427),
.B2(n_1424),
.Y(n_4073)
);

OAI22xp5_ASAP7_75t_L g4074 ( 
.A1(n_3817),
.A2(n_3683),
.B1(n_3628),
.B2(n_3682),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3911),
.Y(n_4075)
);

INVx1_ASAP7_75t_SL g4076 ( 
.A(n_3804),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_3794),
.B(n_3610),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3916),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3785),
.B(n_3610),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3918),
.Y(n_4080)
);

A2O1A1Ixp33_ASAP7_75t_L g4081 ( 
.A1(n_3853),
.A2(n_1432),
.B(n_1435),
.C(n_1429),
.Y(n_4081)
);

BUFx3_ASAP7_75t_L g4082 ( 
.A(n_3840),
.Y(n_4082)
);

INVxp67_ASAP7_75t_L g4083 ( 
.A(n_3790),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3929),
.B(n_3908),
.Y(n_4084)
);

AND2x6_ASAP7_75t_L g4085 ( 
.A(n_3752),
.B(n_3610),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3839),
.Y(n_4086)
);

CKINVDCx5p33_ASAP7_75t_R g4087 ( 
.A(n_3726),
.Y(n_4087)
);

INVx1_ASAP7_75t_SL g4088 ( 
.A(n_3840),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3878),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3743),
.B(n_3628),
.Y(n_4090)
);

AND2x4_ASAP7_75t_L g4091 ( 
.A(n_3698),
.B(n_3628),
.Y(n_4091)
);

AND2x4_ASAP7_75t_L g4092 ( 
.A(n_3698),
.B(n_3682),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3846),
.Y(n_4093)
);

OAI22xp33_ASAP7_75t_L g4094 ( 
.A1(n_3783),
.A2(n_1032),
.B1(n_1038),
.B2(n_1036),
.Y(n_4094)
);

AOI21xp5_ASAP7_75t_L g4095 ( 
.A1(n_3739),
.A2(n_3005),
.B(n_2954),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3755),
.B(n_3682),
.Y(n_4096)
);

NAND2x1_ASAP7_75t_L g4097 ( 
.A(n_3770),
.B(n_2949),
.Y(n_4097)
);

BUFx6f_ASAP7_75t_L g4098 ( 
.A(n_3841),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3786),
.Y(n_4099)
);

INVxp67_ASAP7_75t_L g4100 ( 
.A(n_3811),
.Y(n_4100)
);

AOI33xp33_ASAP7_75t_L g4101 ( 
.A1(n_3900),
.A2(n_1444),
.A3(n_1439),
.B1(n_1446),
.B2(n_1440),
.B3(n_1436),
.Y(n_4101)
);

O2A1O1Ixp33_ASAP7_75t_SL g4102 ( 
.A1(n_3758),
.A2(n_1449),
.B(n_1450),
.C(n_1447),
.Y(n_4102)
);

AOI211xp5_ASAP7_75t_L g4103 ( 
.A1(n_3899),
.A2(n_1041),
.B(n_1052),
.C(n_1048),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_3786),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3928),
.Y(n_4105)
);

NOR2xp33_ASAP7_75t_L g4106 ( 
.A(n_3857),
.B(n_3697),
.Y(n_4106)
);

BUFx6f_ASAP7_75t_L g4107 ( 
.A(n_3841),
.Y(n_4107)
);

BUFx6f_ASAP7_75t_L g4108 ( 
.A(n_3841),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_SL g4109 ( 
.A1(n_3799),
.A2(n_3796),
.B1(n_3821),
.B2(n_3828),
.Y(n_4109)
);

INVx8_ASAP7_75t_L g4110 ( 
.A(n_3797),
.Y(n_4110)
);

OR2x6_ASAP7_75t_L g4111 ( 
.A(n_3830),
.B(n_3697),
.Y(n_4111)
);

AOI22xp5_ASAP7_75t_L g4112 ( 
.A1(n_3927),
.A2(n_1043),
.B1(n_1054),
.B2(n_1053),
.Y(n_4112)
);

INVx5_ASAP7_75t_L g4113 ( 
.A(n_3866),
.Y(n_4113)
);

OAI22xp5_ASAP7_75t_L g4114 ( 
.A1(n_3863),
.A2(n_3697),
.B1(n_3061),
.B2(n_3018),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_3932),
.Y(n_4115)
);

BUFx2_ASAP7_75t_SL g4116 ( 
.A(n_3866),
.Y(n_4116)
);

CKINVDCx8_ASAP7_75t_R g4117 ( 
.A(n_3866),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3907),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3887),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3876),
.Y(n_4120)
);

AOI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_3862),
.A2(n_1056),
.B1(n_1063),
.B2(n_1062),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_3877),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3889),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3901),
.Y(n_4124)
);

BUFx6f_ASAP7_75t_L g4125 ( 
.A(n_3842),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_3891),
.B(n_1451),
.Y(n_4126)
);

INVx3_ASAP7_75t_L g4127 ( 
.A(n_3842),
.Y(n_4127)
);

BUFx6f_ASAP7_75t_L g4128 ( 
.A(n_3842),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3793),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3847),
.Y(n_4130)
);

BUFx3_ASAP7_75t_L g4131 ( 
.A(n_3847),
.Y(n_4131)
);

BUFx6f_ASAP7_75t_L g4132 ( 
.A(n_3847),
.Y(n_4132)
);

AOI21x1_ASAP7_75t_L g4133 ( 
.A1(n_3725),
.A2(n_3897),
.B(n_3917),
.Y(n_4133)
);

OR2x2_ASAP7_75t_L g4134 ( 
.A(n_3861),
.B(n_1454),
.Y(n_4134)
);

AND2x4_ASAP7_75t_L g4135 ( 
.A(n_3930),
.B(n_2949),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3885),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3805),
.B(n_1877),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3791),
.Y(n_4138)
);

NAND3xp33_ASAP7_75t_L g4139 ( 
.A(n_3779),
.B(n_3719),
.C(n_3787),
.Y(n_4139)
);

INVx2_ASAP7_75t_SL g4140 ( 
.A(n_3883),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3858),
.B(n_1877),
.Y(n_4141)
);

AOI22xp5_ASAP7_75t_L g4142 ( 
.A1(n_3855),
.A2(n_1070),
.B1(n_1072),
.B2(n_1068),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3867),
.B(n_1078),
.Y(n_4143)
);

AND2x4_ASAP7_75t_L g4144 ( 
.A(n_3923),
.B(n_2954),
.Y(n_4144)
);

CKINVDCx5p33_ASAP7_75t_R g4145 ( 
.A(n_3883),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3909),
.Y(n_4146)
);

INVx3_ASAP7_75t_L g4147 ( 
.A(n_3883),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_3890),
.B(n_1458),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3745),
.Y(n_4149)
);

BUFx4f_ASAP7_75t_SL g4150 ( 
.A(n_3890),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3829),
.A2(n_2962),
.B(n_2954),
.Y(n_4151)
);

OR2x6_ASAP7_75t_L g4152 ( 
.A(n_3750),
.B(n_2962),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3904),
.Y(n_4153)
);

INVx2_ASAP7_75t_L g4154 ( 
.A(n_3890),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3807),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3832),
.B(n_1079),
.Y(n_4156)
);

OR2x6_ASAP7_75t_L g4157 ( 
.A(n_3923),
.B(n_2962),
.Y(n_4157)
);

INVx4_ASAP7_75t_L g4158 ( 
.A(n_3902),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3809),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3865),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_3777),
.B(n_2993),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3868),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3757),
.Y(n_4163)
);

INVx2_ASAP7_75t_SL g4164 ( 
.A(n_3880),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_SL g4165 ( 
.A(n_3886),
.B(n_2993),
.Y(n_4165)
);

INVx2_ASAP7_75t_SL g4166 ( 
.A(n_3945),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_3969),
.Y(n_4167)
);

AO32x2_ASAP7_75t_L g4168 ( 
.A1(n_4164),
.A2(n_3874),
.A3(n_3834),
.B1(n_3892),
.B2(n_3813),
.Y(n_4168)
);

O2A1O1Ixp33_ASAP7_75t_L g4169 ( 
.A1(n_4066),
.A2(n_3814),
.B(n_3893),
.C(n_3818),
.Y(n_4169)
);

O2A1O1Ixp33_ASAP7_75t_SL g4170 ( 
.A1(n_3994),
.A2(n_3859),
.B(n_3851),
.C(n_3854),
.Y(n_4170)
);

OAI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_3933),
.A2(n_3820),
.B1(n_3926),
.B2(n_3778),
.Y(n_4171)
);

AO32x2_ASAP7_75t_L g4172 ( 
.A1(n_4158),
.A2(n_3706),
.A3(n_1744),
.B1(n_3795),
.B2(n_3849),
.Y(n_4172)
);

AOI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_3961),
.A2(n_4072),
.B1(n_4069),
.B2(n_3967),
.Y(n_4173)
);

AOI22xp5_ASAP7_75t_L g4174 ( 
.A1(n_4106),
.A2(n_1083),
.B1(n_1087),
.B2(n_1084),
.Y(n_4174)
);

A2O1A1Ixp33_ASAP7_75t_L g4175 ( 
.A1(n_4103),
.A2(n_3922),
.B(n_3845),
.C(n_3913),
.Y(n_4175)
);

AO32x2_ASAP7_75t_L g4176 ( 
.A1(n_3978),
.A2(n_1744),
.A3(n_3894),
.B1(n_3879),
.B2(n_3843),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3934),
.Y(n_4177)
);

OR2x2_ASAP7_75t_L g4178 ( 
.A(n_3946),
.B(n_3827),
.Y(n_4178)
);

INVx2_ASAP7_75t_SL g4179 ( 
.A(n_3945),
.Y(n_4179)
);

AO31x2_ASAP7_75t_L g4180 ( 
.A1(n_4124),
.A2(n_3895),
.A3(n_1461),
.B(n_1463),
.Y(n_4180)
);

AOI22xp33_ASAP7_75t_L g4181 ( 
.A1(n_4109),
.A2(n_4136),
.B1(n_4084),
.B2(n_4039),
.Y(n_4181)
);

AOI21xp5_ASAP7_75t_L g4182 ( 
.A1(n_4139),
.A2(n_3036),
.B(n_3035),
.Y(n_4182)
);

INVx3_ASAP7_75t_L g4183 ( 
.A(n_4055),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_3935),
.Y(n_4184)
);

OAI21x1_ASAP7_75t_L g4185 ( 
.A1(n_4133),
.A2(n_3061),
.B(n_2220),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3946),
.B(n_1081),
.Y(n_4186)
);

A2O1A1Ixp33_ASAP7_75t_L g4187 ( 
.A1(n_4005),
.A2(n_1097),
.B(n_1098),
.C(n_1095),
.Y(n_4187)
);

A2O1A1Ixp33_ASAP7_75t_L g4188 ( 
.A1(n_4005),
.A2(n_4101),
.B(n_4142),
.C(n_4024),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4048),
.B(n_4052),
.Y(n_4189)
);

NOR2xp33_ASAP7_75t_L g4190 ( 
.A(n_4083),
.B(n_1104),
.Y(n_4190)
);

OAI21x1_ASAP7_75t_L g4191 ( 
.A1(n_4133),
.A2(n_2229),
.B(n_2217),
.Y(n_4191)
);

AOI221x1_ASAP7_75t_L g4192 ( 
.A1(n_4149),
.A2(n_1467),
.B1(n_1468),
.B2(n_1465),
.C(n_1459),
.Y(n_4192)
);

O2A1O1Ixp33_ASAP7_75t_L g4193 ( 
.A1(n_4156),
.A2(n_1469),
.B(n_1476),
.C(n_1475),
.Y(n_4193)
);

OAI21x1_ASAP7_75t_L g4194 ( 
.A1(n_4046),
.A2(n_3956),
.B(n_4097),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_4011),
.B(n_4089),
.Y(n_4195)
);

AOI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_4155),
.A2(n_3035),
.B(n_3025),
.Y(n_4196)
);

NAND2x1p5_ASAP7_75t_L g4197 ( 
.A(n_4113),
.B(n_2993),
.Y(n_4197)
);

OAI21x1_ASAP7_75t_L g4198 ( 
.A1(n_4097),
.A2(n_2237),
.B(n_2236),
.Y(n_4198)
);

AND2x2_ASAP7_75t_L g4199 ( 
.A(n_4008),
.B(n_1478),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3942),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_3943),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_3944),
.Y(n_4202)
);

OAI21x1_ASAP7_75t_L g4203 ( 
.A1(n_3975),
.A2(n_2237),
.B(n_2236),
.Y(n_4203)
);

OAI211xp5_ASAP7_75t_L g4204 ( 
.A1(n_4031),
.A2(n_1106),
.B(n_1480),
.C(n_1479),
.Y(n_4204)
);

OAI21x1_ASAP7_75t_L g4205 ( 
.A1(n_4095),
.A2(n_2254),
.B(n_2246),
.Y(n_4205)
);

CKINVDCx6p67_ASAP7_75t_R g4206 ( 
.A(n_3937),
.Y(n_4206)
);

AO21x2_ASAP7_75t_L g4207 ( 
.A1(n_4161),
.A2(n_1482),
.B(n_1481),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3950),
.Y(n_4208)
);

A2O1A1Ixp33_ASAP7_75t_L g4209 ( 
.A1(n_3974),
.A2(n_1488),
.B(n_1489),
.C(n_1486),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_4159),
.A2(n_3015),
.B(n_2997),
.Y(n_4210)
);

O2A1O1Ixp33_ASAP7_75t_L g4211 ( 
.A1(n_4094),
.A2(n_1494),
.B(n_1496),
.C(n_1491),
.Y(n_4211)
);

OAI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_3957),
.A2(n_1502),
.B(n_1499),
.Y(n_4212)
);

AO31x2_ASAP7_75t_L g4213 ( 
.A1(n_4153),
.A2(n_4163),
.A3(n_4162),
.B(n_4160),
.Y(n_4213)
);

O2A1O1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_4065),
.A2(n_4081),
.B(n_3977),
.C(n_4019),
.Y(n_4214)
);

AOI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_4129),
.A2(n_3036),
.B(n_3035),
.Y(n_4215)
);

OAI21x1_ASAP7_75t_L g4216 ( 
.A1(n_4044),
.A2(n_2254),
.B(n_2246),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_SL g4217 ( 
.A(n_4027),
.B(n_1506),
.Y(n_4217)
);

OAI21xp5_ASAP7_75t_L g4218 ( 
.A1(n_4051),
.A2(n_1508),
.B(n_1507),
.Y(n_4218)
);

BUFx5_ASAP7_75t_L g4219 ( 
.A(n_4146),
.Y(n_4219)
);

A2O1A1Ixp33_ASAP7_75t_L g4220 ( 
.A1(n_4073),
.A2(n_1514),
.B(n_1515),
.C(n_1511),
.Y(n_4220)
);

O2A1O1Ixp33_ASAP7_75t_SL g4221 ( 
.A1(n_4028),
.A2(n_1519),
.B(n_1530),
.C(n_1518),
.Y(n_4221)
);

AOI21xp5_ASAP7_75t_L g4222 ( 
.A1(n_4151),
.A2(n_3015),
.B(n_2997),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_4007),
.A2(n_3015),
.B(n_2997),
.Y(n_4223)
);

AOI21xp5_ASAP7_75t_L g4224 ( 
.A1(n_3954),
.A2(n_3036),
.B(n_3025),
.Y(n_4224)
);

AOI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_3941),
.A2(n_1533),
.B1(n_1541),
.B2(n_1531),
.Y(n_4225)
);

NOR2xp33_ASAP7_75t_L g4226 ( 
.A(n_4100),
.B(n_993),
.Y(n_4226)
);

INVx2_ASAP7_75t_SL g4227 ( 
.A(n_3970),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_3954),
.A2(n_3044),
.B(n_3025),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_L g4229 ( 
.A1(n_4119),
.A2(n_1088),
.B1(n_1101),
.B2(n_1061),
.Y(n_4229)
);

CKINVDCx11_ASAP7_75t_R g4230 ( 
.A(n_3993),
.Y(n_4230)
);

HB1xp67_ASAP7_75t_L g4231 ( 
.A(n_3952),
.Y(n_4231)
);

AOI22xp33_ASAP7_75t_L g4232 ( 
.A1(n_4004),
.A2(n_1105),
.B1(n_1748),
.B2(n_1742),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4052),
.B(n_6),
.Y(n_4233)
);

AOI22xp33_ASAP7_75t_L g4234 ( 
.A1(n_4138),
.A2(n_1748),
.B1(n_1751),
.B2(n_1742),
.Y(n_4234)
);

AO31x2_ASAP7_75t_L g4235 ( 
.A1(n_3981),
.A2(n_2260),
.A3(n_2271),
.B(n_2265),
.Y(n_4235)
);

AOI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_4012),
.A2(n_1661),
.B1(n_1688),
.B2(n_1684),
.Y(n_4236)
);

O2A1O1Ixp33_ASAP7_75t_SL g4237 ( 
.A1(n_4061),
.A2(n_4049),
.B(n_4059),
.C(n_4010),
.Y(n_4237)
);

AOI22xp33_ASAP7_75t_SL g4238 ( 
.A1(n_4037),
.A2(n_2818),
.B1(n_2835),
.B2(n_2774),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_3954),
.A2(n_3044),
.B(n_2687),
.Y(n_4239)
);

AND2x4_ASAP7_75t_L g4240 ( 
.A(n_4023),
.B(n_3044),
.Y(n_4240)
);

O2A1O1Ixp33_ASAP7_75t_L g4241 ( 
.A1(n_4102),
.A2(n_1697),
.B(n_1755),
.C(n_1751),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_3962),
.Y(n_4242)
);

A2O1A1Ixp33_ASAP7_75t_L g4243 ( 
.A1(n_4058),
.A2(n_2265),
.B(n_2271),
.C(n_2260),
.Y(n_4243)
);

AO31x2_ASAP7_75t_L g4244 ( 
.A1(n_4015),
.A2(n_2277),
.A3(n_2283),
.B(n_2281),
.Y(n_4244)
);

OAI21x1_ASAP7_75t_L g4245 ( 
.A1(n_4021),
.A2(n_2283),
.B(n_2281),
.Y(n_4245)
);

OAI222xp33_ASAP7_75t_L g4246 ( 
.A1(n_4076),
.A2(n_1744),
.B1(n_1782),
.B2(n_1790),
.C1(n_1770),
.C2(n_1755),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_4086),
.B(n_1770),
.Y(n_4247)
);

OAI22xp5_ASAP7_75t_L g4248 ( 
.A1(n_3963),
.A2(n_1804),
.B1(n_1782),
.B2(n_1796),
.Y(n_4248)
);

OA21x2_ASAP7_75t_L g4249 ( 
.A1(n_4165),
.A2(n_1796),
.B(n_1790),
.Y(n_4249)
);

OAI22x1_ASAP7_75t_L g4250 ( 
.A1(n_3989),
.A2(n_11),
.B1(n_7),
.B2(n_8),
.Y(n_4250)
);

O2A1O1Ixp33_ASAP7_75t_SL g4251 ( 
.A1(n_3980),
.A2(n_24),
.B(n_32),
.C(n_13),
.Y(n_4251)
);

NOR2x1_ASAP7_75t_R g4252 ( 
.A(n_3940),
.B(n_1730),
.Y(n_4252)
);

BUFx6f_ASAP7_75t_L g4253 ( 
.A(n_3984),
.Y(n_4253)
);

NOR2xp33_ASAP7_75t_L g4254 ( 
.A(n_3964),
.B(n_13),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_3965),
.Y(n_4255)
);

NOR2xp33_ASAP7_75t_L g4256 ( 
.A(n_4014),
.B(n_14),
.Y(n_4256)
);

INVx3_ASAP7_75t_L g4257 ( 
.A(n_3951),
.Y(n_4257)
);

O2A1O1Ixp33_ASAP7_75t_SL g4258 ( 
.A1(n_4143),
.A2(n_25),
.B(n_33),
.C(n_14),
.Y(n_4258)
);

OAI21x1_ASAP7_75t_L g4259 ( 
.A1(n_4021),
.A2(n_1811),
.B(n_1804),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3966),
.Y(n_4260)
);

HB1xp67_ASAP7_75t_SL g4261 ( 
.A(n_4087),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_3949),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_3953),
.Y(n_4263)
);

CKINVDCx20_ASAP7_75t_R g4264 ( 
.A(n_4002),
.Y(n_4264)
);

CKINVDCx20_ASAP7_75t_R g4265 ( 
.A(n_4041),
.Y(n_4265)
);

OAI21x1_ASAP7_75t_L g4266 ( 
.A1(n_4099),
.A2(n_1811),
.B(n_1897),
.Y(n_4266)
);

OAI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_4001),
.A2(n_1793),
.B1(n_1730),
.B2(n_1750),
.Y(n_4267)
);

O2A1O1Ixp33_ASAP7_75t_L g4268 ( 
.A1(n_4074),
.A2(n_1793),
.B(n_2632),
.C(n_18),
.Y(n_4268)
);

A2O1A1Ixp33_ASAP7_75t_L g4269 ( 
.A1(n_4034),
.A2(n_19),
.B(n_15),
.C(n_16),
.Y(n_4269)
);

OAI21x1_ASAP7_75t_L g4270 ( 
.A1(n_4104),
.A2(n_1902),
.B(n_1897),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_3952),
.Y(n_4271)
);

AOI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_3955),
.A2(n_2687),
.B(n_2657),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_3959),
.Y(n_4273)
);

INVx1_ASAP7_75t_SL g4274 ( 
.A(n_3990),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_SL g4275 ( 
.A(n_4117),
.B(n_2774),
.Y(n_4275)
);

OAI22xp33_ASAP7_75t_L g4276 ( 
.A1(n_4134),
.A2(n_1750),
.B1(n_1760),
.B2(n_1745),
.Y(n_4276)
);

NOR2xp33_ASAP7_75t_L g4277 ( 
.A(n_4000),
.B(n_15),
.Y(n_4277)
);

AOI21x1_ASAP7_75t_L g4278 ( 
.A1(n_4137),
.A2(n_2632),
.B(n_1614),
.Y(n_4278)
);

OA21x2_ASAP7_75t_L g4279 ( 
.A1(n_3973),
.A2(n_2818),
.B(n_2774),
.Y(n_4279)
);

AND2x4_ASAP7_75t_L g4280 ( 
.A(n_4023),
.B(n_454),
.Y(n_4280)
);

A2O1A1Ixp33_ASAP7_75t_L g4281 ( 
.A1(n_3987),
.A2(n_22),
.B(n_16),
.C(n_19),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_3955),
.A2(n_2687),
.B(n_1902),
.Y(n_4282)
);

AND2x4_ASAP7_75t_L g4283 ( 
.A(n_4006),
.B(n_455),
.Y(n_4283)
);

AOI21xp5_ASAP7_75t_L g4284 ( 
.A1(n_3955),
.A2(n_1902),
.B(n_1897),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_3947),
.Y(n_4285)
);

OAI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_4056),
.A2(n_1750),
.B1(n_1760),
.B2(n_1745),
.Y(n_4286)
);

OAI22xp5_ASAP7_75t_L g4287 ( 
.A1(n_3971),
.A2(n_1750),
.B1(n_1760),
.B2(n_1745),
.Y(n_4287)
);

OAI21x1_ASAP7_75t_L g4288 ( 
.A1(n_3991),
.A2(n_1944),
.B(n_1918),
.Y(n_4288)
);

AOI22xp33_ASAP7_75t_L g4289 ( 
.A1(n_3989),
.A2(n_2835),
.B1(n_2818),
.B2(n_1760),
.Y(n_4289)
);

OR2x6_ASAP7_75t_L g4290 ( 
.A(n_4020),
.B(n_1745),
.Y(n_4290)
);

A2O1A1Ixp33_ASAP7_75t_L g4291 ( 
.A1(n_4121),
.A2(n_26),
.B(n_23),
.C(n_24),
.Y(n_4291)
);

NOR3xp33_ASAP7_75t_L g4292 ( 
.A(n_3960),
.B(n_1589),
.C(n_1584),
.Y(n_4292)
);

AOI21xp5_ASAP7_75t_L g4293 ( 
.A1(n_3999),
.A2(n_4113),
.B(n_4122),
.Y(n_4293)
);

CKINVDCx11_ASAP7_75t_R g4294 ( 
.A(n_3984),
.Y(n_4294)
);

AOI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_4113),
.A2(n_1944),
.B(n_1918),
.Y(n_4295)
);

OAI21xp5_ASAP7_75t_L g4296 ( 
.A1(n_4038),
.A2(n_2835),
.B(n_2818),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_L g4297 ( 
.A(n_3939),
.B(n_23),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_3968),
.Y(n_4298)
);

OAI22xp33_ASAP7_75t_L g4299 ( 
.A1(n_3988),
.A2(n_1764),
.B1(n_1771),
.B2(n_1763),
.Y(n_4299)
);

OAI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_4047),
.A2(n_2835),
.B(n_3071),
.Y(n_4300)
);

O2A1O1Ixp33_ASAP7_75t_SL g4301 ( 
.A1(n_4090),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_4301)
);

OAI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4030),
.A2(n_3071),
.B(n_2980),
.Y(n_4302)
);

AOI21x1_ASAP7_75t_L g4303 ( 
.A1(n_4141),
.A2(n_1764),
.B(n_1763),
.Y(n_4303)
);

OAI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_4112),
.A2(n_3071),
.B(n_2980),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4022),
.Y(n_4305)
);

AOI21xp5_ASAP7_75t_L g4306 ( 
.A1(n_4120),
.A2(n_1944),
.B(n_1918),
.Y(n_4306)
);

OAI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_4060),
.A2(n_1764),
.B1(n_1771),
.B2(n_1763),
.Y(n_4307)
);

INVx2_ASAP7_75t_SL g4308 ( 
.A(n_4003),
.Y(n_4308)
);

AOI22xp33_ASAP7_75t_L g4309 ( 
.A1(n_4006),
.A2(n_1764),
.B1(n_1771),
.B2(n_1763),
.Y(n_4309)
);

OAI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4105),
.A2(n_3071),
.B(n_2980),
.Y(n_4310)
);

BUFx10_ASAP7_75t_L g4311 ( 
.A(n_3985),
.Y(n_4311)
);

OR2x2_ASAP7_75t_L g4312 ( 
.A(n_4077),
.B(n_1771),
.Y(n_4312)
);

OAI22xp5_ASAP7_75t_L g4313 ( 
.A1(n_4093),
.A2(n_1773),
.B1(n_1792),
.B2(n_1772),
.Y(n_4313)
);

AOI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_3958),
.A2(n_2967),
.B1(n_2980),
.B2(n_1773),
.Y(n_4314)
);

OAI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_4115),
.A2(n_2967),
.B(n_1972),
.Y(n_4315)
);

A2O1A1Ixp33_ASAP7_75t_L g4316 ( 
.A1(n_3998),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_4316)
);

O2A1O1Ixp33_ASAP7_75t_L g4317 ( 
.A1(n_3948),
.A2(n_33),
.B(n_29),
.C(n_32),
.Y(n_4317)
);

NOR2xp67_ASAP7_75t_R g4318 ( 
.A(n_3938),
.B(n_1772),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_3996),
.Y(n_4319)
);

OR2x2_ASAP7_75t_L g4320 ( 
.A(n_3995),
.B(n_1772),
.Y(n_4320)
);

BUFx3_ASAP7_75t_L g4321 ( 
.A(n_4145),
.Y(n_4321)
);

O2A1O1Ixp33_ASAP7_75t_L g4322 ( 
.A1(n_4114),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_4123),
.B(n_35),
.Y(n_4323)
);

OAI21x1_ASAP7_75t_L g4324 ( 
.A1(n_4009),
.A2(n_1972),
.B(n_1970),
.Y(n_4324)
);

BUFx12f_ASAP7_75t_L g4325 ( 
.A(n_4041),
.Y(n_4325)
);

O2A1O1Ixp33_ASAP7_75t_SL g4326 ( 
.A1(n_4096),
.A2(n_4033),
.B(n_3936),
.C(n_4079),
.Y(n_4326)
);

NOR2xp67_ASAP7_75t_L g4327 ( 
.A(n_4018),
.B(n_37),
.Y(n_4327)
);

OAI22xp5_ASAP7_75t_L g4328 ( 
.A1(n_3988),
.A2(n_1773),
.B1(n_1792),
.B2(n_1772),
.Y(n_4328)
);

BUFx3_ASAP7_75t_L g4329 ( 
.A(n_4082),
.Y(n_4329)
);

AO31x2_ASAP7_75t_L g4330 ( 
.A1(n_4032),
.A2(n_1648),
.A3(n_1547),
.B(n_2967),
.Y(n_4330)
);

NOR2xp33_ASAP7_75t_L g4331 ( 
.A(n_4029),
.B(n_37),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_SL g4332 ( 
.A(n_4057),
.B(n_1773),
.Y(n_4332)
);

OAI21x1_ASAP7_75t_L g4333 ( 
.A1(n_4042),
.A2(n_1972),
.B(n_1970),
.Y(n_4333)
);

AOI22xp33_ASAP7_75t_L g4334 ( 
.A1(n_4050),
.A2(n_1794),
.B1(n_1809),
.B2(n_1792),
.Y(n_4334)
);

AND2x6_ASAP7_75t_L g4335 ( 
.A(n_4063),
.B(n_1792),
.Y(n_4335)
);

A2O1A1Ixp33_ASAP7_75t_L g4336 ( 
.A1(n_4013),
.A2(n_41),
.B(n_38),
.C(n_39),
.Y(n_4336)
);

OAI21xp5_ASAP7_75t_L g4337 ( 
.A1(n_4126),
.A2(n_4148),
.B(n_4118),
.Y(n_4337)
);

A2O1A1Ixp33_ASAP7_75t_L g4338 ( 
.A1(n_4020),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_4338)
);

A2O1A1Ixp33_ASAP7_75t_L g4339 ( 
.A1(n_4110),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4080),
.B(n_44),
.Y(n_4340)
);

OR2x6_ASAP7_75t_L g4341 ( 
.A(n_4110),
.B(n_1794),
.Y(n_4341)
);

A2O1A1Ixp33_ASAP7_75t_L g4342 ( 
.A1(n_3997),
.A2(n_51),
.B(n_47),
.C(n_49),
.Y(n_4342)
);

AOI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_4026),
.A2(n_1986),
.B(n_1970),
.Y(n_4343)
);

AO31x2_ASAP7_75t_L g4344 ( 
.A1(n_4053),
.A2(n_1648),
.A3(n_1547),
.B(n_2967),
.Y(n_4344)
);

O2A1O1Ixp33_ASAP7_75t_L g4345 ( 
.A1(n_4062),
.A2(n_53),
.B(n_49),
.C(n_52),
.Y(n_4345)
);

OAI21xp5_ASAP7_75t_L g4346 ( 
.A1(n_4075),
.A2(n_2001),
.B(n_1986),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_3976),
.B(n_54),
.Y(n_4347)
);

BUFx3_ASAP7_75t_L g4348 ( 
.A(n_4131),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4078),
.A2(n_2001),
.B(n_1986),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_3972),
.B(n_54),
.Y(n_4350)
);

O2A1O1Ixp33_ASAP7_75t_SL g4351 ( 
.A1(n_4054),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_4351)
);

OAI22xp33_ASAP7_75t_L g4352 ( 
.A1(n_4068),
.A2(n_1809),
.B1(n_1815),
.B2(n_1794),
.Y(n_4352)
);

OAI21x1_ASAP7_75t_L g4353 ( 
.A1(n_3983),
.A2(n_2010),
.B(n_2001),
.Y(n_4353)
);

AOI21x1_ASAP7_75t_L g4354 ( 
.A1(n_4135),
.A2(n_1809),
.B(n_1794),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_4026),
.A2(n_2041),
.B(n_2010),
.Y(n_4355)
);

AOI21xp5_ASAP7_75t_L g4356 ( 
.A1(n_4111),
.A2(n_2041),
.B(n_2010),
.Y(n_4356)
);

AND2x4_ASAP7_75t_L g4357 ( 
.A(n_3958),
.B(n_456),
.Y(n_4357)
);

CKINVDCx5p33_ASAP7_75t_R g4358 ( 
.A(n_4043),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_3986),
.Y(n_4359)
);

BUFx10_ASAP7_75t_L g4360 ( 
.A(n_3985),
.Y(n_4360)
);

AOI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_4111),
.A2(n_2073),
.B(n_2041),
.Y(n_4361)
);

AO31x2_ASAP7_75t_L g4362 ( 
.A1(n_4035),
.A2(n_1648),
.A3(n_1547),
.B(n_57),
.Y(n_4362)
);

AO31x2_ASAP7_75t_L g4363 ( 
.A1(n_4040),
.A2(n_59),
.A3(n_55),
.B(n_56),
.Y(n_4363)
);

INVx3_ASAP7_75t_L g4364 ( 
.A(n_3951),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4064),
.Y(n_4365)
);

O2A1O1Ixp33_ASAP7_75t_L g4366 ( 
.A1(n_3979),
.A2(n_64),
.B(n_60),
.C(n_61),
.Y(n_4366)
);

O2A1O1Ixp33_ASAP7_75t_L g4367 ( 
.A1(n_3982),
.A2(n_64),
.B(n_60),
.C(n_61),
.Y(n_4367)
);

AOI22xp5_ASAP7_75t_L g4368 ( 
.A1(n_4063),
.A2(n_1815),
.B1(n_1809),
.B2(n_1681),
.Y(n_4368)
);

BUFx10_ASAP7_75t_L g4369 ( 
.A(n_3992),
.Y(n_4369)
);

A2O1A1Ixp33_ASAP7_75t_L g4370 ( 
.A1(n_4116),
.A2(n_69),
.B(n_65),
.C(n_67),
.Y(n_4370)
);

AOI22xp33_ASAP7_75t_L g4371 ( 
.A1(n_4135),
.A2(n_1815),
.B1(n_1681),
.B2(n_1693),
.Y(n_4371)
);

AOI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_4085),
.A2(n_1815),
.B1(n_1681),
.B2(n_1693),
.Y(n_4372)
);

NOR4xp25_ASAP7_75t_L g4373 ( 
.A(n_4088),
.B(n_71),
.C(n_65),
.D(n_69),
.Y(n_4373)
);

AOI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_4152),
.A2(n_2278),
.B(n_2093),
.Y(n_4374)
);

AOI21xp5_ASAP7_75t_L g4375 ( 
.A1(n_4152),
.A2(n_2278),
.B(n_2093),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4067),
.B(n_71),
.Y(n_4376)
);

NOR2xp33_ASAP7_75t_SL g4377 ( 
.A(n_4150),
.B(n_1683),
.Y(n_4377)
);

OAI21x1_ASAP7_75t_L g4378 ( 
.A1(n_4130),
.A2(n_4154),
.B(n_4036),
.Y(n_4378)
);

AOI21xp33_ASAP7_75t_L g4379 ( 
.A1(n_4091),
.A2(n_1681),
.B(n_1671),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4116),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_3982),
.A2(n_2278),
.B(n_2093),
.Y(n_4381)
);

O2A1O1Ixp33_ASAP7_75t_SL g4382 ( 
.A1(n_4140),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_4382)
);

OAI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4025),
.A2(n_2119),
.B(n_2073),
.Y(n_4383)
);

AO31x2_ASAP7_75t_L g4384 ( 
.A1(n_4085),
.A2(n_77),
.A3(n_75),
.B(n_76),
.Y(n_4384)
);

AO32x2_ASAP7_75t_L g4385 ( 
.A1(n_4085),
.A2(n_79),
.A3(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_3951),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4091),
.B(n_78),
.Y(n_4387)
);

AOI21xp5_ASAP7_75t_L g4388 ( 
.A1(n_4157),
.A2(n_2119),
.B(n_2073),
.Y(n_4388)
);

OAI21x1_ASAP7_75t_L g4389 ( 
.A1(n_4127),
.A2(n_2138),
.B(n_2119),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_3992),
.Y(n_4390)
);

INVxp67_ASAP7_75t_L g4391 ( 
.A(n_4070),
.Y(n_4391)
);

AOI21xp5_ASAP7_75t_L g4392 ( 
.A1(n_4157),
.A2(n_2208),
.B(n_2138),
.Y(n_4392)
);

O2A1O1Ixp33_ASAP7_75t_L g4393 ( 
.A1(n_4147),
.A2(n_83),
.B(n_79),
.C(n_80),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_4092),
.A2(n_4144),
.B(n_4017),
.Y(n_4394)
);

O2A1O1Ixp33_ASAP7_75t_L g4395 ( 
.A1(n_4092),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_4395)
);

BUFx12f_ASAP7_75t_L g4396 ( 
.A(n_4016),
.Y(n_4396)
);

OR2x2_ASAP7_75t_L g4397 ( 
.A(n_4016),
.B(n_1671),
.Y(n_4397)
);

OAI21x1_ASAP7_75t_L g4398 ( 
.A1(n_4017),
.A2(n_2208),
.B(n_2138),
.Y(n_4398)
);

AO31x2_ASAP7_75t_L g4399 ( 
.A1(n_4045),
.A2(n_86),
.A3(n_84),
.B(n_85),
.Y(n_4399)
);

O2A1O1Ixp33_ASAP7_75t_SL g4400 ( 
.A1(n_4045),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_4400)
);

AOI221xp5_ASAP7_75t_L g4401 ( 
.A1(n_4144),
.A2(n_1694),
.B1(n_1693),
.B2(n_1671),
.C(n_89),
.Y(n_4401)
);

BUFx6f_ASAP7_75t_L g4402 ( 
.A(n_4294),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4184),
.Y(n_4403)
);

AOI22xp33_ASAP7_75t_L g4404 ( 
.A1(n_4173),
.A2(n_4071),
.B1(n_4098),
.B2(n_4070),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_4201),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4202),
.Y(n_4406)
);

CKINVDCx8_ASAP7_75t_R g4407 ( 
.A(n_4358),
.Y(n_4407)
);

INVx3_ASAP7_75t_L g4408 ( 
.A(n_4378),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4177),
.Y(n_4409)
);

AOI22xp33_ASAP7_75t_L g4410 ( 
.A1(n_4292),
.A2(n_4132),
.B1(n_4098),
.B2(n_4107),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4200),
.Y(n_4411)
);

BUFx3_ASAP7_75t_L g4412 ( 
.A(n_4264),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_4189),
.B(n_4071),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_4305),
.B(n_4107),
.Y(n_4414)
);

AOI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_4170),
.A2(n_4125),
.B(n_4108),
.Y(n_4415)
);

OAI21xp33_ASAP7_75t_L g4416 ( 
.A1(n_4281),
.A2(n_4373),
.B(n_4291),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4208),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4255),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_4167),
.Y(n_4419)
);

INVx2_ASAP7_75t_SL g4420 ( 
.A(n_4321),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4242),
.Y(n_4421)
);

CKINVDCx11_ASAP7_75t_R g4422 ( 
.A(n_4230),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4260),
.Y(n_4423)
);

CKINVDCx5p33_ASAP7_75t_R g4424 ( 
.A(n_4206),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4319),
.Y(n_4425)
);

INVx2_ASAP7_75t_L g4426 ( 
.A(n_4298),
.Y(n_4426)
);

AOI22xp33_ASAP7_75t_SL g4427 ( 
.A1(n_4171),
.A2(n_4125),
.B1(n_4128),
.B2(n_4108),
.Y(n_4427)
);

OAI22xp5_ASAP7_75t_L g4428 ( 
.A1(n_4181),
.A2(n_4132),
.B1(n_4128),
.B2(n_89),
.Y(n_4428)
);

AOI22xp33_ASAP7_75t_L g4429 ( 
.A1(n_4304),
.A2(n_1694),
.B1(n_1693),
.B2(n_2208),
.Y(n_4429)
);

CKINVDCx9p33_ASAP7_75t_R g4430 ( 
.A(n_4277),
.Y(n_4430)
);

AOI22xp33_ASAP7_75t_L g4431 ( 
.A1(n_4401),
.A2(n_4337),
.B1(n_4296),
.B2(n_4331),
.Y(n_4431)
);

INVx6_ASAP7_75t_L g4432 ( 
.A(n_4325),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_4285),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4178),
.B(n_87),
.Y(n_4434)
);

OAI221xp5_ASAP7_75t_L g4435 ( 
.A1(n_4188),
.A2(n_91),
.B1(n_88),
.B2(n_90),
.C(n_92),
.Y(n_4435)
);

AOI22xp33_ASAP7_75t_L g4436 ( 
.A1(n_4300),
.A2(n_1694),
.B1(n_2209),
.B2(n_1589),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4365),
.Y(n_4437)
);

AND2x4_ASAP7_75t_L g4438 ( 
.A(n_4231),
.B(n_90),
.Y(n_4438)
);

AOI22xp33_ASAP7_75t_L g4439 ( 
.A1(n_4302),
.A2(n_1694),
.B1(n_2209),
.B2(n_1589),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_L g4440 ( 
.A(n_4274),
.B(n_91),
.Y(n_4440)
);

AOI22xp33_ASAP7_75t_L g4441 ( 
.A1(n_4199),
.A2(n_2209),
.B1(n_1584),
.B2(n_1762),
.Y(n_4441)
);

AO21x2_ASAP7_75t_L g4442 ( 
.A1(n_4191),
.A2(n_94),
.B(n_95),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4195),
.B(n_4308),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4262),
.Y(n_4444)
);

NAND2x1p5_ASAP7_75t_L g4445 ( 
.A(n_4380),
.B(n_1683),
.Y(n_4445)
);

AOI222xp33_ASAP7_75t_L g4446 ( 
.A1(n_4250),
.A2(n_4269),
.B1(n_4316),
.B2(n_4336),
.C1(n_4204),
.C2(n_4342),
.Y(n_4446)
);

OAI21xp5_ASAP7_75t_L g4447 ( 
.A1(n_4169),
.A2(n_1683),
.B(n_1584),
.Y(n_4447)
);

INVx5_ASAP7_75t_L g4448 ( 
.A(n_4335),
.Y(n_4448)
);

AOI22xp33_ASAP7_75t_L g4449 ( 
.A1(n_4212),
.A2(n_1762),
.B1(n_1786),
.B2(n_1757),
.Y(n_4449)
);

BUFx3_ASAP7_75t_L g4450 ( 
.A(n_4265),
.Y(n_4450)
);

OAI21xp5_ASAP7_75t_L g4451 ( 
.A1(n_4214),
.A2(n_94),
.B(n_95),
.Y(n_4451)
);

A2O1A1Ixp33_ASAP7_75t_L g4452 ( 
.A1(n_4317),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_4452)
);

OR2x2_ASAP7_75t_L g4453 ( 
.A(n_4271),
.B(n_96),
.Y(n_4453)
);

OAI22xp5_ASAP7_75t_L g4454 ( 
.A1(n_4338),
.A2(n_102),
.B1(n_97),
.B2(n_99),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4263),
.Y(n_4455)
);

OAI221xp5_ASAP7_75t_L g4456 ( 
.A1(n_4339),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.C(n_108),
.Y(n_4456)
);

INVx3_ASAP7_75t_L g4457 ( 
.A(n_4386),
.Y(n_4457)
);

CKINVDCx11_ASAP7_75t_R g4458 ( 
.A(n_4396),
.Y(n_4458)
);

INVx6_ASAP7_75t_L g4459 ( 
.A(n_4311),
.Y(n_4459)
);

BUFx4f_ASAP7_75t_L g4460 ( 
.A(n_4253),
.Y(n_4460)
);

INVx2_ASAP7_75t_L g4461 ( 
.A(n_4273),
.Y(n_4461)
);

CKINVDCx20_ASAP7_75t_R g4462 ( 
.A(n_4227),
.Y(n_4462)
);

OR2x2_ASAP7_75t_L g4463 ( 
.A(n_4213),
.B(n_103),
.Y(n_4463)
);

NAND2x1p5_ASAP7_75t_L g4464 ( 
.A(n_4293),
.B(n_1757),
.Y(n_4464)
);

NOR2xp33_ASAP7_75t_L g4465 ( 
.A(n_4186),
.B(n_109),
.Y(n_4465)
);

NAND2x1p5_ASAP7_75t_L g4466 ( 
.A(n_4329),
.B(n_1757),
.Y(n_4466)
);

AO21x2_ASAP7_75t_L g4467 ( 
.A1(n_4185),
.A2(n_4182),
.B(n_4196),
.Y(n_4467)
);

OAI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4370),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4359),
.Y(n_4469)
);

AOI22xp33_ASAP7_75t_SL g4470 ( 
.A1(n_4254),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_4470)
);

O2A1O1Ixp33_ASAP7_75t_SL g4471 ( 
.A1(n_4367),
.A2(n_117),
.B(n_114),
.C(n_116),
.Y(n_4471)
);

OAI22xp33_ASAP7_75t_L g4472 ( 
.A1(n_4192),
.A2(n_122),
.B1(n_118),
.B2(n_120),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4219),
.Y(n_4473)
);

OAI22xp33_ASAP7_75t_SL g4474 ( 
.A1(n_4385),
.A2(n_122),
.B1(n_118),
.B2(n_120),
.Y(n_4474)
);

AOI22xp33_ASAP7_75t_L g4475 ( 
.A1(n_4190),
.A2(n_4256),
.B1(n_4226),
.B2(n_4238),
.Y(n_4475)
);

A2O1A1Ixp33_ASAP7_75t_L g4476 ( 
.A1(n_4395),
.A2(n_128),
.B(n_124),
.C(n_127),
.Y(n_4476)
);

INVx2_ASAP7_75t_SL g4477 ( 
.A(n_4348),
.Y(n_4477)
);

AOI22xp33_ASAP7_75t_L g4478 ( 
.A1(n_4267),
.A2(n_1762),
.B1(n_1786),
.B2(n_1757),
.Y(n_4478)
);

CKINVDCx5p33_ASAP7_75t_R g4479 ( 
.A(n_4261),
.Y(n_4479)
);

BUFx3_ASAP7_75t_L g4480 ( 
.A(n_4166),
.Y(n_4480)
);

NOR2xp33_ASAP7_75t_L g4481 ( 
.A(n_4179),
.B(n_4237),
.Y(n_4481)
);

AND2x4_ASAP7_75t_L g4482 ( 
.A(n_4257),
.B(n_4364),
.Y(n_4482)
);

OAI22xp33_ASAP7_75t_L g4483 ( 
.A1(n_4327),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4213),
.Y(n_4484)
);

AOI22xp33_ASAP7_75t_L g4485 ( 
.A1(n_4283),
.A2(n_1786),
.B1(n_1762),
.B2(n_1921),
.Y(n_4485)
);

INVx3_ASAP7_75t_L g4486 ( 
.A(n_4369),
.Y(n_4486)
);

AOI22xp33_ASAP7_75t_SL g4487 ( 
.A1(n_4219),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_4487)
);

AOI22xp33_ASAP7_75t_L g4488 ( 
.A1(n_4280),
.A2(n_1786),
.B1(n_1945),
.B2(n_1921),
.Y(n_4488)
);

AOI22xp5_ASAP7_75t_L g4489 ( 
.A1(n_4258),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_4489)
);

OAI221xp5_ASAP7_75t_L g4490 ( 
.A1(n_4187),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_4490)
);

OAI22xp5_ASAP7_75t_L g4491 ( 
.A1(n_4393),
.A2(n_138),
.B1(n_133),
.B2(n_137),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_4219),
.Y(n_4492)
);

O2A1O1Ixp33_ASAP7_75t_L g4493 ( 
.A1(n_4366),
.A2(n_139),
.B(n_137),
.C(n_138),
.Y(n_4493)
);

AOI22xp33_ASAP7_75t_L g4494 ( 
.A1(n_4219),
.A2(n_1945),
.B1(n_1961),
.B2(n_1921),
.Y(n_4494)
);

OAI22xp33_ASAP7_75t_L g4495 ( 
.A1(n_4372),
.A2(n_142),
.B1(n_139),
.B2(n_140),
.Y(n_4495)
);

OAI221xp5_ASAP7_75t_L g4496 ( 
.A1(n_4174),
.A2(n_145),
.B1(n_140),
.B2(n_144),
.C(n_146),
.Y(n_4496)
);

CKINVDCx11_ASAP7_75t_R g4497 ( 
.A(n_4360),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4363),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4233),
.B(n_144),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4363),
.Y(n_4500)
);

OAI22xp5_ASAP7_75t_L g4501 ( 
.A1(n_4322),
.A2(n_4345),
.B1(n_4225),
.B2(n_4232),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4362),
.Y(n_4502)
);

NOR2x1_ASAP7_75t_SL g4503 ( 
.A(n_4290),
.B(n_1612),
.Y(n_4503)
);

BUFx2_ASAP7_75t_SL g4504 ( 
.A(n_4183),
.Y(n_4504)
);

NAND2x1p5_ASAP7_75t_L g4505 ( 
.A(n_4312),
.B(n_1612),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4362),
.Y(n_4506)
);

AOI22xp33_ASAP7_75t_L g4507 ( 
.A1(n_4357),
.A2(n_1961),
.B1(n_1980),
.B2(n_1945),
.Y(n_4507)
);

INVx4_ASAP7_75t_L g4508 ( 
.A(n_4335),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4326),
.B(n_146),
.Y(n_4509)
);

OAI21xp5_ASAP7_75t_L g4510 ( 
.A1(n_4175),
.A2(n_147),
.B(n_148),
.Y(n_4510)
);

INVx6_ASAP7_75t_L g4511 ( 
.A(n_4253),
.Y(n_4511)
);

OAI22xp33_ASAP7_75t_L g4512 ( 
.A1(n_4275),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_SL g4513 ( 
.A(n_4268),
.B(n_1606),
.Y(n_4513)
);

OAI22xp5_ASAP7_75t_L g4514 ( 
.A1(n_4217),
.A2(n_152),
.B1(n_149),
.B2(n_151),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4320),
.Y(n_4515)
);

A2O1A1Ixp33_ASAP7_75t_L g4516 ( 
.A1(n_4193),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_4516)
);

INVx3_ASAP7_75t_L g4517 ( 
.A(n_4240),
.Y(n_4517)
);

OAI22xp5_ASAP7_75t_L g4518 ( 
.A1(n_4340),
.A2(n_158),
.B1(n_154),
.B2(n_155),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4194),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4350),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4323),
.B(n_160),
.Y(n_4521)
);

BUFx2_ASAP7_75t_L g4522 ( 
.A(n_4390),
.Y(n_4522)
);

OAI22xp33_ASAP7_75t_L g4523 ( 
.A1(n_4387),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_4523)
);

O2A1O1Ixp33_ASAP7_75t_SL g4524 ( 
.A1(n_4376),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_4176),
.Y(n_4525)
);

AOI22xp33_ASAP7_75t_L g4526 ( 
.A1(n_4347),
.A2(n_1961),
.B1(n_1980),
.B2(n_1945),
.Y(n_4526)
);

AOI22xp33_ASAP7_75t_L g4527 ( 
.A1(n_4297),
.A2(n_1980),
.B1(n_1995),
.B2(n_1961),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4176),
.Y(n_4528)
);

INVxp67_ASAP7_75t_L g4529 ( 
.A(n_4247),
.Y(n_4529)
);

AOI22xp33_ASAP7_75t_SL g4530 ( 
.A1(n_4385),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_4530)
);

AOI22xp5_ASAP7_75t_L g4531 ( 
.A1(n_4251),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_4531)
);

AOI22xp33_ASAP7_75t_L g4532 ( 
.A1(n_4207),
.A2(n_1995),
.B1(n_2013),
.B2(n_1980),
.Y(n_4532)
);

OR2x6_ASAP7_75t_L g4533 ( 
.A(n_4210),
.B(n_4215),
.Y(n_4533)
);

A2O1A1Ixp33_ASAP7_75t_L g4534 ( 
.A1(n_4211),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_4534)
);

OAI22xp5_ASAP7_75t_L g4535 ( 
.A1(n_4314),
.A2(n_172),
.B1(n_169),
.B2(n_171),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4385),
.Y(n_4536)
);

HB1xp67_ASAP7_75t_L g4537 ( 
.A(n_4180),
.Y(n_4537)
);

AND2x4_ASAP7_75t_L g4538 ( 
.A(n_4394),
.B(n_171),
.Y(n_4538)
);

HB1xp67_ASAP7_75t_L g4539 ( 
.A(n_4180),
.Y(n_4539)
);

OAI22xp5_ASAP7_75t_L g4540 ( 
.A1(n_4391),
.A2(n_177),
.B1(n_174),
.B2(n_175),
.Y(n_4540)
);

OAI22xp5_ASAP7_75t_L g4541 ( 
.A1(n_4229),
.A2(n_178),
.B1(n_174),
.B2(n_175),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4399),
.Y(n_4542)
);

AOI21xp5_ASAP7_75t_L g4543 ( 
.A1(n_4246),
.A2(n_2013),
.B(n_1995),
.Y(n_4543)
);

OAI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4289),
.A2(n_4334),
.B1(n_4309),
.B2(n_4371),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_4176),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4399),
.Y(n_4546)
);

INVx2_ASAP7_75t_L g4547 ( 
.A(n_4235),
.Y(n_4547)
);

AOI22xp33_ASAP7_75t_L g4548 ( 
.A1(n_4310),
.A2(n_2013),
.B1(n_2018),
.B2(n_1995),
.Y(n_4548)
);

AOI21xp33_ASAP7_75t_L g4549 ( 
.A1(n_4397),
.A2(n_178),
.B(n_180),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4384),
.Y(n_4550)
);

HB1xp67_ASAP7_75t_L g4551 ( 
.A(n_4235),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4384),
.Y(n_4552)
);

AOI22xp5_ASAP7_75t_L g4553 ( 
.A1(n_4351),
.A2(n_183),
.B1(n_180),
.B2(n_182),
.Y(n_4553)
);

AOI22xp33_ASAP7_75t_L g4554 ( 
.A1(n_4218),
.A2(n_4332),
.B1(n_4349),
.B2(n_4346),
.Y(n_4554)
);

A2O1A1Ixp33_ASAP7_75t_L g4555 ( 
.A1(n_4306),
.A2(n_185),
.B(n_182),
.C(n_184),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_SL g4556 ( 
.A(n_4335),
.B(n_186),
.Y(n_4556)
);

AND2x4_ASAP7_75t_L g4557 ( 
.A(n_4270),
.B(n_186),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4353),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4168),
.Y(n_4559)
);

BUFx3_ASAP7_75t_L g4560 ( 
.A(n_4197),
.Y(n_4560)
);

AOI22xp33_ASAP7_75t_L g4561 ( 
.A1(n_4286),
.A2(n_2018),
.B1(n_2036),
.B2(n_2013),
.Y(n_4561)
);

AND2x4_ASAP7_75t_L g4562 ( 
.A(n_4245),
.B(n_4290),
.Y(n_4562)
);

AOI22xp33_ASAP7_75t_L g4563 ( 
.A1(n_4307),
.A2(n_2036),
.B1(n_2042),
.B2(n_2018),
.Y(n_4563)
);

OAI21xp33_ASAP7_75t_L g4564 ( 
.A1(n_4209),
.A2(n_187),
.B(n_188),
.Y(n_4564)
);

OAI22xp5_ASAP7_75t_L g4565 ( 
.A1(n_4368),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_4565)
);

AOI22xp33_ASAP7_75t_L g4566 ( 
.A1(n_4383),
.A2(n_2036),
.B1(n_2042),
.B2(n_2018),
.Y(n_4566)
);

OAI22xp33_ASAP7_75t_L g4567 ( 
.A1(n_4377),
.A2(n_4341),
.B1(n_4328),
.B2(n_4299),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4168),
.B(n_189),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4168),
.Y(n_4569)
);

AOI22xp33_ASAP7_75t_L g4570 ( 
.A1(n_4276),
.A2(n_2042),
.B1(n_2059),
.B2(n_2036),
.Y(n_4570)
);

OAI22xp5_ASAP7_75t_L g4571 ( 
.A1(n_4315),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_4571)
);

CKINVDCx8_ASAP7_75t_R g4572 ( 
.A(n_4341),
.Y(n_4572)
);

BUFx2_ASAP7_75t_L g4573 ( 
.A(n_4279),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4330),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4330),
.Y(n_4575)
);

AOI22xp33_ASAP7_75t_L g4576 ( 
.A1(n_4248),
.A2(n_2059),
.B1(n_2070),
.B2(n_2042),
.Y(n_4576)
);

CKINVDCx20_ASAP7_75t_R g4577 ( 
.A(n_4236),
.Y(n_4577)
);

AND2x4_ASAP7_75t_L g4578 ( 
.A(n_4288),
.B(n_192),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4344),
.Y(n_4579)
);

OAI221xp5_ASAP7_75t_L g4580 ( 
.A1(n_4382),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.C(n_199),
.Y(n_4580)
);

OAI221xp5_ASAP7_75t_L g4581 ( 
.A1(n_4301),
.A2(n_200),
.B1(n_194),
.B2(n_199),
.C(n_201),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4249),
.Y(n_4582)
);

AND2x2_ASAP7_75t_L g4583 ( 
.A(n_4279),
.B(n_4324),
.Y(n_4583)
);

AND2x4_ASAP7_75t_L g4584 ( 
.A(n_4333),
.B(n_200),
.Y(n_4584)
);

AOI22xp33_ASAP7_75t_SL g4585 ( 
.A1(n_4400),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_4585)
);

AOI22xp33_ASAP7_75t_L g4586 ( 
.A1(n_4379),
.A2(n_2070),
.B1(n_2074),
.B2(n_2059),
.Y(n_4586)
);

HB1xp67_ASAP7_75t_L g4587 ( 
.A(n_4249),
.Y(n_4587)
);

AO31x2_ASAP7_75t_L g4588 ( 
.A1(n_4484),
.A2(n_4313),
.A3(n_4287),
.B(n_4223),
.Y(n_4588)
);

OR2x6_ASAP7_75t_L g4589 ( 
.A(n_4533),
.B(n_4222),
.Y(n_4589)
);

BUFx6f_ASAP7_75t_L g4590 ( 
.A(n_4402),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4409),
.Y(n_4591)
);

AOI21xp5_ASAP7_75t_L g4592 ( 
.A1(n_4510),
.A2(n_4272),
.B(n_4352),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4411),
.Y(n_4593)
);

OR2x6_ASAP7_75t_L g4594 ( 
.A(n_4533),
.B(n_4343),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4417),
.Y(n_4595)
);

HB1xp67_ASAP7_75t_L g4596 ( 
.A(n_4498),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4457),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4421),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4559),
.B(n_4344),
.Y(n_4599)
);

INVx4_ASAP7_75t_L g4600 ( 
.A(n_4402),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4457),
.Y(n_4601)
);

O2A1O1Ixp33_ASAP7_75t_L g4602 ( 
.A1(n_4435),
.A2(n_4221),
.B(n_4220),
.C(n_4243),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4423),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4425),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4437),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4403),
.Y(n_4606)
);

INVx2_ASAP7_75t_L g4607 ( 
.A(n_4405),
.Y(n_4607)
);

AO21x1_ASAP7_75t_SL g4608 ( 
.A1(n_4536),
.A2(n_4318),
.B(n_4172),
.Y(n_4608)
);

HB1xp67_ASAP7_75t_L g4609 ( 
.A(n_4500),
.Y(n_4609)
);

AOI21x1_ASAP7_75t_L g4610 ( 
.A1(n_4568),
.A2(n_4354),
.B(n_4303),
.Y(n_4610)
);

HB1xp67_ASAP7_75t_L g4611 ( 
.A(n_4550),
.Y(n_4611)
);

AOI22xp33_ASAP7_75t_L g4612 ( 
.A1(n_4416),
.A2(n_4234),
.B1(n_4355),
.B2(n_4381),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4406),
.Y(n_4613)
);

OR2x2_ASAP7_75t_L g4614 ( 
.A(n_4426),
.B(n_4244),
.Y(n_4614)
);

BUFx2_ASAP7_75t_L g4615 ( 
.A(n_4482),
.Y(n_4615)
);

HB1xp67_ASAP7_75t_L g4616 ( 
.A(n_4552),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4418),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4419),
.Y(n_4618)
);

OAI22xp5_ASAP7_75t_L g4619 ( 
.A1(n_4530),
.A2(n_4224),
.B1(n_4228),
.B2(n_4278),
.Y(n_4619)
);

INVx4_ASAP7_75t_L g4620 ( 
.A(n_4402),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4469),
.Y(n_4621)
);

BUFx3_ASAP7_75t_L g4622 ( 
.A(n_4462),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4444),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4455),
.Y(n_4624)
);

BUFx2_ASAP7_75t_L g4625 ( 
.A(n_4482),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4443),
.B(n_4515),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4461),
.Y(n_4627)
);

OR2x6_ASAP7_75t_L g4628 ( 
.A(n_4533),
.B(n_4259),
.Y(n_4628)
);

HB1xp67_ASAP7_75t_L g4629 ( 
.A(n_4542),
.Y(n_4629)
);

AO21x2_ASAP7_75t_L g4630 ( 
.A1(n_4519),
.A2(n_4203),
.B(n_4216),
.Y(n_4630)
);

AND2x4_ASAP7_75t_L g4631 ( 
.A(n_4408),
.B(n_4244),
.Y(n_4631)
);

AND2x4_ASAP7_75t_L g4632 ( 
.A(n_4408),
.B(n_4398),
.Y(n_4632)
);

AOI21x1_ASAP7_75t_L g4633 ( 
.A1(n_4509),
.A2(n_4284),
.B(n_4295),
.Y(n_4633)
);

OAI21x1_ASAP7_75t_L g4634 ( 
.A1(n_4574),
.A2(n_4266),
.B(n_4198),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4433),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4546),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4414),
.Y(n_4637)
);

INVx2_ASAP7_75t_SL g4638 ( 
.A(n_4432),
.Y(n_4638)
);

HB1xp67_ASAP7_75t_L g4639 ( 
.A(n_4502),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4413),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4506),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4463),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4569),
.B(n_4389),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4504),
.B(n_4172),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4520),
.Y(n_4645)
);

INVx2_ASAP7_75t_L g4646 ( 
.A(n_4473),
.Y(n_4646)
);

BUFx3_ASAP7_75t_L g4647 ( 
.A(n_4422),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4492),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4525),
.B(n_4205),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4477),
.B(n_4172),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4537),
.Y(n_4651)
);

NOR2xp33_ASAP7_75t_L g4652 ( 
.A(n_4434),
.B(n_4252),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_4517),
.Y(n_4653)
);

INVx4_ASAP7_75t_L g4654 ( 
.A(n_4432),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4517),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_4573),
.Y(n_4656)
);

BUFx4f_ASAP7_75t_SL g4657 ( 
.A(n_4450),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4539),
.Y(n_4658)
);

BUFx2_ASAP7_75t_SL g4659 ( 
.A(n_4407),
.Y(n_4659)
);

INVx3_ASAP7_75t_L g4660 ( 
.A(n_4480),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4453),
.Y(n_4661)
);

AND2x2_ASAP7_75t_L g4662 ( 
.A(n_4420),
.B(n_4356),
.Y(n_4662)
);

HB1xp67_ASAP7_75t_L g4663 ( 
.A(n_4528),
.Y(n_4663)
);

OAI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_4510),
.A2(n_4361),
.B(n_4241),
.Y(n_4664)
);

HB1xp67_ASAP7_75t_L g4665 ( 
.A(n_4545),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4529),
.Y(n_4666)
);

INVx3_ASAP7_75t_L g4667 ( 
.A(n_4486),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4522),
.B(n_4486),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4558),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4438),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4551),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4438),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4587),
.B(n_204),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4575),
.Y(n_4674)
);

INVx2_ASAP7_75t_L g4675 ( 
.A(n_4583),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4579),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4547),
.Y(n_4677)
);

NOR2xp33_ASAP7_75t_L g4678 ( 
.A(n_4521),
.B(n_204),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4412),
.B(n_4282),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4467),
.Y(n_4680)
);

HB1xp67_ASAP7_75t_L g4681 ( 
.A(n_4582),
.Y(n_4681)
);

O2A1O1Ixp33_ASAP7_75t_SL g4682 ( 
.A1(n_4452),
.A2(n_4239),
.B(n_209),
.C(n_206),
.Y(n_4682)
);

HB1xp67_ASAP7_75t_L g4683 ( 
.A(n_4467),
.Y(n_4683)
);

O2A1O1Ixp5_ASAP7_75t_L g4684 ( 
.A1(n_4451),
.A2(n_4472),
.B(n_4476),
.C(n_4468),
.Y(n_4684)
);

HB1xp67_ASAP7_75t_L g4685 ( 
.A(n_4442),
.Y(n_4685)
);

INVx3_ASAP7_75t_L g4686 ( 
.A(n_4560),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4538),
.Y(n_4687)
);

INVx3_ASAP7_75t_L g4688 ( 
.A(n_4511),
.Y(n_4688)
);

BUFx3_ASAP7_75t_L g4689 ( 
.A(n_4424),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4442),
.Y(n_4690)
);

INVx3_ASAP7_75t_SL g4691 ( 
.A(n_4479),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4562),
.Y(n_4692)
);

HB1xp67_ASAP7_75t_L g4693 ( 
.A(n_4464),
.Y(n_4693)
);

CKINVDCx14_ASAP7_75t_R g4694 ( 
.A(n_4458),
.Y(n_4694)
);

OR2x2_ASAP7_75t_L g4695 ( 
.A(n_4538),
.B(n_4374),
.Y(n_4695)
);

OR2x2_ASAP7_75t_L g4696 ( 
.A(n_4499),
.B(n_4375),
.Y(n_4696)
);

OAI21x1_ASAP7_75t_L g4697 ( 
.A1(n_4445),
.A2(n_4392),
.B(n_4388),
.Y(n_4697)
);

CKINVDCx20_ASAP7_75t_R g4698 ( 
.A(n_4497),
.Y(n_4698)
);

CKINVDCx11_ASAP7_75t_R g4699 ( 
.A(n_4572),
.Y(n_4699)
);

OR2x6_ASAP7_75t_L g4700 ( 
.A(n_4508),
.B(n_4562),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4474),
.Y(n_4701)
);

BUFx3_ASAP7_75t_L g4702 ( 
.A(n_4511),
.Y(n_4702)
);

INVx4_ASAP7_75t_SL g4703 ( 
.A(n_4459),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4474),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4557),
.Y(n_4705)
);

INVx3_ASAP7_75t_L g4706 ( 
.A(n_4459),
.Y(n_4706)
);

HB1xp67_ASAP7_75t_L g4707 ( 
.A(n_4557),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4578),
.Y(n_4708)
);

HB1xp67_ASAP7_75t_L g4709 ( 
.A(n_4578),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4584),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4584),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4481),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4427),
.Y(n_4713)
);

OAI211xp5_ASAP7_75t_SL g4714 ( 
.A1(n_4416),
.A2(n_209),
.B(n_206),
.C(n_207),
.Y(n_4714)
);

HB1xp67_ASAP7_75t_L g4715 ( 
.A(n_4448),
.Y(n_4715)
);

OR2x6_ASAP7_75t_L g4716 ( 
.A(n_4508),
.B(n_2059),
.Y(n_4716)
);

INVx5_ASAP7_75t_L g4717 ( 
.A(n_4448),
.Y(n_4717)
);

BUFx6f_ASAP7_75t_L g4718 ( 
.A(n_4460),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4505),
.Y(n_4719)
);

AND2x4_ASAP7_75t_L g4720 ( 
.A(n_4448),
.B(n_207),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4440),
.Y(n_4721)
);

OAI21x1_ASAP7_75t_L g4722 ( 
.A1(n_4415),
.A2(n_1633),
.B(n_1606),
.Y(n_4722)
);

AO31x2_ASAP7_75t_L g4723 ( 
.A1(n_4503),
.A2(n_212),
.A3(n_210),
.B(n_211),
.Y(n_4723)
);

INVx2_ASAP7_75t_SL g4724 ( 
.A(n_4460),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4524),
.Y(n_4725)
);

INVx3_ASAP7_75t_L g4726 ( 
.A(n_4466),
.Y(n_4726)
);

AOI221xp5_ASAP7_75t_L g4727 ( 
.A1(n_4496),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.C(n_214),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4430),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4531),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4531),
.Y(n_4730)
);

OAI21x1_ASAP7_75t_L g4731 ( 
.A1(n_4447),
.A2(n_1633),
.B(n_1606),
.Y(n_4731)
);

AOI22xp33_ASAP7_75t_L g4732 ( 
.A1(n_4701),
.A2(n_4456),
.B1(n_4501),
.B2(n_4490),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4611),
.Y(n_4733)
);

AOI22xp33_ASAP7_75t_L g4734 ( 
.A1(n_4704),
.A2(n_4581),
.B1(n_4454),
.B2(n_4580),
.Y(n_4734)
);

OAI22xp5_ASAP7_75t_L g4735 ( 
.A1(n_4729),
.A2(n_4431),
.B1(n_4489),
.B2(n_4553),
.Y(n_4735)
);

AOI22xp33_ASAP7_75t_L g4736 ( 
.A1(n_4730),
.A2(n_4446),
.B1(n_4577),
.B2(n_4564),
.Y(n_4736)
);

AOI22xp33_ASAP7_75t_L g4737 ( 
.A1(n_4727),
.A2(n_4446),
.B1(n_4564),
.B2(n_4491),
.Y(n_4737)
);

OAI221xp5_ASAP7_75t_L g4738 ( 
.A1(n_4684),
.A2(n_4470),
.B1(n_4475),
.B2(n_4465),
.C(n_4489),
.Y(n_4738)
);

AOI33xp33_ASAP7_75t_L g4739 ( 
.A1(n_4725),
.A2(n_4523),
.A3(n_4487),
.B1(n_4585),
.B2(n_4483),
.B3(n_4471),
.Y(n_4739)
);

BUFx6f_ASAP7_75t_L g4740 ( 
.A(n_4590),
.Y(n_4740)
);

O2A1O1Ixp33_ASAP7_75t_L g4741 ( 
.A1(n_4714),
.A2(n_4493),
.B(n_4516),
.C(n_4534),
.Y(n_4741)
);

OAI221xp5_ASAP7_75t_L g4742 ( 
.A1(n_4684),
.A2(n_4553),
.B1(n_4518),
.B2(n_4428),
.C(n_4556),
.Y(n_4742)
);

OAI221xp5_ASAP7_75t_L g4743 ( 
.A1(n_4727),
.A2(n_4556),
.B1(n_4541),
.B2(n_4404),
.C(n_4555),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4611),
.Y(n_4744)
);

NAND3xp33_ASAP7_75t_L g4745 ( 
.A(n_4685),
.B(n_4549),
.C(n_4514),
.Y(n_4745)
);

AOI22xp33_ASAP7_75t_SL g4746 ( 
.A1(n_4728),
.A2(n_4447),
.B1(n_4565),
.B2(n_4571),
.Y(n_4746)
);

OAI22xp5_ASAP7_75t_L g4747 ( 
.A1(n_4712),
.A2(n_4410),
.B1(n_4512),
.B2(n_4495),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4615),
.B(n_4527),
.Y(n_4748)
);

AOI221xp5_ASAP7_75t_L g4749 ( 
.A1(n_4714),
.A2(n_4540),
.B1(n_4535),
.B2(n_4513),
.C(n_4567),
.Y(n_4749)
);

OAI22xp5_ASAP7_75t_L g4750 ( 
.A1(n_4713),
.A2(n_4554),
.B1(n_4526),
.B2(n_4548),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4642),
.B(n_4429),
.Y(n_4751)
);

AOI222xp33_ASAP7_75t_L g4752 ( 
.A1(n_4678),
.A2(n_4544),
.B1(n_4449),
.B2(n_4439),
.C1(n_4436),
.C2(n_215),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_L g4753 ( 
.A(n_4666),
.B(n_4532),
.Y(n_4753)
);

INVx2_ASAP7_75t_L g4754 ( 
.A(n_4708),
.Y(n_4754)
);

CKINVDCx6p67_ASAP7_75t_R g4755 ( 
.A(n_4647),
.Y(n_4755)
);

NOR2xp33_ASAP7_75t_L g4756 ( 
.A(n_4654),
.B(n_213),
.Y(n_4756)
);

AOI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_4592),
.A2(n_4543),
.B(n_4488),
.Y(n_4757)
);

AOI22xp33_ASAP7_75t_L g4758 ( 
.A1(n_4664),
.A2(n_4441),
.B1(n_4485),
.B2(n_4507),
.Y(n_4758)
);

AOI22xp33_ASAP7_75t_L g4759 ( 
.A1(n_4664),
.A2(n_4566),
.B1(n_4494),
.B2(n_4576),
.Y(n_4759)
);

AOI22xp33_ASAP7_75t_L g4760 ( 
.A1(n_4687),
.A2(n_4586),
.B1(n_4561),
.B2(n_4563),
.Y(n_4760)
);

CKINVDCx5p33_ASAP7_75t_R g4761 ( 
.A(n_4694),
.Y(n_4761)
);

NOR2xp33_ASAP7_75t_L g4762 ( 
.A(n_4654),
.B(n_214),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4707),
.B(n_4645),
.Y(n_4763)
);

AOI21xp5_ASAP7_75t_L g4764 ( 
.A1(n_4592),
.A2(n_4570),
.B(n_4478),
.Y(n_4764)
);

AND2x4_ASAP7_75t_L g4765 ( 
.A(n_4700),
.B(n_216),
.Y(n_4765)
);

INVx8_ASAP7_75t_L g4766 ( 
.A(n_4590),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4710),
.Y(n_4767)
);

OAI221xp5_ASAP7_75t_L g4768 ( 
.A1(n_4678),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.C(n_221),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4707),
.B(n_219),
.Y(n_4769)
);

OAI221xp5_ASAP7_75t_L g4770 ( 
.A1(n_4705),
.A2(n_223),
.B1(n_220),
.B2(n_221),
.C(n_225),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4709),
.B(n_226),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4616),
.Y(n_4772)
);

CKINVDCx5p33_ASAP7_75t_R g4773 ( 
.A(n_4659),
.Y(n_4773)
);

HB1xp67_ASAP7_75t_L g4774 ( 
.A(n_4616),
.Y(n_4774)
);

NAND3xp33_ASAP7_75t_L g4775 ( 
.A(n_4685),
.B(n_227),
.C(n_228),
.Y(n_4775)
);

OAI221xp5_ASAP7_75t_L g4776 ( 
.A1(n_4652),
.A2(n_231),
.B1(n_227),
.B2(n_229),
.C(n_233),
.Y(n_4776)
);

AOI21xp33_ASAP7_75t_L g4777 ( 
.A1(n_4594),
.A2(n_231),
.B(n_234),
.Y(n_4777)
);

INVx2_ASAP7_75t_L g4778 ( 
.A(n_4711),
.Y(n_4778)
);

OR2x2_ASAP7_75t_L g4779 ( 
.A(n_4661),
.B(n_235),
.Y(n_4779)
);

OAI22xp5_ASAP7_75t_L g4780 ( 
.A1(n_4696),
.A2(n_239),
.B1(n_236),
.B2(n_238),
.Y(n_4780)
);

OAI21xp5_ASAP7_75t_L g4781 ( 
.A1(n_4682),
.A2(n_238),
.B(n_239),
.Y(n_4781)
);

OAI22xp33_ASAP7_75t_L g4782 ( 
.A1(n_4717),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4625),
.B(n_241),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4709),
.B(n_242),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4640),
.B(n_243),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4641),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4692),
.B(n_244),
.Y(n_4787)
);

NAND3xp33_ASAP7_75t_L g4788 ( 
.A(n_4690),
.B(n_4673),
.C(n_4612),
.Y(n_4788)
);

AOI22xp33_ASAP7_75t_L g4789 ( 
.A1(n_4652),
.A2(n_2074),
.B1(n_2077),
.B2(n_2070),
.Y(n_4789)
);

OAI211xp5_ASAP7_75t_L g4790 ( 
.A1(n_4673),
.A2(n_247),
.B(n_244),
.C(n_246),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4596),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4637),
.B(n_248),
.Y(n_4792)
);

AOI222xp33_ASAP7_75t_L g4793 ( 
.A1(n_4721),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.C1(n_252),
.C2(n_254),
.Y(n_4793)
);

OAI22xp33_ASAP7_75t_L g4794 ( 
.A1(n_4717),
.A2(n_257),
.B1(n_254),
.B2(n_255),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4596),
.Y(n_4795)
);

AOI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_4602),
.A2(n_257),
.B(n_258),
.Y(n_4796)
);

OAI22xp33_ASAP7_75t_L g4797 ( 
.A1(n_4717),
.A2(n_262),
.B1(n_258),
.B2(n_261),
.Y(n_4797)
);

AOI22xp33_ASAP7_75t_L g4798 ( 
.A1(n_4679),
.A2(n_2074),
.B1(n_2077),
.B2(n_2070),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4646),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4686),
.B(n_264),
.Y(n_4800)
);

AOI21xp5_ASAP7_75t_L g4801 ( 
.A1(n_4602),
.A2(n_264),
.B(n_265),
.Y(n_4801)
);

AOI221xp5_ASAP7_75t_L g4802 ( 
.A1(n_4619),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.C(n_268),
.Y(n_4802)
);

AOI22xp33_ASAP7_75t_L g4803 ( 
.A1(n_4594),
.A2(n_2077),
.B1(n_2083),
.B2(n_2074),
.Y(n_4803)
);

AOI22xp5_ASAP7_75t_L g4804 ( 
.A1(n_4619),
.A2(n_1635),
.B1(n_1633),
.B2(n_270),
.Y(n_4804)
);

AOI22xp33_ASAP7_75t_SL g4805 ( 
.A1(n_4657),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_4805)
);

OAI221xp5_ASAP7_75t_L g4806 ( 
.A1(n_4695),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_4806)
);

OAI21x1_ASAP7_75t_L g4807 ( 
.A1(n_4680),
.A2(n_1635),
.B(n_275),
.Y(n_4807)
);

BUFx8_ASAP7_75t_SL g4808 ( 
.A(n_4698),
.Y(n_4808)
);

AOI21x1_ASAP7_75t_L g4809 ( 
.A1(n_4715),
.A2(n_4683),
.B(n_4629),
.Y(n_4809)
);

AOI22xp33_ASAP7_75t_L g4810 ( 
.A1(n_4594),
.A2(n_2077),
.B1(n_2087),
.B2(n_2083),
.Y(n_4810)
);

AOI211xp5_ASAP7_75t_L g4811 ( 
.A1(n_4720),
.A2(n_285),
.B(n_278),
.C(n_280),
.Y(n_4811)
);

AOI221xp5_ASAP7_75t_L g4812 ( 
.A1(n_4651),
.A2(n_4658),
.B1(n_4636),
.B2(n_4593),
.C(n_4598),
.Y(n_4812)
);

AOI221xp5_ASAP7_75t_L g4813 ( 
.A1(n_4591),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4609),
.Y(n_4814)
);

OAI211xp5_ASAP7_75t_L g4815 ( 
.A1(n_4612),
.A2(n_291),
.B(n_287),
.C(n_289),
.Y(n_4815)
);

OAI21xp5_ASAP7_75t_L g4816 ( 
.A1(n_4720),
.A2(n_292),
.B(n_293),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4609),
.Y(n_4817)
);

INVx2_ASAP7_75t_L g4818 ( 
.A(n_4648),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4650),
.B(n_293),
.Y(n_4819)
);

INVxp67_ASAP7_75t_L g4820 ( 
.A(n_4595),
.Y(n_4820)
);

AOI22xp33_ASAP7_75t_L g4821 ( 
.A1(n_4589),
.A2(n_2083),
.B1(n_2115),
.B2(n_2087),
.Y(n_4821)
);

INVx1_ASAP7_75t_SL g4822 ( 
.A(n_4715),
.Y(n_4822)
);

AOI22xp33_ASAP7_75t_L g4823 ( 
.A1(n_4589),
.A2(n_2083),
.B1(n_2115),
.B2(n_2087),
.Y(n_4823)
);

OAI22xp33_ASAP7_75t_L g4824 ( 
.A1(n_4717),
.A2(n_298),
.B1(n_294),
.B2(n_297),
.Y(n_4824)
);

OAI22xp33_ASAP7_75t_L g4825 ( 
.A1(n_4589),
.A2(n_299),
.B1(n_294),
.B2(n_298),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4626),
.B(n_299),
.Y(n_4826)
);

AOI22xp33_ASAP7_75t_L g4827 ( 
.A1(n_4693),
.A2(n_2087),
.B1(n_2117),
.B2(n_2115),
.Y(n_4827)
);

AOI221xp5_ASAP7_75t_L g4828 ( 
.A1(n_4603),
.A2(n_300),
.B1(n_301),
.B2(n_304),
.C(n_305),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4639),
.Y(n_4829)
);

INVxp67_ASAP7_75t_L g4830 ( 
.A(n_4604),
.Y(n_4830)
);

INVx11_ASAP7_75t_L g4831 ( 
.A(n_4657),
.Y(n_4831)
);

AOI222xp33_ASAP7_75t_L g4832 ( 
.A1(n_4600),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.C1(n_309),
.C2(n_311),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4639),
.Y(n_4833)
);

AOI22xp5_ASAP7_75t_L g4834 ( 
.A1(n_4693),
.A2(n_1635),
.B1(n_311),
.B2(n_306),
.Y(n_4834)
);

OAI21x1_ASAP7_75t_L g4835 ( 
.A1(n_4599),
.A2(n_309),
.B(n_312),
.Y(n_4835)
);

OAI22xp33_ASAP7_75t_L g4836 ( 
.A1(n_4700),
.A2(n_316),
.B1(n_312),
.B2(n_314),
.Y(n_4836)
);

AOI22xp33_ASAP7_75t_L g4837 ( 
.A1(n_4670),
.A2(n_2117),
.B1(n_2150),
.B2(n_2115),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4686),
.B(n_318),
.Y(n_4838)
);

AOI22xp33_ASAP7_75t_L g4839 ( 
.A1(n_4672),
.A2(n_4662),
.B1(n_4620),
.B2(n_4600),
.Y(n_4839)
);

AOI22xp5_ASAP7_75t_L g4840 ( 
.A1(n_4620),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4629),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4674),
.Y(n_4842)
);

HB1xp67_ASAP7_75t_L g4843 ( 
.A(n_4671),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4597),
.Y(n_4844)
);

BUFx4f_ASAP7_75t_SL g4845 ( 
.A(n_4689),
.Y(n_4845)
);

AOI22xp33_ASAP7_75t_SL g4846 ( 
.A1(n_4590),
.A2(n_322),
.B1(n_319),
.B2(n_320),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_4621),
.B(n_322),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_L g4848 ( 
.A(n_4606),
.B(n_323),
.Y(n_4848)
);

AOI22xp33_ASAP7_75t_L g4849 ( 
.A1(n_4638),
.A2(n_2150),
.B1(n_2167),
.B2(n_2117),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4601),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4676),
.Y(n_4851)
);

AOI22xp5_ASAP7_75t_L g4852 ( 
.A1(n_4668),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4613),
.B(n_326),
.Y(n_4853)
);

AOI22xp5_ASAP7_75t_L g4854 ( 
.A1(n_4700),
.A2(n_329),
.B1(n_326),
.B2(n_328),
.Y(n_4854)
);

INVx11_ASAP7_75t_L g4855 ( 
.A(n_4703),
.Y(n_4855)
);

BUFx3_ASAP7_75t_L g4856 ( 
.A(n_4622),
.Y(n_4856)
);

INVx3_ASAP7_75t_L g4857 ( 
.A(n_4706),
.Y(n_4857)
);

OAI22xp33_ASAP7_75t_L g4858 ( 
.A1(n_4716),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4656),
.Y(n_4859)
);

NOR2xp33_ASAP7_75t_L g4860 ( 
.A(n_4691),
.B(n_331),
.Y(n_4860)
);

OAI22xp33_ASAP7_75t_L g4861 ( 
.A1(n_4716),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_4861)
);

CKINVDCx11_ASAP7_75t_R g4862 ( 
.A(n_4699),
.Y(n_4862)
);

BUFx4f_ASAP7_75t_SL g4863 ( 
.A(n_4718),
.Y(n_4863)
);

AOI211xp5_ASAP7_75t_L g4864 ( 
.A1(n_4644),
.A2(n_337),
.B(n_333),
.C(n_334),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4617),
.B(n_4618),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_4857),
.B(n_4660),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4786),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4809),
.Y(n_4868)
);

INVx6_ASAP7_75t_L g4869 ( 
.A(n_4766),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4842),
.Y(n_4870)
);

BUFx3_ASAP7_75t_L g4871 ( 
.A(n_4808),
.Y(n_4871)
);

BUFx3_ASAP7_75t_L g4872 ( 
.A(n_4862),
.Y(n_4872)
);

AND2x2_ASAP7_75t_L g4873 ( 
.A(n_4857),
.B(n_4660),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4822),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4839),
.B(n_4748),
.Y(n_4875)
);

HB1xp67_ASAP7_75t_L g4876 ( 
.A(n_4774),
.Y(n_4876)
);

OAI22xp33_ASAP7_75t_L g4877 ( 
.A1(n_4738),
.A2(n_4706),
.B1(n_4718),
.B2(n_4724),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4851),
.Y(n_4878)
);

OR2x2_ASAP7_75t_L g4879 ( 
.A(n_4763),
.B(n_4643),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4843),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4754),
.B(n_4667),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4788),
.B(n_4605),
.Y(n_4882)
);

AND2x2_ASAP7_75t_L g4883 ( 
.A(n_4767),
.B(n_4667),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4865),
.Y(n_4884)
);

AND2x4_ASAP7_75t_L g4885 ( 
.A(n_4822),
.B(n_4703),
.Y(n_4885)
);

AND2x4_ASAP7_75t_L g4886 ( 
.A(n_4733),
.B(n_4744),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4820),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4830),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4819),
.B(n_4675),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4778),
.B(n_4688),
.Y(n_4890)
);

HB1xp67_ASAP7_75t_L g4891 ( 
.A(n_4772),
.Y(n_4891)
);

AOI22xp33_ASAP7_75t_L g4892 ( 
.A1(n_4737),
.A2(n_4742),
.B1(n_4732),
.B2(n_4735),
.Y(n_4892)
);

OR2x2_ASAP7_75t_L g4893 ( 
.A(n_4753),
.B(n_4643),
.Y(n_4893)
);

AND2x4_ASAP7_75t_L g4894 ( 
.A(n_4791),
.B(n_4703),
.Y(n_4894)
);

INVx2_ASAP7_75t_L g4895 ( 
.A(n_4859),
.Y(n_4895)
);

AND2x4_ASAP7_75t_L g4896 ( 
.A(n_4795),
.B(n_4631),
.Y(n_4896)
);

BUFx3_ASAP7_75t_L g4897 ( 
.A(n_4755),
.Y(n_4897)
);

AND2x4_ASAP7_75t_L g4898 ( 
.A(n_4814),
.B(n_4631),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4817),
.Y(n_4899)
);

HB1xp67_ASAP7_75t_L g4900 ( 
.A(n_4829),
.Y(n_4900)
);

INVx2_ASAP7_75t_L g4901 ( 
.A(n_4844),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4850),
.B(n_4688),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4787),
.B(n_4653),
.Y(n_4903)
);

INVx2_ASAP7_75t_SL g4904 ( 
.A(n_4855),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4833),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4841),
.B(n_4655),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4799),
.B(n_4663),
.Y(n_4907)
);

AND2x4_ASAP7_75t_L g4908 ( 
.A(n_4765),
.B(n_4632),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4818),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4848),
.Y(n_4910)
);

OR2x2_ASAP7_75t_L g4911 ( 
.A(n_4751),
.B(n_4623),
.Y(n_4911)
);

AND2x2_ASAP7_75t_L g4912 ( 
.A(n_4783),
.B(n_4702),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4853),
.Y(n_4913)
);

AND2x4_ASAP7_75t_L g4914 ( 
.A(n_4765),
.B(n_4632),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4740),
.B(n_4784),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4740),
.B(n_4607),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4740),
.B(n_4624),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4792),
.B(n_4635),
.Y(n_4918)
);

BUFx2_ASAP7_75t_L g4919 ( 
.A(n_4761),
.Y(n_4919)
);

INVx1_ASAP7_75t_SL g4920 ( 
.A(n_4863),
.Y(n_4920)
);

BUFx3_ASAP7_75t_L g4921 ( 
.A(n_4766),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_SL g4922 ( 
.A(n_4745),
.B(n_4718),
.Y(n_4922)
);

HB1xp67_ASAP7_75t_L g4923 ( 
.A(n_4769),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4771),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4835),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4779),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4847),
.Y(n_4927)
);

INVxp67_ASAP7_75t_L g4928 ( 
.A(n_4775),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4812),
.B(n_4663),
.Y(n_4929)
);

BUFx2_ASAP7_75t_L g4930 ( 
.A(n_4766),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4785),
.Y(n_4931)
);

AND2x2_ASAP7_75t_L g4932 ( 
.A(n_4800),
.B(n_4627),
.Y(n_4932)
);

AND2x2_ASAP7_75t_L g4933 ( 
.A(n_4838),
.B(n_4665),
.Y(n_4933)
);

AOI33xp33_ASAP7_75t_L g4934 ( 
.A1(n_4736),
.A2(n_4669),
.A3(n_4677),
.B1(n_340),
.B2(n_342),
.B3(n_343),
.Y(n_4934)
);

INVxp67_ASAP7_75t_SL g4935 ( 
.A(n_4864),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4807),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4856),
.B(n_4665),
.Y(n_4937)
);

AND2x2_ASAP7_75t_L g4938 ( 
.A(n_4826),
.B(n_4719),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4804),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4757),
.B(n_4599),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4780),
.Y(n_4941)
);

OR2x2_ASAP7_75t_L g4942 ( 
.A(n_4750),
.B(n_4649),
.Y(n_4942)
);

AND2x2_ASAP7_75t_L g4943 ( 
.A(n_4773),
.B(n_4726),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4834),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4747),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4747),
.Y(n_4946)
);

OR2x6_ASAP7_75t_L g4947 ( 
.A(n_4781),
.B(n_4716),
.Y(n_4947)
);

BUFx2_ASAP7_75t_L g4948 ( 
.A(n_4845),
.Y(n_4948)
);

INVx3_ASAP7_75t_L g4949 ( 
.A(n_4831),
.Y(n_4949)
);

INVx2_ASAP7_75t_L g4950 ( 
.A(n_4756),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4816),
.Y(n_4951)
);

AO21x2_ASAP7_75t_L g4952 ( 
.A1(n_4825),
.A2(n_4683),
.B(n_4649),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4816),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4790),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4854),
.Y(n_4955)
);

INVx2_ASAP7_75t_L g4956 ( 
.A(n_4762),
.Y(n_4956)
);

AND2x2_ASAP7_75t_L g4957 ( 
.A(n_4860),
.B(n_4726),
.Y(n_4957)
);

OR2x6_ASAP7_75t_L g4958 ( 
.A(n_4781),
.B(n_4796),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4806),
.Y(n_4959)
);

BUFx6f_ASAP7_75t_L g4960 ( 
.A(n_4802),
.Y(n_4960)
);

INVx2_ASAP7_75t_L g4961 ( 
.A(n_4852),
.Y(n_4961)
);

NOR2xp33_ASAP7_75t_L g4962 ( 
.A(n_4768),
.B(n_4633),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4770),
.Y(n_4963)
);

HB1xp67_ASAP7_75t_L g4964 ( 
.A(n_4777),
.Y(n_4964)
);

AND2x4_ASAP7_75t_L g4965 ( 
.A(n_4821),
.B(n_4614),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4739),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4823),
.B(n_4681),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4746),
.B(n_4681),
.Y(n_4968)
);

BUFx3_ASAP7_75t_L g4969 ( 
.A(n_4840),
.Y(n_4969)
);

NOR2x1_ASAP7_75t_L g4970 ( 
.A(n_4836),
.B(n_4628),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4866),
.B(n_4734),
.Y(n_4971)
);

NOR2xp33_ASAP7_75t_L g4972 ( 
.A(n_4872),
.B(n_4949),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4891),
.Y(n_4973)
);

AOI22xp33_ASAP7_75t_L g4974 ( 
.A1(n_4960),
.A2(n_4743),
.B1(n_4801),
.B2(n_4749),
.Y(n_4974)
);

INVx3_ASAP7_75t_L g4975 ( 
.A(n_4897),
.Y(n_4975)
);

OAI221xp5_ASAP7_75t_L g4976 ( 
.A1(n_4892),
.A2(n_4776),
.B1(n_4811),
.B2(n_4805),
.C(n_4741),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4964),
.B(n_4945),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4873),
.B(n_4803),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4930),
.B(n_4810),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4891),
.Y(n_4980)
);

AOI22xp33_ASAP7_75t_SL g4981 ( 
.A1(n_4935),
.A2(n_4815),
.B1(n_4764),
.B2(n_4832),
.Y(n_4981)
);

AO21x2_ASAP7_75t_L g4982 ( 
.A1(n_4868),
.A2(n_4794),
.B(n_4782),
.Y(n_4982)
);

AOI22xp5_ASAP7_75t_L g4983 ( 
.A1(n_4935),
.A2(n_4832),
.B1(n_4813),
.B2(n_4828),
.Y(n_4983)
);

OR2x2_ASAP7_75t_L g4984 ( 
.A(n_4911),
.B(n_4760),
.Y(n_4984)
);

OAI33xp33_ASAP7_75t_L g4985 ( 
.A1(n_4966),
.A2(n_4824),
.A3(n_4797),
.B1(n_4861),
.B2(n_4858),
.B3(n_4793),
.Y(n_4985)
);

AO21x2_ASAP7_75t_L g4986 ( 
.A1(n_4868),
.A2(n_4722),
.B(n_4793),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4964),
.B(n_4723),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4946),
.B(n_4923),
.Y(n_4988)
);

AO21x2_ASAP7_75t_L g4989 ( 
.A1(n_4922),
.A2(n_4610),
.B(n_4697),
.Y(n_4989)
);

OR2x2_ASAP7_75t_L g4990 ( 
.A(n_4893),
.B(n_4759),
.Y(n_4990)
);

INVx2_ASAP7_75t_L g4991 ( 
.A(n_4885),
.Y(n_4991)
);

OAI322xp33_ASAP7_75t_L g4992 ( 
.A1(n_4928),
.A2(n_4846),
.A3(n_4752),
.B1(n_343),
.B2(n_344),
.C1(n_346),
.C2(n_348),
.Y(n_4992)
);

INVx2_ASAP7_75t_L g4993 ( 
.A(n_4885),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4908),
.B(n_4798),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4900),
.Y(n_4995)
);

OAI33xp33_ASAP7_75t_L g4996 ( 
.A1(n_4928),
.A2(n_338),
.A3(n_339),
.B1(n_346),
.B2(n_348),
.B3(n_349),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4908),
.B(n_4827),
.Y(n_4997)
);

AND2x2_ASAP7_75t_L g4998 ( 
.A(n_4908),
.B(n_4723),
.Y(n_4998)
);

OAI22xp33_ASAP7_75t_L g4999 ( 
.A1(n_4958),
.A2(n_4628),
.B1(n_4752),
.B2(n_4758),
.Y(n_4999)
);

OAI22xp5_ASAP7_75t_L g5000 ( 
.A1(n_4892),
.A2(n_4789),
.B1(n_4837),
.B2(n_4849),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4914),
.B(n_4723),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_SL g5002 ( 
.A(n_4877),
.B(n_4731),
.Y(n_5002)
);

AOI221xp5_ASAP7_75t_L g5003 ( 
.A1(n_4960),
.A2(n_4954),
.B1(n_4922),
.B2(n_4951),
.C(n_4953),
.Y(n_5003)
);

NAND3xp33_ASAP7_75t_L g5004 ( 
.A(n_4960),
.B(n_4628),
.C(n_4608),
.Y(n_5004)
);

AOI22xp5_ASAP7_75t_SL g5005 ( 
.A1(n_4969),
.A2(n_4588),
.B1(n_350),
.B2(n_338),
.Y(n_5005)
);

AOI222xp33_ASAP7_75t_L g5006 ( 
.A1(n_4960),
.A2(n_4959),
.B1(n_4963),
.B2(n_4969),
.C1(n_4955),
.C2(n_4961),
.Y(n_5006)
);

OA21x2_ASAP7_75t_L g5007 ( 
.A1(n_4968),
.A2(n_4634),
.B(n_4630),
.Y(n_5007)
);

AOI221xp5_ASAP7_75t_L g5008 ( 
.A1(n_4959),
.A2(n_4963),
.B1(n_4962),
.B2(n_4877),
.C(n_4939),
.Y(n_5008)
);

AND2x2_ASAP7_75t_L g5009 ( 
.A(n_4914),
.B(n_4588),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4900),
.Y(n_5010)
);

OAI31xp33_ASAP7_75t_SL g5011 ( 
.A1(n_4970),
.A2(n_4588),
.A3(n_352),
.B(n_349),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4876),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4876),
.Y(n_5013)
);

BUFx3_ASAP7_75t_L g5014 ( 
.A(n_4872),
.Y(n_5014)
);

NAND3xp33_ASAP7_75t_L g5015 ( 
.A(n_4958),
.B(n_351),
.C(n_353),
.Y(n_5015)
);

AOI22xp5_ASAP7_75t_L g5016 ( 
.A1(n_4958),
.A2(n_4630),
.B1(n_356),
.B2(n_354),
.Y(n_5016)
);

OR2x2_ASAP7_75t_L g5017 ( 
.A(n_4923),
.B(n_354),
.Y(n_5017)
);

OAI221xp5_ASAP7_75t_SL g5018 ( 
.A1(n_4934),
.A2(n_355),
.B1(n_357),
.B2(n_358),
.C(n_359),
.Y(n_5018)
);

AOI221xp5_ASAP7_75t_L g5019 ( 
.A1(n_4962),
.A2(n_355),
.B1(n_358),
.B2(n_361),
.C(n_364),
.Y(n_5019)
);

HB1xp67_ASAP7_75t_L g5020 ( 
.A(n_4874),
.Y(n_5020)
);

OA21x2_ASAP7_75t_L g5021 ( 
.A1(n_4940),
.A2(n_361),
.B(n_364),
.Y(n_5021)
);

OAI21xp5_ASAP7_75t_L g5022 ( 
.A1(n_4934),
.A2(n_366),
.B(n_367),
.Y(n_5022)
);

NOR2xp33_ASAP7_75t_L g5023 ( 
.A(n_4949),
.B(n_367),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4867),
.Y(n_5024)
);

HB1xp67_ASAP7_75t_L g5025 ( 
.A(n_4874),
.Y(n_5025)
);

HB1xp67_ASAP7_75t_L g5026 ( 
.A(n_4933),
.Y(n_5026)
);

OA21x2_ASAP7_75t_L g5027 ( 
.A1(n_4885),
.A2(n_369),
.B(n_370),
.Y(n_5027)
);

AND2x2_ASAP7_75t_L g5028 ( 
.A(n_4914),
.B(n_4902),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4870),
.Y(n_5029)
);

OAI211xp5_ASAP7_75t_L g5030 ( 
.A1(n_4961),
.A2(n_4944),
.B(n_4941),
.C(n_4925),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4897),
.Y(n_5031)
);

AOI22xp33_ASAP7_75t_L g5032 ( 
.A1(n_4942),
.A2(n_369),
.B1(n_370),
.B2(n_372),
.Y(n_5032)
);

INVx2_ASAP7_75t_L g5033 ( 
.A(n_4915),
.Y(n_5033)
);

OAI22xp5_ASAP7_75t_L g5034 ( 
.A1(n_4947),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_5034)
);

OR2x2_ASAP7_75t_L g5035 ( 
.A(n_4882),
.B(n_373),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4878),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_4894),
.Y(n_5037)
);

NOR2xp33_ASAP7_75t_L g5038 ( 
.A(n_4949),
.B(n_374),
.Y(n_5038)
);

AOI211xp5_ASAP7_75t_L g5039 ( 
.A1(n_4929),
.A2(n_375),
.B(n_376),
.C(n_377),
.Y(n_5039)
);

INVx2_ASAP7_75t_L g5040 ( 
.A(n_4894),
.Y(n_5040)
);

INVx2_ASAP7_75t_L g5041 ( 
.A(n_5027),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4973),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4980),
.Y(n_5043)
);

NAND2x1_ASAP7_75t_L g5044 ( 
.A(n_5027),
.B(n_4894),
.Y(n_5044)
);

INVx2_ASAP7_75t_L g5045 ( 
.A(n_5014),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4975),
.B(n_4929),
.Y(n_5046)
);

INVx2_ASAP7_75t_L g5047 ( 
.A(n_4975),
.Y(n_5047)
);

AND2x2_ASAP7_75t_L g5048 ( 
.A(n_5028),
.B(n_4875),
.Y(n_5048)
);

HB1xp67_ASAP7_75t_L g5049 ( 
.A(n_5026),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4981),
.B(n_4925),
.Y(n_5050)
);

INVx2_ASAP7_75t_L g5051 ( 
.A(n_4991),
.Y(n_5051)
);

OR2x2_ASAP7_75t_L g5052 ( 
.A(n_4977),
.B(n_4880),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4995),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4993),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_5010),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_5020),
.Y(n_5056)
);

AND2x2_ASAP7_75t_L g5057 ( 
.A(n_5037),
.B(n_4952),
.Y(n_5057)
);

AND2x2_ASAP7_75t_L g5058 ( 
.A(n_5040),
.B(n_4952),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_5025),
.Y(n_5059)
);

BUFx2_ASAP7_75t_L g5060 ( 
.A(n_5031),
.Y(n_5060)
);

AND2x4_ASAP7_75t_L g5061 ( 
.A(n_5033),
.B(n_4886),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_5012),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_5013),
.Y(n_5063)
);

BUFx2_ASAP7_75t_L g5064 ( 
.A(n_4982),
.Y(n_5064)
);

OR2x2_ASAP7_75t_L g5065 ( 
.A(n_4977),
.B(n_4909),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_5024),
.Y(n_5066)
);

BUFx2_ASAP7_75t_L g5067 ( 
.A(n_4982),
.Y(n_5067)
);

BUFx2_ASAP7_75t_L g5068 ( 
.A(n_5021),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_5029),
.Y(n_5069)
);

AND2x2_ASAP7_75t_L g5070 ( 
.A(n_4971),
.B(n_4896),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_5036),
.Y(n_5071)
);

AND2x2_ASAP7_75t_L g5072 ( 
.A(n_4997),
.B(n_4896),
.Y(n_5072)
);

BUFx2_ASAP7_75t_L g5073 ( 
.A(n_5021),
.Y(n_5073)
);

INVx2_ASAP7_75t_L g5074 ( 
.A(n_4998),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_5001),
.B(n_4896),
.Y(n_5075)
);

INVx1_ASAP7_75t_SL g5076 ( 
.A(n_5017),
.Y(n_5076)
);

INVx2_ASAP7_75t_L g5077 ( 
.A(n_5009),
.Y(n_5077)
);

AND2x2_ASAP7_75t_L g5078 ( 
.A(n_4994),
.B(n_4898),
.Y(n_5078)
);

INVx2_ASAP7_75t_SL g5079 ( 
.A(n_4972),
.Y(n_5079)
);

AND2x2_ASAP7_75t_L g5080 ( 
.A(n_4978),
.B(n_4979),
.Y(n_5080)
);

BUFx2_ASAP7_75t_L g5081 ( 
.A(n_4988),
.Y(n_5081)
);

INVx1_ASAP7_75t_SL g5082 ( 
.A(n_4988),
.Y(n_5082)
);

OR2x2_ASAP7_75t_L g5083 ( 
.A(n_4987),
.B(n_4909),
.Y(n_5083)
);

AND2x2_ASAP7_75t_L g5084 ( 
.A(n_5011),
.B(n_4898),
.Y(n_5084)
);

OR2x2_ASAP7_75t_L g5085 ( 
.A(n_4987),
.B(n_4984),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_5049),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_5056),
.Y(n_5087)
);

OAI322xp33_ASAP7_75t_L g5088 ( 
.A1(n_5050),
.A2(n_4983),
.A3(n_4999),
.B1(n_4976),
.B2(n_5005),
.C1(n_5016),
.C2(n_5034),
.Y(n_5088)
);

NOR3xp33_ASAP7_75t_L g5089 ( 
.A(n_5079),
.B(n_5003),
.C(n_5030),
.Y(n_5089)
);

AND2x2_ASAP7_75t_SL g5090 ( 
.A(n_5064),
.B(n_5003),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_5084),
.B(n_5006),
.Y(n_5091)
);

OR2x2_ASAP7_75t_L g5092 ( 
.A(n_5076),
.B(n_4990),
.Y(n_5092)
);

NOR2xp33_ASAP7_75t_SL g5093 ( 
.A(n_5079),
.B(n_5018),
.Y(n_5093)
);

INVxp67_ASAP7_75t_SL g5094 ( 
.A(n_5044),
.Y(n_5094)
);

NAND3xp33_ASAP7_75t_L g5095 ( 
.A(n_5064),
.B(n_5011),
.C(n_5006),
.Y(n_5095)
);

OR2x2_ASAP7_75t_L g5096 ( 
.A(n_5068),
.B(n_5030),
.Y(n_5096)
);

OAI321xp33_ASAP7_75t_L g5097 ( 
.A1(n_5067),
.A2(n_5022),
.A3(n_4976),
.B1(n_5008),
.B2(n_4974),
.C(n_5039),
.Y(n_5097)
);

INVx2_ASAP7_75t_L g5098 ( 
.A(n_5067),
.Y(n_5098)
);

AOI33xp33_ASAP7_75t_L g5099 ( 
.A1(n_5082),
.A2(n_5008),
.A3(n_5019),
.B1(n_5032),
.B2(n_4985),
.B3(n_4927),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_5056),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_5060),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5059),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_5059),
.Y(n_5103)
);

BUFx2_ASAP7_75t_L g5104 ( 
.A(n_5060),
.Y(n_5104)
);

AND2x2_ASAP7_75t_L g5105 ( 
.A(n_5084),
.B(n_5048),
.Y(n_5105)
);

NOR2x1_ASAP7_75t_SL g5106 ( 
.A(n_5041),
.B(n_4947),
.Y(n_5106)
);

INVxp67_ASAP7_75t_L g5107 ( 
.A(n_5068),
.Y(n_5107)
);

INVx2_ASAP7_75t_SL g5108 ( 
.A(n_5061),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_5062),
.Y(n_5109)
);

NAND3xp33_ASAP7_75t_L g5110 ( 
.A(n_5073),
.B(n_5022),
.C(n_5015),
.Y(n_5110)
);

AND2x2_ASAP7_75t_L g5111 ( 
.A(n_5048),
.B(n_4904),
.Y(n_5111)
);

HB1xp67_ASAP7_75t_L g5112 ( 
.A(n_5044),
.Y(n_5112)
);

OAI22xp5_ASAP7_75t_L g5113 ( 
.A1(n_5073),
.A2(n_4947),
.B1(n_5004),
.B2(n_5034),
.Y(n_5113)
);

INVx2_ASAP7_75t_L g5114 ( 
.A(n_5047),
.Y(n_5114)
);

AOI22xp33_ASAP7_75t_L g5115 ( 
.A1(n_5080),
.A2(n_4992),
.B1(n_5019),
.B2(n_4996),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_5062),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_5104),
.Y(n_5117)
);

AOI32xp33_ASAP7_75t_L g5118 ( 
.A1(n_5091),
.A2(n_5041),
.A3(n_5046),
.B1(n_5081),
.B2(n_5080),
.Y(n_5118)
);

AOI22xp5_ASAP7_75t_L g5119 ( 
.A1(n_5095),
.A2(n_5041),
.B1(n_5081),
.B2(n_5000),
.Y(n_5119)
);

OAI21xp33_ASAP7_75t_L g5120 ( 
.A1(n_5093),
.A2(n_5046),
.B(n_5085),
.Y(n_5120)
);

AND2x4_ASAP7_75t_L g5121 ( 
.A(n_5108),
.B(n_5047),
.Y(n_5121)
);

OR2x2_ASAP7_75t_L g5122 ( 
.A(n_5092),
.B(n_5085),
.Y(n_5122)
);

AND2x4_ASAP7_75t_L g5123 ( 
.A(n_5108),
.B(n_5045),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_5101),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_5101),
.Y(n_5125)
);

BUFx2_ASAP7_75t_L g5126 ( 
.A(n_5094),
.Y(n_5126)
);

INVx2_ASAP7_75t_L g5127 ( 
.A(n_5111),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_L g5128 ( 
.A(n_5090),
.B(n_5051),
.Y(n_5128)
);

NOR2x1_ASAP7_75t_L g5129 ( 
.A(n_5096),
.B(n_5045),
.Y(n_5129)
);

AND2x2_ASAP7_75t_L g5130 ( 
.A(n_5105),
.B(n_5070),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_5098),
.Y(n_5131)
);

AND2x2_ASAP7_75t_L g5132 ( 
.A(n_5105),
.B(n_5070),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_5098),
.Y(n_5133)
);

OR2x2_ASAP7_75t_L g5134 ( 
.A(n_5086),
.B(n_5052),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_5091),
.B(n_5051),
.Y(n_5135)
);

AND2x2_ASAP7_75t_L g5136 ( 
.A(n_5111),
.B(n_5078),
.Y(n_5136)
);

AND2x2_ASAP7_75t_L g5137 ( 
.A(n_5106),
.B(n_5078),
.Y(n_5137)
);

NAND2xp5_ASAP7_75t_L g5138 ( 
.A(n_5090),
.B(n_5054),
.Y(n_5138)
);

AND2x4_ASAP7_75t_L g5139 ( 
.A(n_5121),
.B(n_5123),
.Y(n_5139)
);

BUFx3_ASAP7_75t_L g5140 ( 
.A(n_5123),
.Y(n_5140)
);

OR2x2_ASAP7_75t_L g5141 ( 
.A(n_5135),
.B(n_5096),
.Y(n_5141)
);

OR2x2_ASAP7_75t_L g5142 ( 
.A(n_5117),
.B(n_5110),
.Y(n_5142)
);

INVx1_ASAP7_75t_SL g5143 ( 
.A(n_5130),
.Y(n_5143)
);

AOI211xp5_ASAP7_75t_L g5144 ( 
.A1(n_5120),
.A2(n_5088),
.B(n_5097),
.C(n_5089),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5129),
.Y(n_5145)
);

AND2x2_ASAP7_75t_L g5146 ( 
.A(n_5132),
.B(n_5072),
.Y(n_5146)
);

AND2x2_ASAP7_75t_L g5147 ( 
.A(n_5136),
.B(n_5072),
.Y(n_5147)
);

NAND2x1p5_ASAP7_75t_L g5148 ( 
.A(n_5137),
.B(n_4871),
.Y(n_5148)
);

INVx1_ASAP7_75t_L g5149 ( 
.A(n_5126),
.Y(n_5149)
);

INVxp67_ASAP7_75t_L g5150 ( 
.A(n_5128),
.Y(n_5150)
);

AND2x4_ASAP7_75t_L g5151 ( 
.A(n_5121),
.B(n_5114),
.Y(n_5151)
);

OR2x2_ASAP7_75t_L g5152 ( 
.A(n_5122),
.B(n_5052),
.Y(n_5152)
);

NOR3xp33_ASAP7_75t_L g5153 ( 
.A(n_5120),
.B(n_5138),
.C(n_5128),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5138),
.Y(n_5154)
);

BUFx3_ASAP7_75t_L g5155 ( 
.A(n_5127),
.Y(n_5155)
);

OR2x2_ASAP7_75t_L g5156 ( 
.A(n_5134),
.B(n_5054),
.Y(n_5156)
);

OAI211xp5_ASAP7_75t_SL g5157 ( 
.A1(n_5119),
.A2(n_5099),
.B(n_5115),
.C(n_5107),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_5124),
.Y(n_5158)
);

NOR2xp67_ASAP7_75t_SL g5159 ( 
.A(n_5125),
.B(n_4871),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5131),
.Y(n_5160)
);

OR2x2_ASAP7_75t_L g5161 ( 
.A(n_5119),
.B(n_5065),
.Y(n_5161)
);

NOR2xp33_ASAP7_75t_L g5162 ( 
.A(n_5148),
.B(n_4948),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_5139),
.B(n_5118),
.Y(n_5163)
);

INVxp67_ASAP7_75t_SL g5164 ( 
.A(n_5140),
.Y(n_5164)
);

INVx2_ASAP7_75t_L g5165 ( 
.A(n_5139),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_5151),
.Y(n_5166)
);

INVx1_ASAP7_75t_SL g5167 ( 
.A(n_5152),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5146),
.B(n_5114),
.Y(n_5168)
);

AND2x2_ASAP7_75t_L g5169 ( 
.A(n_5147),
.B(n_5143),
.Y(n_5169)
);

O2A1O1Ixp33_ASAP7_75t_SL g5170 ( 
.A1(n_5144),
.A2(n_5112),
.B(n_4904),
.C(n_5113),
.Y(n_5170)
);

AND2x2_ASAP7_75t_L g5171 ( 
.A(n_5155),
.B(n_4919),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_L g5172 ( 
.A(n_5153),
.B(n_5115),
.Y(n_5172)
);

OAI31xp33_ASAP7_75t_L g5173 ( 
.A1(n_5157),
.A2(n_5023),
.A3(n_5038),
.B(n_5035),
.Y(n_5173)
);

OR2x2_ASAP7_75t_L g5174 ( 
.A(n_5141),
.B(n_5065),
.Y(n_5174)
);

AND2x4_ASAP7_75t_L g5175 ( 
.A(n_5151),
.B(n_5133),
.Y(n_5175)
);

INVx1_ASAP7_75t_SL g5176 ( 
.A(n_5145),
.Y(n_5176)
);

NAND2xp5_ASAP7_75t_L g5177 ( 
.A(n_5149),
.B(n_5099),
.Y(n_5177)
);

HB1xp67_ASAP7_75t_L g5178 ( 
.A(n_5175),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_5175),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_5164),
.B(n_5149),
.Y(n_5180)
);

OR2x2_ASAP7_75t_L g5181 ( 
.A(n_5165),
.B(n_5161),
.Y(n_5181)
);

INVxp67_ASAP7_75t_L g5182 ( 
.A(n_5162),
.Y(n_5182)
);

OR2x2_ASAP7_75t_L g5183 ( 
.A(n_5167),
.B(n_5142),
.Y(n_5183)
);

HB1xp67_ASAP7_75t_L g5184 ( 
.A(n_5166),
.Y(n_5184)
);

AND2x2_ASAP7_75t_L g5185 ( 
.A(n_5171),
.B(n_5159),
.Y(n_5185)
);

AOI22xp33_ASAP7_75t_SL g5186 ( 
.A1(n_5172),
.A2(n_5154),
.B1(n_5150),
.B2(n_5058),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_5169),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_5168),
.B(n_5154),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_5178),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_5181),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_5184),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5179),
.Y(n_5192)
);

NAND2xp5_ASAP7_75t_SL g5193 ( 
.A(n_5183),
.B(n_5173),
.Y(n_5193)
);

INVx2_ASAP7_75t_L g5194 ( 
.A(n_5185),
.Y(n_5194)
);

OAI21xp33_ASAP7_75t_SL g5195 ( 
.A1(n_5188),
.A2(n_5173),
.B(n_5177),
.Y(n_5195)
);

INVx2_ASAP7_75t_L g5196 ( 
.A(n_5187),
.Y(n_5196)
);

OR2x2_ASAP7_75t_L g5197 ( 
.A(n_5180),
.B(n_5156),
.Y(n_5197)
);

OR2x2_ASAP7_75t_L g5198 ( 
.A(n_5188),
.B(n_5174),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_5186),
.B(n_5176),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_5182),
.Y(n_5200)
);

AOI221xp5_ASAP7_75t_L g5201 ( 
.A1(n_5186),
.A2(n_5170),
.B1(n_5176),
.B2(n_5163),
.C(n_5102),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_5178),
.Y(n_5202)
);

OR2x2_ASAP7_75t_L g5203 ( 
.A(n_5189),
.B(n_5158),
.Y(n_5203)
);

AND3x2_ASAP7_75t_L g5204 ( 
.A(n_5189),
.B(n_5202),
.C(n_5191),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_5194),
.B(n_5192),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_5198),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_5197),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_5190),
.Y(n_5208)
);

INVxp67_ASAP7_75t_SL g5209 ( 
.A(n_5193),
.Y(n_5209)
);

AOI31xp33_ASAP7_75t_SL g5210 ( 
.A1(n_5201),
.A2(n_5074),
.A3(n_5077),
.B(n_5083),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_5196),
.B(n_5160),
.Y(n_5211)
);

OAI22xp5_ASAP7_75t_L g5212 ( 
.A1(n_5199),
.A2(n_5063),
.B1(n_5061),
.B2(n_5074),
.Y(n_5212)
);

AND2x2_ASAP7_75t_L g5213 ( 
.A(n_5200),
.B(n_5087),
.Y(n_5213)
);

OAI21xp33_ASAP7_75t_SL g5214 ( 
.A1(n_5209),
.A2(n_5058),
.B(n_5057),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5206),
.B(n_5100),
.Y(n_5215)
);

O2A1O1Ixp33_ASAP7_75t_SL g5216 ( 
.A1(n_5203),
.A2(n_5103),
.B(n_5116),
.C(n_5109),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_5204),
.B(n_5195),
.Y(n_5217)
);

OR2x2_ASAP7_75t_L g5218 ( 
.A(n_5205),
.B(n_5063),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_5212),
.Y(n_5219)
);

INVx2_ASAP7_75t_SL g5220 ( 
.A(n_5213),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_5208),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_5210),
.Y(n_5222)
);

NAND2xp5_ASAP7_75t_L g5223 ( 
.A(n_5215),
.B(n_5207),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_5217),
.Y(n_5224)
);

A2O1A1Ixp33_ASAP7_75t_L g5225 ( 
.A1(n_5214),
.A2(n_5211),
.B(n_5042),
.C(n_5053),
.Y(n_5225)
);

XNOR2x1_ASAP7_75t_L g5226 ( 
.A(n_5222),
.B(n_4920),
.Y(n_5226)
);

NOR2xp33_ASAP7_75t_L g5227 ( 
.A(n_5220),
.B(n_5042),
.Y(n_5227)
);

NOR2x1_ASAP7_75t_L g5228 ( 
.A(n_5218),
.B(n_5043),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_5216),
.Y(n_5229)
);

OR2x2_ASAP7_75t_L g5230 ( 
.A(n_5219),
.B(n_5043),
.Y(n_5230)
);

OAI22xp5_ASAP7_75t_L g5231 ( 
.A1(n_5221),
.A2(n_5055),
.B1(n_5053),
.B2(n_5066),
.Y(n_5231)
);

CKINVDCx14_ASAP7_75t_R g5232 ( 
.A(n_5215),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5217),
.Y(n_5233)
);

AND2x2_ASAP7_75t_L g5234 ( 
.A(n_5222),
.B(n_5061),
.Y(n_5234)
);

NAND3xp33_ASAP7_75t_L g5235 ( 
.A(n_5217),
.B(n_5055),
.C(n_5066),
.Y(n_5235)
);

AOI22xp5_ASAP7_75t_L g5236 ( 
.A1(n_5222),
.A2(n_5061),
.B1(n_5071),
.B2(n_5069),
.Y(n_5236)
);

INVxp67_ASAP7_75t_L g5237 ( 
.A(n_5217),
.Y(n_5237)
);

AOI22xp5_ASAP7_75t_L g5238 ( 
.A1(n_5222),
.A2(n_5071),
.B1(n_5069),
.B2(n_5057),
.Y(n_5238)
);

AOI22xp33_ASAP7_75t_L g5239 ( 
.A1(n_5222),
.A2(n_5077),
.B1(n_5083),
.B2(n_5075),
.Y(n_5239)
);

NOR2xp33_ASAP7_75t_L g5240 ( 
.A(n_5232),
.B(n_4950),
.Y(n_5240)
);

NOR2x1_ASAP7_75t_L g5241 ( 
.A(n_5229),
.B(n_4950),
.Y(n_5241)
);

A2O1A1Ixp33_ASAP7_75t_L g5242 ( 
.A1(n_5227),
.A2(n_4956),
.B(n_5075),
.C(n_4921),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5234),
.Y(n_5243)
);

NOR2x1_ASAP7_75t_L g5244 ( 
.A(n_5223),
.B(n_4956),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5226),
.Y(n_5245)
);

OR2x2_ASAP7_75t_L g5246 ( 
.A(n_5230),
.B(n_4924),
.Y(n_5246)
);

NAND3xp33_ASAP7_75t_SL g5247 ( 
.A(n_5238),
.B(n_5002),
.C(n_4943),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5228),
.Y(n_5248)
);

NOR3xp33_ASAP7_75t_L g5249 ( 
.A(n_5237),
.B(n_4913),
.C(n_4910),
.Y(n_5249)
);

AO22x2_ASAP7_75t_L g5250 ( 
.A1(n_5224),
.A2(n_4931),
.B1(n_5000),
.B2(n_4888),
.Y(n_5250)
);

NOR2x1p5_ASAP7_75t_L g5251 ( 
.A(n_5233),
.B(n_4921),
.Y(n_5251)
);

HB1xp67_ASAP7_75t_L g5252 ( 
.A(n_5231),
.Y(n_5252)
);

NOR2xp33_ASAP7_75t_L g5253 ( 
.A(n_5236),
.B(n_4869),
.Y(n_5253)
);

NOR2xp33_ASAP7_75t_L g5254 ( 
.A(n_5235),
.B(n_4869),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_5239),
.B(n_4887),
.Y(n_5255)
);

AND2x4_ASAP7_75t_L g5256 ( 
.A(n_5225),
.B(n_4912),
.Y(n_5256)
);

NAND3xp33_ASAP7_75t_L g5257 ( 
.A(n_5226),
.B(n_5007),
.C(n_4936),
.Y(n_5257)
);

NOR3xp33_ASAP7_75t_L g5258 ( 
.A(n_5232),
.B(n_4957),
.C(n_4926),
.Y(n_5258)
);

NAND3xp33_ASAP7_75t_SL g5259 ( 
.A(n_5229),
.B(n_4937),
.C(n_4905),
.Y(n_5259)
);

NOR2xp33_ASAP7_75t_SL g5260 ( 
.A(n_5234),
.B(n_4869),
.Y(n_5260)
);

NAND2x1_ASAP7_75t_SL g5261 ( 
.A(n_5228),
.B(n_5007),
.Y(n_5261)
);

NOR3x1_ASAP7_75t_L g5262 ( 
.A(n_5235),
.B(n_4899),
.C(n_4918),
.Y(n_5262)
);

NAND3xp33_ASAP7_75t_L g5263 ( 
.A(n_5226),
.B(n_4886),
.C(n_4884),
.Y(n_5263)
);

INVx2_ASAP7_75t_L g5264 ( 
.A(n_5226),
.Y(n_5264)
);

OAI21xp33_ASAP7_75t_L g5265 ( 
.A1(n_5260),
.A2(n_4886),
.B(n_4938),
.Y(n_5265)
);

AOI22xp5_ASAP7_75t_L g5266 ( 
.A1(n_5258),
.A2(n_4986),
.B1(n_4989),
.B2(n_4898),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_L g5267 ( 
.A(n_5256),
.B(n_4986),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_5241),
.Y(n_5268)
);

NOR3xp33_ASAP7_75t_L g5269 ( 
.A(n_5243),
.B(n_5245),
.C(n_5264),
.Y(n_5269)
);

OAI21xp33_ASAP7_75t_L g5270 ( 
.A1(n_5253),
.A2(n_4889),
.B(n_4917),
.Y(n_5270)
);

O2A1O1Ixp33_ASAP7_75t_L g5271 ( 
.A1(n_5248),
.A2(n_4989),
.B(n_4895),
.C(n_381),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_5250),
.Y(n_5272)
);

NOR2xp33_ASAP7_75t_L g5273 ( 
.A(n_5259),
.B(n_4895),
.Y(n_5273)
);

AOI21xp5_ASAP7_75t_L g5274 ( 
.A1(n_5240),
.A2(n_4901),
.B(n_4916),
.Y(n_5274)
);

OAI221xp5_ASAP7_75t_L g5275 ( 
.A1(n_5242),
.A2(n_4901),
.B1(n_4879),
.B2(n_4967),
.C(n_4890),
.Y(n_5275)
);

OAI31xp33_ASAP7_75t_L g5276 ( 
.A1(n_5250),
.A2(n_5251),
.A3(n_5254),
.B(n_5257),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_SL g5277 ( 
.A(n_5244),
.B(n_5255),
.Y(n_5277)
);

INVx1_ASAP7_75t_SL g5278 ( 
.A(n_5246),
.Y(n_5278)
);

INVx2_ASAP7_75t_L g5279 ( 
.A(n_5261),
.Y(n_5279)
);

AOI321xp33_ASAP7_75t_L g5280 ( 
.A1(n_5249),
.A2(n_5247),
.A3(n_5252),
.B1(n_5263),
.B2(n_5262),
.C(n_4965),
.Y(n_5280)
);

O2A1O1Ixp33_ASAP7_75t_L g5281 ( 
.A1(n_5248),
.A2(n_376),
.B(n_379),
.C(n_382),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5256),
.Y(n_5282)
);

AOI21xp5_ASAP7_75t_L g5283 ( 
.A1(n_5240),
.A2(n_4932),
.B(n_4903),
.Y(n_5283)
);

O2A1O1Ixp33_ASAP7_75t_L g5284 ( 
.A1(n_5248),
.A2(n_384),
.B(n_388),
.C(n_390),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5256),
.Y(n_5285)
);

AO22x2_ASAP7_75t_L g5286 ( 
.A1(n_5248),
.A2(n_4907),
.B1(n_4906),
.B2(n_4883),
.Y(n_5286)
);

INVx2_ASAP7_75t_SL g5287 ( 
.A(n_5251),
.Y(n_5287)
);

INVxp67_ASAP7_75t_SL g5288 ( 
.A(n_5241),
.Y(n_5288)
);

AOI21xp5_ASAP7_75t_L g5289 ( 
.A1(n_5240),
.A2(n_4907),
.B(n_4881),
.Y(n_5289)
);

AOI221xp5_ASAP7_75t_L g5290 ( 
.A1(n_5259),
.A2(n_4965),
.B1(n_4906),
.B2(n_390),
.C(n_391),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_5256),
.Y(n_5291)
);

O2A1O1Ixp33_ASAP7_75t_L g5292 ( 
.A1(n_5288),
.A2(n_384),
.B(n_388),
.C(n_391),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5267),
.Y(n_5293)
);

AND2x2_ASAP7_75t_L g5294 ( 
.A(n_5282),
.B(n_4965),
.Y(n_5294)
);

NOR2xp67_ASAP7_75t_L g5295 ( 
.A(n_5268),
.B(n_393),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5272),
.Y(n_5296)
);

NOR2x1_ASAP7_75t_L g5297 ( 
.A(n_5279),
.B(n_393),
.Y(n_5297)
);

NOR2xp33_ASAP7_75t_L g5298 ( 
.A(n_5285),
.B(n_394),
.Y(n_5298)
);

NOR4xp75_ASAP7_75t_L g5299 ( 
.A(n_5277),
.B(n_395),
.C(n_397),
.D(n_398),
.Y(n_5299)
);

NOR3xp33_ASAP7_75t_L g5300 ( 
.A(n_5269),
.B(n_398),
.C(n_399),
.Y(n_5300)
);

NAND3xp33_ASAP7_75t_L g5301 ( 
.A(n_5276),
.B(n_401),
.C(n_402),
.Y(n_5301)
);

NOR2x1_ASAP7_75t_L g5302 ( 
.A(n_5281),
.B(n_401),
.Y(n_5302)
);

NAND3x1_ASAP7_75t_L g5303 ( 
.A(n_5291),
.B(n_402),
.C(n_403),
.Y(n_5303)
);

OAI21xp5_ASAP7_75t_L g5304 ( 
.A1(n_5290),
.A2(n_403),
.B(n_404),
.Y(n_5304)
);

NAND4xp75_ASAP7_75t_L g5305 ( 
.A(n_5287),
.B(n_404),
.C(n_408),
.D(n_409),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5265),
.B(n_408),
.Y(n_5306)
);

NOR3x1_ASAP7_75t_L g5307 ( 
.A(n_5280),
.B(n_410),
.C(n_411),
.Y(n_5307)
);

NOR3xp33_ASAP7_75t_L g5308 ( 
.A(n_5278),
.B(n_411),
.C(n_413),
.Y(n_5308)
);

NOR2x1_ASAP7_75t_L g5309 ( 
.A(n_5284),
.B(n_413),
.Y(n_5309)
);

NOR3xp33_ASAP7_75t_L g5310 ( 
.A(n_5273),
.B(n_414),
.C(n_415),
.Y(n_5310)
);

NAND3xp33_ASAP7_75t_L g5311 ( 
.A(n_5271),
.B(n_414),
.C(n_416),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_5283),
.B(n_419),
.Y(n_5312)
);

OAI211xp5_ASAP7_75t_L g5313 ( 
.A1(n_5270),
.A2(n_420),
.B(n_422),
.C(n_423),
.Y(n_5313)
);

NOR3xp33_ASAP7_75t_L g5314 ( 
.A(n_5274),
.B(n_423),
.C(n_424),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5289),
.B(n_425),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_5303),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_5294),
.Y(n_5317)
);

OAI22xp5_ASAP7_75t_SL g5318 ( 
.A1(n_5311),
.A2(n_5266),
.B1(n_5275),
.B2(n_5286),
.Y(n_5318)
);

AOI22xp5_ASAP7_75t_L g5319 ( 
.A1(n_5300),
.A2(n_5286),
.B1(n_428),
.B2(n_430),
.Y(n_5319)
);

AOI221xp5_ASAP7_75t_L g5320 ( 
.A1(n_5296),
.A2(n_427),
.B1(n_428),
.B2(n_431),
.C(n_432),
.Y(n_5320)
);

OR2x2_ASAP7_75t_L g5321 ( 
.A(n_5306),
.B(n_431),
.Y(n_5321)
);

XNOR2xp5_ASAP7_75t_L g5322 ( 
.A(n_5299),
.B(n_432),
.Y(n_5322)
);

OAI211xp5_ASAP7_75t_SL g5323 ( 
.A1(n_5304),
.A2(n_433),
.B(n_434),
.C(n_436),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_5297),
.Y(n_5324)
);

NAND4xp25_ASAP7_75t_L g5325 ( 
.A(n_5307),
.B(n_434),
.C(n_436),
.D(n_437),
.Y(n_5325)
);

OAI211xp5_ASAP7_75t_L g5326 ( 
.A1(n_5313),
.A2(n_5301),
.B(n_5292),
.C(n_5295),
.Y(n_5326)
);

NOR2x1_ASAP7_75t_L g5327 ( 
.A(n_5305),
.B(n_437),
.Y(n_5327)
);

AOI211xp5_ASAP7_75t_L g5328 ( 
.A1(n_5314),
.A2(n_438),
.B(n_439),
.C(n_440),
.Y(n_5328)
);

XNOR2x1_ASAP7_75t_L g5329 ( 
.A(n_5302),
.B(n_438),
.Y(n_5329)
);

NAND4xp25_ASAP7_75t_L g5330 ( 
.A(n_5310),
.B(n_439),
.C(n_440),
.D(n_442),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_5298),
.B(n_442),
.Y(n_5331)
);

AOI221xp5_ASAP7_75t_L g5332 ( 
.A1(n_5293),
.A2(n_443),
.B1(n_444),
.B2(n_445),
.C(n_446),
.Y(n_5332)
);

AOI21xp33_ASAP7_75t_SL g5333 ( 
.A1(n_5308),
.A2(n_444),
.B(n_447),
.Y(n_5333)
);

INVx2_ASAP7_75t_L g5334 ( 
.A(n_5321),
.Y(n_5334)
);

NOR3xp33_ASAP7_75t_L g5335 ( 
.A(n_5317),
.B(n_5312),
.C(n_5315),
.Y(n_5335)
);

NOR3xp33_ASAP7_75t_L g5336 ( 
.A(n_5331),
.B(n_5309),
.C(n_449),
.Y(n_5336)
);

NAND4xp25_ASAP7_75t_L g5337 ( 
.A(n_5325),
.B(n_447),
.C(n_450),
.D(n_458),
.Y(n_5337)
);

NOR2x1_ASAP7_75t_L g5338 ( 
.A(n_5316),
.B(n_459),
.Y(n_5338)
);

NAND5xp2_ASAP7_75t_L g5339 ( 
.A(n_5326),
.B(n_463),
.C(n_468),
.D(n_472),
.E(n_474),
.Y(n_5339)
);

BUFx2_ASAP7_75t_L g5340 ( 
.A(n_5327),
.Y(n_5340)
);

OAI22xp5_ASAP7_75t_L g5341 ( 
.A1(n_5319),
.A2(n_2167),
.B1(n_2259),
.B2(n_2257),
.Y(n_5341)
);

NOR3x1_ASAP7_75t_L g5342 ( 
.A(n_5330),
.B(n_476),
.C(n_477),
.Y(n_5342)
);

CKINVDCx5p33_ASAP7_75t_R g5343 ( 
.A(n_5324),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_5322),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_5329),
.Y(n_5345)
);

OR2x2_ASAP7_75t_L g5346 ( 
.A(n_5333),
.B(n_478),
.Y(n_5346)
);

INVx2_ASAP7_75t_L g5347 ( 
.A(n_5318),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5328),
.Y(n_5348)
);

AOI211xp5_ASAP7_75t_L g5349 ( 
.A1(n_5323),
.A2(n_479),
.B(n_483),
.C(n_484),
.Y(n_5349)
);

NOR3xp33_ASAP7_75t_L g5350 ( 
.A(n_5347),
.B(n_5332),
.C(n_5320),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_5338),
.B(n_486),
.Y(n_5351)
);

INVx2_ASAP7_75t_L g5352 ( 
.A(n_5346),
.Y(n_5352)
);

INVxp67_ASAP7_75t_L g5353 ( 
.A(n_5340),
.Y(n_5353)
);

NAND3xp33_ASAP7_75t_L g5354 ( 
.A(n_5336),
.B(n_2167),
.C(n_2259),
.Y(n_5354)
);

NAND5xp2_ASAP7_75t_L g5355 ( 
.A(n_5335),
.B(n_489),
.C(n_491),
.D(n_492),
.E(n_493),
.Y(n_5355)
);

OAI221xp5_ASAP7_75t_L g5356 ( 
.A1(n_5337),
.A2(n_494),
.B1(n_495),
.B2(n_496),
.C(n_498),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5344),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_5343),
.Y(n_5358)
);

OAI221xp5_ASAP7_75t_L g5359 ( 
.A1(n_5349),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.C(n_502),
.Y(n_5359)
);

OAI22xp5_ASAP7_75t_L g5360 ( 
.A1(n_5345),
.A2(n_2167),
.B1(n_2259),
.B2(n_2257),
.Y(n_5360)
);

AOI21xp33_ASAP7_75t_SL g5361 ( 
.A1(n_5348),
.A2(n_505),
.B(n_506),
.Y(n_5361)
);

NAND2xp5_ASAP7_75t_SL g5362 ( 
.A(n_5334),
.B(n_2117),
.Y(n_5362)
);

NOR3xp33_ASAP7_75t_L g5363 ( 
.A(n_5341),
.B(n_508),
.C(n_509),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5342),
.Y(n_5364)
);

NOR3xp33_ASAP7_75t_L g5365 ( 
.A(n_5339),
.B(n_510),
.C(n_512),
.Y(n_5365)
);

OAI22x1_ASAP7_75t_L g5366 ( 
.A1(n_5340),
.A2(n_514),
.B1(n_516),
.B2(n_517),
.Y(n_5366)
);

AOI22x1_ASAP7_75t_L g5367 ( 
.A1(n_5357),
.A2(n_519),
.B1(n_522),
.B2(n_524),
.Y(n_5367)
);

AOI21xp5_ASAP7_75t_L g5368 ( 
.A1(n_5353),
.A2(n_1624),
.B(n_1634),
.Y(n_5368)
);

BUFx2_ASAP7_75t_L g5369 ( 
.A(n_5351),
.Y(n_5369)
);

A2O1A1Ixp33_ASAP7_75t_L g5370 ( 
.A1(n_5358),
.A2(n_525),
.B(n_526),
.C(n_529),
.Y(n_5370)
);

XOR2xp5_ASAP7_75t_L g5371 ( 
.A(n_5364),
.B(n_532),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_5365),
.Y(n_5372)
);

AOI221xp5_ASAP7_75t_L g5373 ( 
.A1(n_5350),
.A2(n_2173),
.B1(n_2259),
.B2(n_2257),
.C(n_2252),
.Y(n_5373)
);

AND2x4_ASAP7_75t_L g5374 ( 
.A(n_5352),
.B(n_537),
.Y(n_5374)
);

INVx2_ASAP7_75t_L g5375 ( 
.A(n_5366),
.Y(n_5375)
);

INVxp67_ASAP7_75t_L g5376 ( 
.A(n_5356),
.Y(n_5376)
);

NAND4xp25_ASAP7_75t_L g5377 ( 
.A(n_5359),
.B(n_5363),
.C(n_5355),
.D(n_5354),
.Y(n_5377)
);

NAND5xp2_ASAP7_75t_L g5378 ( 
.A(n_5361),
.B(n_538),
.C(n_539),
.D(n_540),
.E(n_541),
.Y(n_5378)
);

BUFx6f_ASAP7_75t_L g5379 ( 
.A(n_5362),
.Y(n_5379)
);

OR4x1_ASAP7_75t_L g5380 ( 
.A(n_5372),
.B(n_5360),
.C(n_545),
.D(n_546),
.Y(n_5380)
);

INVx2_ASAP7_75t_SL g5381 ( 
.A(n_5374),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_5375),
.Y(n_5382)
);

CKINVDCx20_ASAP7_75t_R g5383 ( 
.A(n_5369),
.Y(n_5383)
);

NAND2xp5_ASAP7_75t_L g5384 ( 
.A(n_5371),
.B(n_542),
.Y(n_5384)
);

OAI22xp5_ASAP7_75t_L g5385 ( 
.A1(n_5376),
.A2(n_5379),
.B1(n_5373),
.B2(n_5367),
.Y(n_5385)
);

AND3x4_ASAP7_75t_L g5386 ( 
.A(n_5377),
.B(n_548),
.C(n_549),
.Y(n_5386)
);

XNOR2xp5_ASAP7_75t_L g5387 ( 
.A(n_5383),
.B(n_5368),
.Y(n_5387)
);

INVx2_ASAP7_75t_L g5388 ( 
.A(n_5380),
.Y(n_5388)
);

XNOR2xp5_ASAP7_75t_L g5389 ( 
.A(n_5382),
.B(n_5378),
.Y(n_5389)
);

XOR2x1_ASAP7_75t_L g5390 ( 
.A(n_5381),
.B(n_5379),
.Y(n_5390)
);

INVx2_ASAP7_75t_L g5391 ( 
.A(n_5386),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5384),
.Y(n_5392)
);

HB1xp67_ASAP7_75t_L g5393 ( 
.A(n_5385),
.Y(n_5393)
);

OAI22xp5_ASAP7_75t_SL g5394 ( 
.A1(n_5388),
.A2(n_5370),
.B1(n_554),
.B2(n_555),
.Y(n_5394)
);

INVx4_ASAP7_75t_L g5395 ( 
.A(n_5393),
.Y(n_5395)
);

AOI21xp33_ASAP7_75t_L g5396 ( 
.A1(n_5389),
.A2(n_552),
.B(n_556),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5391),
.Y(n_5397)
);

NAND4xp25_ASAP7_75t_L g5398 ( 
.A(n_5392),
.B(n_561),
.C(n_562),
.D(n_566),
.Y(n_5398)
);

XNOR2xp5_ASAP7_75t_L g5399 ( 
.A(n_5390),
.B(n_5387),
.Y(n_5399)
);

CKINVDCx20_ASAP7_75t_R g5400 ( 
.A(n_5399),
.Y(n_5400)
);

OAI22xp5_ASAP7_75t_SL g5401 ( 
.A1(n_5395),
.A2(n_567),
.B1(n_568),
.B2(n_569),
.Y(n_5401)
);

OAI22xp5_ASAP7_75t_L g5402 ( 
.A1(n_5397),
.A2(n_572),
.B1(n_575),
.B2(n_578),
.Y(n_5402)
);

AOI22xp5_ASAP7_75t_L g5403 ( 
.A1(n_5394),
.A2(n_5398),
.B1(n_5396),
.B2(n_2173),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_5399),
.Y(n_5404)
);

NOR3xp33_ASAP7_75t_L g5405 ( 
.A(n_5404),
.B(n_579),
.C(n_581),
.Y(n_5405)
);

XNOR2xp5_ASAP7_75t_L g5406 ( 
.A(n_5400),
.B(n_583),
.Y(n_5406)
);

INVx1_ASAP7_75t_L g5407 ( 
.A(n_5403),
.Y(n_5407)
);

HB1xp67_ASAP7_75t_L g5408 ( 
.A(n_5401),
.Y(n_5408)
);

NAND2xp5_ASAP7_75t_L g5409 ( 
.A(n_5408),
.B(n_5402),
.Y(n_5409)
);

NAND3xp33_ASAP7_75t_L g5410 ( 
.A(n_5407),
.B(n_2173),
.C(n_2257),
.Y(n_5410)
);

AOI21xp33_ASAP7_75t_L g5411 ( 
.A1(n_5406),
.A2(n_584),
.B(n_587),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_5405),
.Y(n_5412)
);

OAI21xp5_ASAP7_75t_L g5413 ( 
.A1(n_5408),
.A2(n_588),
.B(n_591),
.Y(n_5413)
);

AOI21xp5_ASAP7_75t_L g5414 ( 
.A1(n_5409),
.A2(n_1662),
.B(n_1639),
.Y(n_5414)
);

OAI21xp5_ASAP7_75t_L g5415 ( 
.A1(n_5412),
.A2(n_592),
.B(n_594),
.Y(n_5415)
);

AOI21x1_ASAP7_75t_L g5416 ( 
.A1(n_5410),
.A2(n_595),
.B(n_600),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_5413),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5411),
.Y(n_5418)
);

AOI22xp33_ASAP7_75t_L g5419 ( 
.A1(n_5412),
.A2(n_2150),
.B1(n_2252),
.B2(n_2240),
.Y(n_5419)
);

AOI222xp33_ASAP7_75t_L g5420 ( 
.A1(n_5412),
.A2(n_601),
.B1(n_602),
.B2(n_603),
.C1(n_604),
.C2(n_606),
.Y(n_5420)
);

OAI22xp5_ASAP7_75t_L g5421 ( 
.A1(n_5409),
.A2(n_609),
.B1(n_611),
.B2(n_613),
.Y(n_5421)
);

AOI222xp33_ASAP7_75t_L g5422 ( 
.A1(n_5412),
.A2(n_614),
.B1(n_615),
.B2(n_616),
.C1(n_617),
.C2(n_618),
.Y(n_5422)
);

BUFx2_ASAP7_75t_L g5423 ( 
.A(n_5412),
.Y(n_5423)
);

OAI21x1_ASAP7_75t_L g5424 ( 
.A1(n_5414),
.A2(n_620),
.B(n_623),
.Y(n_5424)
);

OAI21xp33_ASAP7_75t_L g5425 ( 
.A1(n_5417),
.A2(n_2150),
.B(n_2252),
.Y(n_5425)
);

AO21x2_ASAP7_75t_L g5426 ( 
.A1(n_5418),
.A2(n_627),
.B(n_631),
.Y(n_5426)
);

AOI22xp33_ASAP7_75t_SL g5427 ( 
.A1(n_5423),
.A2(n_2173),
.B1(n_2205),
.B2(n_2222),
.Y(n_5427)
);

AOI21xp5_ASAP7_75t_L g5428 ( 
.A1(n_5419),
.A2(n_1634),
.B(n_1624),
.Y(n_5428)
);

AOI21xp5_ASAP7_75t_L g5429 ( 
.A1(n_5415),
.A2(n_1634),
.B(n_1624),
.Y(n_5429)
);

OAI21xp5_ASAP7_75t_SL g5430 ( 
.A1(n_5416),
.A2(n_634),
.B(n_635),
.Y(n_5430)
);

NAND2xp5_ASAP7_75t_L g5431 ( 
.A(n_5422),
.B(n_637),
.Y(n_5431)
);

AOI21xp5_ASAP7_75t_L g5432 ( 
.A1(n_5421),
.A2(n_1639),
.B(n_1649),
.Y(n_5432)
);

NAND2xp5_ASAP7_75t_L g5433 ( 
.A(n_5420),
.B(n_640),
.Y(n_5433)
);

NOR2xp67_ASAP7_75t_SL g5434 ( 
.A(n_5431),
.B(n_1649),
.Y(n_5434)
);

NAND2xp5_ASAP7_75t_L g5435 ( 
.A(n_5433),
.B(n_642),
.Y(n_5435)
);

XNOR2xp5_ASAP7_75t_L g5436 ( 
.A(n_5432),
.B(n_645),
.Y(n_5436)
);

AO21x2_ASAP7_75t_L g5437 ( 
.A1(n_5429),
.A2(n_1653),
.B(n_1666),
.Y(n_5437)
);

OAI22xp5_ASAP7_75t_L g5438 ( 
.A1(n_5430),
.A2(n_649),
.B1(n_2252),
.B2(n_2240),
.Y(n_5438)
);

XNOR2xp5_ASAP7_75t_L g5439 ( 
.A(n_5427),
.B(n_2205),
.Y(n_5439)
);

XNOR2xp5_ASAP7_75t_L g5440 ( 
.A(n_5424),
.B(n_2205),
.Y(n_5440)
);

OA21x2_ASAP7_75t_L g5441 ( 
.A1(n_5428),
.A2(n_2205),
.B(n_2240),
.Y(n_5441)
);

OR2x2_ASAP7_75t_L g5442 ( 
.A(n_5435),
.B(n_5425),
.Y(n_5442)
);

NAND2xp5_ASAP7_75t_L g5443 ( 
.A(n_5434),
.B(n_5426),
.Y(n_5443)
);

OR2x6_ASAP7_75t_L g5444 ( 
.A(n_5438),
.B(n_2222),
.Y(n_5444)
);

OR2x6_ASAP7_75t_L g5445 ( 
.A(n_5440),
.B(n_2222),
.Y(n_5445)
);

AOI221xp5_ASAP7_75t_L g5446 ( 
.A1(n_5443),
.A2(n_5436),
.B1(n_5439),
.B2(n_5437),
.C(n_5441),
.Y(n_5446)
);

AOI211xp5_ASAP7_75t_L g5447 ( 
.A1(n_5446),
.A2(n_5442),
.B(n_5445),
.C(n_5444),
.Y(n_5447)
);


endmodule