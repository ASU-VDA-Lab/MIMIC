module fake_jpeg_30481_n_213 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_213);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_30),
.B(n_48),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_34),
.Y(n_88)
);

CKINVDCx10_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_48),
.B1(n_50),
.B2(n_28),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_39),
.B(n_23),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_3),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_25),
.B1(n_12),
.B2(n_15),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_54),
.A2(n_68),
.B1(n_33),
.B2(n_43),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_63),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_29),
.B1(n_47),
.B2(n_46),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_27),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_25),
.B1(n_15),
.B2(n_12),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_79),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_34),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_16),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_55),
.B(n_73),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_70),
.B1(n_44),
.B2(n_33),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_116),
.B1(n_88),
.B2(n_6),
.Y(n_139)
);

OR2x4_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_23),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_109),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_112),
.B1(n_76),
.B2(n_77),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_83),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_3),
.B(n_4),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_26),
.C(n_5),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_80),
.C(n_78),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_60),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_88),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_56),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_131),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_85),
.B1(n_53),
.B2(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_139),
.B1(n_96),
.B2(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_125),
.Y(n_144)
);

OAI22x1_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_116),
.B1(n_111),
.B2(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_66),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_66),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_56),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_82),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_71),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_99),
.B(n_101),
.C(n_92),
.D(n_114),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_90),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_121),
.B1(n_137),
.B2(n_91),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_116),
.B(n_102),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_150),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_129),
.B(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_154),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

CKINVDCx10_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_125),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_117),
.B1(n_139),
.B2(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_162),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_117),
.B1(n_122),
.B2(n_136),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_126),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_118),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_124),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_153),
.B1(n_154),
.B2(n_143),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_145),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_176),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_149),
.B1(n_155),
.B2(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_181),
.B1(n_163),
.B2(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_177),
.Y(n_185)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_144),
.A3(n_156),
.B1(n_162),
.B2(n_160),
.C1(n_145),
.C2(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_179),
.Y(n_191)
);

OA21x2_ASAP7_75t_SL g179 ( 
.A1(n_159),
.A2(n_156),
.B(n_144),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_142),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_170),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_184),
.A2(n_187),
.B1(n_182),
.B2(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_190),
.B1(n_174),
.B2(n_189),
.Y(n_192)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_90),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_170),
.B1(n_165),
.B2(n_137),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_193),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_180),
.B1(n_182),
.B2(n_172),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_178),
.B1(n_173),
.B2(n_133),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_135),
.B(n_115),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_189),
.C(n_188),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_186),
.C(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_200),
.B(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_193),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_207),
.A2(n_208),
.B(n_187),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_199),
.B(n_197),
.C(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_209),
.B(n_97),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_210),
.B(n_95),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_98),
.Y(n_213)
);


endmodule