module fake_netlist_5_467_n_1121 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1121);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1121;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_1032;
wire n_929;
wire n_981;
wire n_941;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_1104;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1096;
wire n_976;
wire n_1095;
wire n_234;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_1114;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_1069;
wire n_236;
wire n_969;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_1091;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_857;
wire n_832;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_77),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_136),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_26),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_98),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_32),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_146),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_78),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_41),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_68),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_95),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_115),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_66),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_71),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_90),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_117),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_85),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_63),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_47),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_96),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_70),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_30),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_49),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_23),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_7),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_24),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_190),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_112),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_130),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_202),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_169),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_100),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_109),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_23),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_194),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_37),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_179),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_32),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_133),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_129),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_38),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_82),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_196),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_120),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_12),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_176),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_43),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_186),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_147),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_50),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_175),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_87),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_43),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_49),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_220),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_222),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_204),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_205),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_215),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_205),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_208),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_223),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_218),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_221),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_226),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_228),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_227),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_233),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_269),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_242),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_272),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_207),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_230),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_258),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_207),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_212),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_213),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_245),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_257),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_217),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_214),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_203),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_225),
.B(n_224),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_203),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_287),
.B(n_206),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_285),
.A2(n_253),
.B1(n_270),
.B2(n_214),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

AND2x4_ASAP7_75t_SL g336 ( 
.A(n_324),
.B(n_304),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_276),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_229),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_296),
.B(n_234),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_206),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_209),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_292),
.A2(n_297),
.B(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_280),
.B(n_256),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_279),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_209),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_238),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_275),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_281),
.B(n_210),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_299),
.A2(n_270),
.B1(n_253),
.B2(n_255),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_314),
.A2(n_240),
.B1(n_241),
.B2(n_236),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_303),
.A2(n_248),
.B1(n_243),
.B2(n_211),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_283),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_283),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_326),
.Y(n_363)
);

BUFx12f_ASAP7_75t_L g364 ( 
.A(n_284),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

AOI22x1_ASAP7_75t_SL g366 ( 
.A1(n_307),
.A2(n_210),
.B1(n_266),
.B2(n_211),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_216),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g373 ( 
.A(n_321),
.B(n_260),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_280),
.B(n_216),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_252),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_252),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

AND2x2_ASAP7_75t_SL g379 ( 
.A(n_325),
.B(n_264),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_314),
.A2(n_254),
.B1(n_266),
.B2(n_263),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_286),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_301),
.B(n_254),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_379),
.B(n_302),
.Y(n_385)
);

BUFx6f_ASAP7_75t_SL g386 ( 
.A(n_379),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_315),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_380),
.A2(n_291),
.B1(n_318),
.B2(n_311),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

CKINVDCx8_ASAP7_75t_R g394 ( 
.A(n_330),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_364),
.B(n_312),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_333),
.A2(n_310),
.B1(n_380),
.B2(n_355),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_383),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_336),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_333),
.A2(n_355),
.B1(n_359),
.B2(n_330),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_341),
.B(n_271),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

BUFx6f_ASAP7_75t_SL g407 ( 
.A(n_339),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_334),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

BUFx6f_ASAP7_75t_SL g414 ( 
.A(n_339),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_341),
.B(n_237),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_347),
.B(n_280),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_288),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_365),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_341),
.B(n_239),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_SL g425 ( 
.A(n_347),
.B(n_262),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_288),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_365),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_334),
.B(n_354),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_336),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_356),
.Y(n_434)
);

INVx8_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

BUFx6f_ASAP7_75t_SL g436 ( 
.A(n_339),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_361),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

CKINVDCx8_ASAP7_75t_R g443 ( 
.A(n_353),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_375),
.B(n_288),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_361),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_373),
.B(n_246),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_337),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_340),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_359),
.A2(n_294),
.B1(n_277),
.B2(n_278),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_337),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_336),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_337),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_332),
.A2(n_316),
.B1(n_311),
.B2(n_303),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_363),
.A2(n_278),
.B1(n_294),
.B2(n_277),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_362),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_362),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_327),
.A2(n_316),
.B(n_293),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_373),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_373),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_409),
.B(n_327),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_393),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_331),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_397),
.Y(n_467)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_372),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_416),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_387),
.B(n_389),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_331),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_387),
.B(n_339),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_400),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_342),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_426),
.B(n_363),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_389),
.B(n_342),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_425),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

NOR3xp33_ASAP7_75t_L g483 ( 
.A(n_396),
.B(n_360),
.C(n_372),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_403),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_389),
.B(n_410),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_432),
.Y(n_486)
);

BUFx5_ASAP7_75t_L g487 ( 
.A(n_447),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_410),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_425),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_401),
.A2(n_352),
.B1(n_329),
.B2(n_350),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_443),
.B(n_364),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_435),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_376),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_389),
.B(n_343),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_444),
.B(n_343),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_446),
.B(n_352),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_385),
.B(n_376),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_385),
.B(n_360),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_401),
.B(n_352),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_418),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_352),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_392),
.B(n_377),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_415),
.B(n_377),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_443),
.B(n_354),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_405),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_415),
.B(n_262),
.Y(n_510)
);

INVx8_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_424),
.B(n_366),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_408),
.B(n_350),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_411),
.B(n_335),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_424),
.B(n_366),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_458),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_398),
.B(n_317),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_421),
.B(n_335),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_422),
.B(n_335),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_406),
.B(n_368),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_430),
.B(n_263),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_431),
.B(n_437),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_458),
.B(n_346),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_449),
.B(n_306),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_386),
.A2(n_249),
.B1(n_250),
.B2(n_247),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_458),
.B(n_346),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_399),
.B(n_251),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_406),
.B(n_346),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_406),
.B(n_368),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_448),
.B(n_368),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_452),
.B(n_317),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_451),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_349),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_478),
.B(n_394),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_471),
.B(n_448),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_519),
.B(n_394),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

AO22x2_ASAP7_75t_L g544 ( 
.A1(n_483),
.A2(n_386),
.B1(n_395),
.B2(n_450),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

AO22x2_ASAP7_75t_L g546 ( 
.A1(n_495),
.A2(n_386),
.B1(n_455),
.B2(n_432),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_481),
.A2(n_308),
.B1(n_309),
.B2(n_306),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_489),
.A2(n_309),
.B1(n_308),
.B2(n_2),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_462),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_475),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_477),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_R g553 ( 
.A(n_491),
.B(n_435),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_465),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_479),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_472),
.B(n_476),
.Y(n_556)
);

AO22x2_ASAP7_75t_L g557 ( 
.A1(n_501),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_485),
.B(n_453),
.Y(n_558)
);

AO22x2_ASAP7_75t_L g559 ( 
.A1(n_517),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_435),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_L g562 ( 
.A(n_507),
.B(n_456),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_493),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_486),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_494),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_469),
.B(n_289),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_497),
.B(n_418),
.Y(n_567)
);

OR2x6_ASAP7_75t_SL g568 ( 
.A(n_513),
.B(n_289),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_506),
.A2(n_407),
.B1(n_436),
.B2(n_414),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_509),
.Y(n_570)
);

AND3x1_ASAP7_75t_L g571 ( 
.A(n_532),
.B(n_295),
.C(n_293),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_518),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_529),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_508),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_498),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_529),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_515),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_500),
.A2(n_407),
.B1(n_436),
.B2(n_414),
.Y(n_579)
);

AO22x2_ASAP7_75t_L g580 ( 
.A1(n_517),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_515),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_468),
.B(n_418),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

OAI221xp5_ASAP7_75t_L g585 ( 
.A1(n_512),
.A2(n_295),
.B1(n_298),
.B2(n_300),
.C(n_381),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_516),
.B(n_414),
.Y(n_586)
);

OAI221xp5_ASAP7_75t_L g587 ( 
.A1(n_510),
.A2(n_298),
.B1(n_300),
.B2(n_381),
.C(n_384),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_486),
.Y(n_588)
);

OAI221xp5_ASAP7_75t_L g589 ( 
.A1(n_510),
.A2(n_384),
.B1(n_381),
.B2(n_457),
.C(n_441),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_492),
.B(n_384),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_459),
.A2(n_436),
.B1(n_434),
.B2(n_441),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_529),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_511),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_471),
.B(n_419),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_492),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_460),
.A2(n_445),
.B1(n_440),
.B2(n_329),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_526),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_520),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_523),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_470),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_523),
.Y(n_601)
);

AO22x2_ASAP7_75t_L g602 ( 
.A1(n_470),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_602)
);

OAI21xp33_ASAP7_75t_L g603 ( 
.A1(n_527),
.A2(n_445),
.B(n_371),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_466),
.A2(n_329),
.B1(n_442),
.B2(n_429),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_511),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_534),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_534),
.Y(n_607)
);

CKINVDCx10_ASAP7_75t_R g608 ( 
.A(n_564),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_567),
.A2(n_471),
.B(n_474),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_556),
.A2(n_471),
.B(n_474),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_558),
.A2(n_496),
.B(n_480),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_542),
.B(n_575),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_575),
.B(n_530),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_558),
.A2(n_464),
.B(n_499),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_561),
.Y(n_615)
);

AO22x1_ASAP7_75t_L g616 ( 
.A1(n_540),
.A2(n_473),
.B1(n_484),
.B2(n_482),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_560),
.B(n_505),
.Y(n_617)
);

OAI21xp33_ASAP7_75t_L g618 ( 
.A1(n_597),
.A2(n_490),
.B(n_502),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_557),
.A2(n_482),
.B1(n_484),
.B2(n_473),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_604),
.A2(n_464),
.B(n_499),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_543),
.Y(n_621)
);

AO21x1_ASAP7_75t_L g622 ( 
.A1(n_591),
.A2(n_502),
.B(n_514),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_557),
.A2(n_488),
.B1(n_464),
.B2(n_531),
.Y(n_623)
);

AOI21xp33_ASAP7_75t_L g624 ( 
.A1(n_586),
.A2(n_524),
.B(n_522),
.Y(n_624)
);

OA21x2_ASAP7_75t_L g625 ( 
.A1(n_596),
.A2(n_528),
.B(n_533),
.Y(n_625)
);

BUFx2_ASAP7_75t_SL g626 ( 
.A(n_605),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_566),
.B(n_538),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_545),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_547),
.B(n_538),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_551),
.B(n_552),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_590),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_562),
.B(n_504),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_555),
.B(n_487),
.Y(n_633)
);

A2O1A1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_574),
.A2(n_592),
.B(n_577),
.C(n_565),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_544),
.A2(n_505),
.B1(n_511),
.B2(n_487),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g636 ( 
.A1(n_594),
.A2(n_539),
.B(n_504),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_563),
.A2(n_511),
.B(n_536),
.C(n_525),
.Y(n_637)
);

AOI21x1_ASAP7_75t_L g638 ( 
.A1(n_562),
.A2(n_583),
.B(n_535),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_541),
.A2(n_535),
.B(n_525),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_568),
.B(n_505),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_571),
.A2(n_505),
.B1(n_504),
.B2(n_536),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_576),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_588),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_570),
.B(n_487),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_593),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_596),
.A2(n_503),
.B(n_603),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_581),
.Y(n_647)
);

O2A1O1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_585),
.A2(n_349),
.B(n_362),
.C(n_371),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_595),
.B(n_374),
.C(n_349),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_572),
.B(n_487),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_573),
.B(n_487),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_571),
.A2(n_503),
.B1(n_329),
.B2(n_433),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_548),
.B(n_582),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_548),
.B(n_329),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_584),
.Y(n_656)
);

O2A1O1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_587),
.A2(n_371),
.B(n_374),
.C(n_370),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_544),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_598),
.Y(n_659)
);

BUFx4f_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

AOI21x1_ASAP7_75t_L g661 ( 
.A1(n_601),
.A2(n_351),
.B(n_369),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_600),
.A2(n_503),
.B1(n_442),
.B2(n_433),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_603),
.A2(n_503),
.B(n_427),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_606),
.A2(n_607),
.B(n_351),
.Y(n_664)
);

AOI21xp33_ASAP7_75t_L g665 ( 
.A1(n_600),
.A2(n_13),
.B(n_14),
.Y(n_665)
);

AOI221x1_ASAP7_75t_L g666 ( 
.A1(n_602),
.A2(n_419),
.B1(n_442),
.B2(n_433),
.C(n_429),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_579),
.B(n_419),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_647),
.Y(n_668)
);

NAND2x1_ASAP7_75t_L g669 ( 
.A(n_656),
.B(n_591),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_654),
.B(n_569),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_613),
.A2(n_546),
.B1(n_602),
.B2(n_549),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_579),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_612),
.A2(n_546),
.B1(n_549),
.B2(n_554),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_SL g674 ( 
.A1(n_658),
.A2(n_569),
.B1(n_554),
.B2(n_550),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_664),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_643),
.B(n_589),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_628),
.B(n_553),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_655),
.B(n_550),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_608),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_615),
.B(n_559),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_642),
.B(n_559),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_611),
.A2(n_351),
.B(n_369),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_619),
.B(n_487),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_636),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_659),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_631),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_627),
.B(n_487),
.Y(n_687)
);

AND3x1_ASAP7_75t_SL g688 ( 
.A(n_621),
.B(n_580),
.C(n_13),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_653),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_638),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_661),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_618),
.A2(n_580),
.B1(n_374),
.B2(n_370),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_631),
.B(n_419),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_645),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_619),
.A2(n_374),
.B1(n_369),
.B2(n_370),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_631),
.B(n_427),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_624),
.A2(n_610),
.B(n_634),
.C(n_637),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_625),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_630),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_629),
.B(n_442),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_646),
.A2(n_429),
.B(n_427),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_625),
.Y(n_702)
);

AOI211xp5_ASAP7_75t_L g703 ( 
.A1(n_665),
.A2(n_623),
.B(n_622),
.C(n_624),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_617),
.B(n_427),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_614),
.A2(n_433),
.B(n_429),
.C(n_368),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_616),
.B(n_14),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_650),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_SL g708 ( 
.A1(n_662),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_SL g709 ( 
.A1(n_640),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_660),
.Y(n_710)
);

BUFx8_ASAP7_75t_SL g711 ( 
.A(n_645),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_650),
.Y(n_712)
);

CKINVDCx8_ASAP7_75t_R g713 ( 
.A(n_645),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_632),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_667),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_660),
.B(n_18),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_633),
.B(n_19),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_656),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_667),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_644),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_635),
.B(n_368),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_665),
.B(n_368),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_651),
.B(n_19),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_623),
.B(n_54),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_632),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_648),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_652),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_649),
.B(n_641),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_641),
.B(n_20),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_715),
.B(n_719),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_697),
.A2(n_620),
.B(n_609),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_SL g732 ( 
.A(n_679),
.B(n_626),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_698),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_708),
.A2(n_662),
.B1(n_652),
.B2(n_666),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_694),
.B(n_639),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_685),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_670),
.B(n_699),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_686),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_694),
.Y(n_739)
);

BUFx12f_ASAP7_75t_L g740 ( 
.A(n_679),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_715),
.B(n_663),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_671),
.B(n_20),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_699),
.B(n_21),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_707),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_694),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_672),
.B(n_55),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_685),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_713),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_698),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_677),
.B(n_21),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_673),
.B(n_22),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_716),
.A2(n_657),
.B(n_24),
.C(n_25),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_689),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_705),
.A2(n_712),
.B(n_707),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_714),
.B(n_22),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_668),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_670),
.B(n_26),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_702),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_672),
.B(n_56),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_713),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_729),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_702),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_689),
.B(n_27),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_720),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_712),
.A2(n_58),
.B(n_57),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_715),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_674),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_720),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_729),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_715),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_683),
.A2(n_60),
.B(n_59),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_683),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_675),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_674),
.B(n_35),
.C(n_36),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_719),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_724),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_678),
.B(n_38),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_669),
.A2(n_138),
.B(n_200),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_703),
.A2(n_39),
.B(n_40),
.C(n_42),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_675),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_714),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_719),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_719),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_725),
.B(n_39),
.Y(n_785)
);

OAI221xp5_ASAP7_75t_L g786 ( 
.A1(n_709),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.C(n_45),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_725),
.B(n_44),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_672),
.B(n_61),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_669),
.A2(n_201),
.B(n_140),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_719),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_672),
.A2(n_710),
.B1(n_676),
.B2(n_728),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_693),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_680),
.Y(n_793)
);

AND2x6_ASAP7_75t_L g794 ( 
.A(n_724),
.B(n_62),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_703),
.B(n_45),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_718),
.Y(n_796)
);

BUFx4f_ASAP7_75t_SL g797 ( 
.A(n_680),
.Y(n_797)
);

CKINVDCx14_ASAP7_75t_R g798 ( 
.A(n_678),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_690),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_780),
.A2(n_709),
.B(n_727),
.C(n_728),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_744),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_780),
.A2(n_727),
.B(n_706),
.C(n_692),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_778),
.B(n_681),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_795),
.A2(n_723),
.B(n_717),
.C(n_726),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_737),
.B(n_681),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_744),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_795),
.A2(n_726),
.B(n_721),
.C(n_704),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_SL g808 ( 
.A1(n_786),
.A2(n_767),
.B1(n_777),
.B2(n_748),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_798),
.B(n_722),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_782),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_793),
.B(n_722),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_767),
.A2(n_718),
.B1(n_692),
.B2(n_687),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_784),
.B(n_721),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_782),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_740),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_791),
.B(n_743),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_796),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_736),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_734),
.A2(n_688),
.B(n_700),
.C(n_701),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_764),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_777),
.A2(n_696),
.B1(n_695),
.B2(n_690),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_775),
.A2(n_701),
.B(n_690),
.C(n_682),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_784),
.B(n_684),
.Y(n_823)
);

AOI221x1_ASAP7_75t_L g824 ( 
.A1(n_775),
.A2(n_684),
.B1(n_682),
.B2(n_691),
.C(n_50),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_742),
.B(n_695),
.Y(n_825)
);

O2A1O1Ixp5_ASAP7_75t_L g826 ( 
.A1(n_772),
.A2(n_684),
.B(n_691),
.C(n_48),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_750),
.B(n_64),
.Y(n_827)
);

O2A1O1Ixp5_ASAP7_75t_L g828 ( 
.A1(n_731),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_764),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_798),
.B(n_773),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_757),
.B(n_46),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_754),
.A2(n_143),
.B(n_198),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_748),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_761),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_792),
.B(n_51),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_773),
.A2(n_144),
.B(n_65),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_SL g838 ( 
.A(n_769),
.B(n_67),
.Y(n_838)
);

NOR2x1_ASAP7_75t_SL g839 ( 
.A(n_741),
.B(n_69),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_783),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_SL g841 ( 
.A1(n_752),
.A2(n_52),
.B(n_72),
.C(n_73),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_74),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_755),
.B(n_785),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_747),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_770),
.A2(n_75),
.B(n_76),
.C(n_79),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_787),
.B(n_751),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_797),
.B(n_80),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_768),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_768),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_756),
.B(n_81),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_788),
.B(n_83),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_749),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_SL g853 ( 
.A1(n_760),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_745),
.B(n_89),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_738),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_797),
.Y(n_856)
);

AOI211xp5_ASAP7_75t_L g857 ( 
.A1(n_770),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_753),
.B(n_94),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_749),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_733),
.B(n_97),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_788),
.B(n_99),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_760),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_783),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_788),
.B(n_101),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_732),
.Y(n_865)
);

O2A1O1Ixp5_ASAP7_75t_L g866 ( 
.A1(n_779),
.A2(n_102),
.B(n_103),
.C(n_104),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_739),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_855),
.B(n_769),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_808),
.A2(n_794),
.B1(n_759),
.B2(n_746),
.Y(n_869)
);

OAI21xp33_ASAP7_75t_L g870 ( 
.A1(n_835),
.A2(n_771),
.B(n_763),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_800),
.A2(n_746),
.B1(n_759),
.B2(n_730),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_816),
.A2(n_794),
.B1(n_765),
.B2(n_735),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_846),
.A2(n_794),
.B1(n_735),
.B2(n_789),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_830),
.B(n_790),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_840),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_SL g876 ( 
.A1(n_815),
.A2(n_794),
.B1(n_790),
.B2(n_766),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_843),
.A2(n_794),
.B1(n_741),
.B2(n_740),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_853),
.A2(n_741),
.B1(n_730),
.B2(n_776),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_801),
.Y(n_879)
);

OAI222xp33_ASAP7_75t_L g880 ( 
.A1(n_807),
.A2(n_730),
.B1(n_776),
.B2(n_766),
.C1(n_799),
.C2(n_774),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_809),
.A2(n_783),
.B1(n_799),
.B2(n_762),
.Y(n_881)
);

OAI21xp33_ASAP7_75t_L g882 ( 
.A1(n_835),
.A2(n_800),
.B(n_857),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_830),
.B(n_733),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_865),
.A2(n_781),
.B1(n_762),
.B2(n_758),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_827),
.A2(n_758),
.B1(n_106),
.B2(n_107),
.Y(n_885)
);

BUFx4f_ASAP7_75t_L g886 ( 
.A(n_840),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_815),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_806),
.Y(n_888)
);

OAI21xp33_ASAP7_75t_L g889 ( 
.A1(n_838),
.A2(n_105),
.B(n_108),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_818),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_825),
.A2(n_831),
.B1(n_803),
.B2(n_812),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_850),
.B(n_110),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_834),
.B(n_111),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_840),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_821),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_810),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_802),
.A2(n_862),
.B1(n_856),
.B2(n_847),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_837),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_804),
.B(n_122),
.C(n_123),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_867),
.Y(n_900)
);

BUFx8_ASAP7_75t_L g901 ( 
.A(n_851),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_SL g902 ( 
.A1(n_839),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_814),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_802),
.A2(n_127),
.B1(n_131),
.B2(n_134),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_836),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_847),
.A2(n_141),
.B1(n_142),
.B2(n_145),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_867),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_810),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_861),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_SL g910 ( 
.A1(n_864),
.A2(n_832),
.B1(n_824),
.B2(n_813),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_820),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_817),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_813),
.A2(n_805),
.B1(n_811),
.B2(n_860),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_822),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_813),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_882),
.A2(n_828),
.B(n_845),
.C(n_841),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_890),
.B(n_823),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_883),
.B(n_811),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_912),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_869),
.A2(n_842),
.B1(n_854),
.B2(n_860),
.Y(n_920)
);

NAND2x1_ASAP7_75t_L g921 ( 
.A(n_879),
.B(n_820),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_889),
.A2(n_841),
.B(n_822),
.C(n_826),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_911),
.B(n_896),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_888),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_874),
.B(n_863),
.Y(n_925)
);

NOR2x1_ASAP7_75t_R g926 ( 
.A(n_887),
.B(n_858),
.Y(n_926)
);

AOI211xp5_ASAP7_75t_L g927 ( 
.A1(n_914),
.A2(n_897),
.B(n_904),
.C(n_870),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_903),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_908),
.B(n_823),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_907),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_913),
.B(n_859),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_871),
.B(n_823),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_895),
.A2(n_819),
.B1(n_844),
.B2(n_833),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_899),
.A2(n_866),
.B(n_819),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_913),
.B(n_900),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_875),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_877),
.B(n_891),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_895),
.A2(n_849),
.B1(n_848),
.B2(n_840),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_884),
.Y(n_939)
);

AOI221xp5_ASAP7_75t_L g940 ( 
.A1(n_891),
.A2(n_829),
.B1(n_820),
.B2(n_852),
.C(n_859),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_875),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_894),
.B(n_875),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_877),
.B(n_852),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_892),
.B(n_829),
.Y(n_944)
);

OA21x2_ASAP7_75t_L g945 ( 
.A1(n_880),
.A2(n_829),
.B(n_159),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_868),
.B(n_158),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_924),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_926),
.B(n_901),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_917),
.B(n_876),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_924),
.B(n_881),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_942),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_939),
.B(n_875),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_919),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_921),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_917),
.B(n_918),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_928),
.Y(n_956)
);

NOR2x1_ASAP7_75t_SL g957 ( 
.A(n_932),
.B(n_894),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_917),
.B(n_910),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_918),
.B(n_873),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_937),
.A2(n_934),
.B1(n_932),
.B2(n_872),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_923),
.B(n_929),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_921),
.Y(n_962)
);

BUFx4f_ASAP7_75t_L g963 ( 
.A(n_945),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_923),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_939),
.B(n_873),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_935),
.B(n_872),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_937),
.A2(n_898),
.B1(n_909),
.B2(n_905),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_923),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_947),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_963),
.A2(n_927),
.B(n_916),
.C(n_922),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_963),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_963),
.A2(n_933),
.B(n_932),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_963),
.A2(n_935),
.B(n_898),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_947),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_953),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_953),
.B(n_925),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_960),
.B(n_930),
.Y(n_977)
);

INVx4_ASAP7_75t_SL g978 ( 
.A(n_951),
.Y(n_978)
);

OA21x2_ASAP7_75t_L g979 ( 
.A1(n_954),
.A2(n_940),
.B(n_936),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_964),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_956),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_951),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_966),
.B(n_925),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_948),
.B(n_930),
.Y(n_984)
);

OA21x2_ASAP7_75t_L g985 ( 
.A1(n_954),
.A2(n_936),
.B(n_943),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_971),
.B(n_962),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_978),
.B(n_957),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_975),
.B(n_966),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_981),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_970),
.B(n_959),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_971),
.B(n_961),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_985),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_978),
.B(n_957),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_971),
.B(n_961),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_978),
.B(n_954),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_983),
.B(n_959),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_976),
.B(n_959),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_989),
.Y(n_998)
);

NOR3xp33_ASAP7_75t_L g999 ( 
.A(n_990),
.B(n_977),
.C(n_973),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_987),
.B(n_993),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_993),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_988),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_993),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_987),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_995),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_992),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_999),
.A2(n_972),
.B1(n_971),
.B2(n_967),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_999),
.A2(n_971),
.B1(n_965),
.B2(n_945),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_1000),
.B(n_991),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_1005),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_1005),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_1000),
.B(n_994),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_1007),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_1010),
.B(n_1002),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1011),
.B(n_1001),
.Y(n_1015)
);

AOI22x1_ASAP7_75t_L g1016 ( 
.A1(n_1009),
.A2(n_1001),
.B1(n_1004),
.B2(n_1012),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_1008),
.B(n_996),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1008),
.Y(n_1018)
);

AO22x1_ASAP7_75t_L g1019 ( 
.A1(n_1007),
.A2(n_1003),
.B1(n_1005),
.B2(n_1004),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_1010),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1009),
.B(n_1003),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_1010),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1022),
.B(n_998),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1020),
.Y(n_1024)
);

BUFx8_ASAP7_75t_SL g1025 ( 
.A(n_1021),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1014),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1022),
.B(n_998),
.Y(n_1027)
);

AO22x1_ASAP7_75t_L g1028 ( 
.A1(n_1018),
.A2(n_1003),
.B1(n_995),
.B2(n_982),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1015),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_1013),
.B(n_984),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1030),
.B(n_1019),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1024),
.B(n_1017),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_1030),
.B(n_1025),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1023),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1027),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1028),
.B(n_997),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_1031),
.B(n_1016),
.C(n_1003),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1035),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_1033),
.A2(n_1032),
.B(n_1036),
.C(n_1034),
.Y(n_1040)
);

OAI211xp5_ASAP7_75t_L g1041 ( 
.A1(n_1032),
.A2(n_1003),
.B(n_986),
.C(n_1006),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_L g1042 ( 
.A(n_1037),
.B(n_1006),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1042),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1039),
.B(n_1003),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1040),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1038),
.B(n_982),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1041),
.B(n_978),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1038),
.B(n_995),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

NAND4xp25_ASAP7_75t_L g1050 ( 
.A(n_1046),
.B(n_946),
.C(n_893),
.D(n_902),
.Y(n_1050)
);

AOI211xp5_ASAP7_75t_SL g1051 ( 
.A1(n_1045),
.A2(n_1047),
.B(n_1043),
.C(n_1048),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_1044),
.B(n_906),
.C(n_965),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_1045),
.A2(n_992),
.B(n_905),
.C(n_909),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_R g1054 ( 
.A(n_1045),
.B(n_161),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_SL g1055 ( 
.A(n_1051),
.B(n_952),
.C(n_950),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_1053),
.A2(n_1049),
.B(n_1052),
.C(n_1050),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1054),
.B(n_980),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1052),
.B(n_978),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1049),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1051),
.B(n_915),
.C(n_979),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1051),
.B(n_980),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1049),
.B(n_980),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_L g1063 ( 
.A(n_1059),
.B(n_885),
.C(n_952),
.Y(n_1063)
);

CKINVDCx6p67_ASAP7_75t_R g1064 ( 
.A(n_1061),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_1060),
.A2(n_985),
.B1(n_979),
.B2(n_981),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1055),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1062),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_SL g1068 ( 
.A(n_1058),
.B(n_958),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_1056),
.B(n_985),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1057),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1064),
.B(n_985),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1068),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1069),
.Y(n_1073)
);

AOI31xp33_ASAP7_75t_L g1074 ( 
.A1(n_1066),
.A2(n_1067),
.A3(n_1070),
.B(n_1065),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_1063),
.B(n_979),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_L g1076 ( 
.A(n_1070),
.B(n_979),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1068),
.Y(n_1077)
);

AOI322xp5_ASAP7_75t_L g1078 ( 
.A1(n_1066),
.A2(n_915),
.A3(n_958),
.B1(n_920),
.B2(n_878),
.C1(n_949),
.C2(n_969),
.Y(n_1078)
);

NAND3xp33_ASAP7_75t_SL g1079 ( 
.A(n_1066),
.B(n_958),
.C(n_878),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1072),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1073),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1077),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1074),
.B(n_974),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1071),
.B(n_974),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1079),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_1076),
.Y(n_1086)
);

OA22x2_ASAP7_75t_L g1087 ( 
.A1(n_1075),
.A2(n_969),
.B1(n_974),
.B2(n_962),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1078),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1073),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1077),
.Y(n_1090)
);

BUFx8_ASAP7_75t_L g1091 ( 
.A(n_1077),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1073),
.Y(n_1092)
);

NAND4xp75_ASAP7_75t_L g1093 ( 
.A(n_1082),
.B(n_945),
.C(n_949),
.D(n_950),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_1091),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_1091),
.B(n_901),
.C(n_956),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_1086),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1083),
.B(n_964),
.Y(n_1097)
);

AOI221xp5_ASAP7_75t_L g1098 ( 
.A1(n_1090),
.A2(n_949),
.B1(n_968),
.B2(n_964),
.C(n_942),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_1080),
.Y(n_1099)
);

OAI32xp33_ASAP7_75t_L g1100 ( 
.A1(n_1081),
.A2(n_941),
.A3(n_968),
.B1(n_944),
.B2(n_955),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_1089),
.B(n_942),
.C(n_945),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_1094),
.B(n_1092),
.C(n_1085),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1099),
.A2(n_1088),
.B1(n_1087),
.B2(n_1084),
.Y(n_1103)
);

OAI211xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1096),
.A2(n_162),
.B(n_164),
.C(n_165),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1095),
.A2(n_941),
.B1(n_886),
.B2(n_932),
.Y(n_1105)
);

XNOR2xp5_ASAP7_75t_L g1106 ( 
.A(n_1097),
.B(n_166),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1100),
.A2(n_938),
.B(n_168),
.C(n_170),
.Y(n_1107)
);

AOI211xp5_ASAP7_75t_L g1108 ( 
.A1(n_1102),
.A2(n_1104),
.B(n_1106),
.C(n_1107),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1103),
.A2(n_1101),
.B1(n_1093),
.B2(n_1098),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_L g1110 ( 
.A(n_1105),
.B(n_167),
.C(n_171),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1110),
.A2(n_1109),
.B1(n_1108),
.B2(n_886),
.Y(n_1111)
);

XNOR2xp5_ASAP7_75t_L g1112 ( 
.A(n_1111),
.B(n_172),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1112),
.A2(n_955),
.B(n_943),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1112),
.A2(n_174),
.B(n_177),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_1114),
.B(n_1113),
.Y(n_1115)
);

FAx1_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_178),
.CI(n_181),
.CON(n_1116),
.SN(n_1116)
);

AOI21xp33_ASAP7_75t_L g1117 ( 
.A1(n_1114),
.A2(n_182),
.B(n_183),
.Y(n_1117)
);

AO21x2_ASAP7_75t_L g1118 ( 
.A1(n_1117),
.A2(n_185),
.B(n_187),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_1115),
.B(n_189),
.Y(n_1119)
);

OAI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1119),
.A2(n_1116),
.B1(n_931),
.B2(n_955),
.Y(n_1120)
);

AOI211xp5_ASAP7_75t_L g1121 ( 
.A1(n_1120),
.A2(n_1118),
.B(n_191),
.C(n_192),
.Y(n_1121)
);


endmodule