module fake_ariane_3164_n_1568 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1568);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1568;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_208;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_93),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_16),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_104),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_36),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_54),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_4),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_88),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_9),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_36),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_2),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_2),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_85),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_51),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_12),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_29),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_33),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_69),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_39),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_40),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_58),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_139),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_123),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_121),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_0),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_47),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_49),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_72),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_68),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_23),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_1),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_111),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_20),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_100),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_33),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_21),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_3),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_18),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_81),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_0),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_110),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_91),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_56),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_70),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_92),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_76),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_19),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_60),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_13),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_82),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_51),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_35),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_79),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_37),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_47),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_55),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_35),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_39),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_73),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_40),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_67),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_115),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_113),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_25),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_18),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_61),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_11),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_6),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_109),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_5),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_10),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_107),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_41),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_20),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_94),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_78),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_42),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_86),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_27),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_37),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_53),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_31),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_57),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_96),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_8),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_90),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_41),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_87),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_64),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_62),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_114),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_99),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_136),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_97),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_135),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_66),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_3),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_102),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_80),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_5),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_52),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_50),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_17),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_16),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_130),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_125),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_75),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_74),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_157),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_R g291 ( 
.A(n_147),
.B(n_160),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_152),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_152),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_152),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_172),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_176),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_194),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_152),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_152),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_183),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_244),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_202),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_183),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_243),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_202),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_167),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_186),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_202),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_202),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_262),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_156),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_275),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_163),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_199),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_202),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_149),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_186),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_169),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_171),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_239),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_239),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_239),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_173),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_285),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_166),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_199),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_285),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_266),
.B(n_6),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_174),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_159),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_159),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_175),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_272),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_185),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_242),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_155),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_242),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_181),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_177),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_187),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_177),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_195),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_190),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_190),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_242),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_273),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_220),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_273),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_196),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_204),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_292),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_291),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_295),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_293),
.Y(n_369)
);

CKINVDCx11_ASAP7_75t_R g370 ( 
.A(n_311),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_209),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_298),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_313),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_320),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_294),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_294),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_324),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_299),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_296),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_297),
.B(n_184),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_316),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_299),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_300),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_307),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_162),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_302),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_303),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_303),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_306),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_306),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_310),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_339),
.B(n_231),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_341),
.B(n_182),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_327),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_314),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_340),
.B(n_209),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_343),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_349),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_331),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_341),
.B(n_188),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_351),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

INVx6_ASAP7_75t_L g418 ( 
.A(n_297),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_192),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_338),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_360),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_317),
.B(n_219),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_362),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_301),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_344),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_348),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_329),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_356),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_357),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_408),
.B(n_359),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_418),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_364),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_371),
.B(n_304),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_365),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_290),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_373),
.B(n_333),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_346),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_366),
.B(n_201),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_393),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_337),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_414),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_342),
.Y(n_456)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_371),
.B(n_225),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_410),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_389),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_371),
.B(n_350),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_318),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_423),
.B(n_151),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_402),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_371),
.B(n_345),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_418),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_309),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_397),
.A2(n_250),
.B1(n_232),
.B2(n_238),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_363),
.B(n_321),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_363),
.A2(n_161),
.B1(n_280),
.B2(n_150),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_350),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_398),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_371),
.B(n_332),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_386),
.B(n_332),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_378),
.B(n_151),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_378),
.B(n_153),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_387),
.B(n_153),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_386),
.A2(n_245),
.B1(n_278),
.B2(n_254),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_387),
.A2(n_150),
.B1(n_148),
.B2(n_280),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_403),
.B(n_203),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_L g490 ( 
.A(n_403),
.B(n_212),
.Y(n_490)
);

CKINVDCx6p67_ASAP7_75t_R g491 ( 
.A(n_370),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_381),
.A2(n_412),
.B1(n_420),
.B2(n_398),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_413),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_415),
.B(n_154),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_415),
.B(n_334),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_374),
.B(n_148),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_412),
.B(n_352),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_367),
.B(n_154),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_368),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_420),
.A2(n_286),
.B1(n_246),
.B2(n_361),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_368),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_419),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_372),
.A2(n_228),
.B1(n_264),
.B2(n_253),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_334),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_382),
.B(n_161),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_L g510 ( 
.A1(n_376),
.A2(n_281),
.B1(n_284),
.B2(n_283),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_431),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_374),
.B(n_335),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_390),
.B(n_354),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_368),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_379),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_379),
.Y(n_517)
);

A2O1A1Ixp33_ASAP7_75t_L g518 ( 
.A1(n_390),
.A2(n_235),
.B(n_258),
.C(n_261),
.Y(n_518)
);

AO21x2_ASAP7_75t_L g519 ( 
.A1(n_392),
.A2(n_269),
.B(n_218),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_430),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_429),
.B(n_158),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_392),
.A2(n_361),
.B1(n_358),
.B2(n_355),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_395),
.B(n_234),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_395),
.B(n_335),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_401),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_401),
.B(n_355),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_379),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_404),
.B(n_336),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_380),
.B(n_385),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_432),
.B(n_282),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_404),
.B(n_358),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_416),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_416),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_417),
.B(n_427),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g535 ( 
.A1(n_417),
.A2(n_284),
.B1(n_206),
.B2(n_207),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_427),
.A2(n_211),
.B1(n_229),
.B2(n_241),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_368),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_383),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_383),
.B(n_158),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_368),
.B(n_208),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_383),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_368),
.B(n_212),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_391),
.B(n_221),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_391),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_391),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_396),
.B(n_164),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_399),
.B(n_273),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_396),
.B(n_336),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_405),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_405),
.B(n_277),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_405),
.B(n_164),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_394),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_409),
.B(n_165),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_409),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_409),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_422),
.B(n_234),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_370),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_422),
.B(n_165),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_422),
.B(n_217),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_426),
.A2(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_394),
.B(n_224),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_426),
.B(n_224),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_394),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_394),
.B(n_274),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_394),
.B(n_274),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_394),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_407),
.B(n_276),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_407),
.B(n_276),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_407),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_407),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_407),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_407),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_411),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_465),
.B(n_421),
.Y(n_575)
);

AO221x1_ASAP7_75t_L g576 ( 
.A1(n_510),
.A2(n_520),
.B1(n_488),
.B2(n_476),
.C(n_492),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_478),
.B(n_287),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_443),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_459),
.B(n_287),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_540),
.A2(n_249),
.B1(n_248),
.B2(n_252),
.Y(n_580)
);

A2O1A1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_469),
.A2(n_288),
.B(n_289),
.C(n_170),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_494),
.B(n_457),
.Y(n_582)
);

NOR3xp33_ASAP7_75t_L g583 ( 
.A(n_494),
.B(n_288),
.C(n_289),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_516),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_497),
.B(n_457),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_493),
.B(n_168),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_444),
.B(n_433),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_497),
.B(n_10),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_438),
.B(n_178),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_R g590 ( 
.A(n_458),
.B(n_557),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_540),
.B(n_212),
.Y(n_591)
);

NOR2xp67_ASAP7_75t_L g592 ( 
.A(n_444),
.B(n_440),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_517),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_455),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_438),
.B(n_179),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_443),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_517),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_480),
.B(n_180),
.Y(n_599)
);

O2A1O1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_452),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_527),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_527),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_490),
.A2(n_271),
.B1(n_268),
.B2(n_267),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_465),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_490),
.A2(n_265),
.B1(n_263),
.B2(n_260),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_480),
.B(n_189),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_480),
.B(n_191),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_511),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_438),
.B(n_193),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_499),
.A2(n_255),
.B(n_197),
.C(n_251),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_474),
.B(n_198),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_559),
.B(n_200),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_474),
.B(n_205),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_449),
.B(n_15),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_559),
.B(n_247),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_449),
.B(n_210),
.Y(n_617)
);

AND2x6_ASAP7_75t_SL g618 ( 
.A(n_496),
.B(n_17),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_532),
.A2(n_227),
.B1(n_240),
.B2(n_237),
.Y(n_619)
);

INVxp33_ASAP7_75t_L g620 ( 
.A(n_441),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_482),
.B(n_21),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_458),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_460),
.B(n_216),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_538),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_466),
.B(n_230),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_545),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_519),
.A2(n_252),
.B1(n_212),
.B2(n_215),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_556),
.B(n_214),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_473),
.B(n_236),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_545),
.Y(n_630)
);

BUFx8_ASAP7_75t_L g631 ( 
.A(n_473),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_483),
.B(n_22),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_523),
.B(n_215),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_486),
.B(n_22),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_489),
.B(n_233),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_555),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_547),
.B(n_446),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_434),
.B(n_213),
.C(n_24),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_489),
.B(n_23),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_447),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_496),
.A2(n_215),
.B1(n_212),
.B2(n_252),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_456),
.B(n_212),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_455),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_496),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_479),
.B(n_212),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_448),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_507),
.B(n_252),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_523),
.B(n_215),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_479),
.B(n_215),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_525),
.Y(n_651)
);

CKINVDCx14_ASAP7_75t_R g652 ( 
.A(n_441),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_L g653 ( 
.A(n_495),
.B(n_530),
.C(n_464),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_508),
.B(n_215),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_519),
.A2(n_215),
.B1(n_25),
.B2(n_26),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_500),
.B(n_24),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_523),
.B(n_215),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_574),
.B(n_26),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_491),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_513),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_513),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_467),
.B(n_28),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_535),
.B(n_28),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_463),
.B(n_30),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_461),
.B(n_31),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_463),
.B(n_34),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_513),
.Y(n_667)
);

NOR2x1p5_ASAP7_75t_L g668 ( 
.A(n_491),
.B(n_38),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_519),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_448),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_467),
.B(n_43),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_467),
.B(n_477),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_511),
.B(n_44),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_525),
.B(n_45),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_436),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_437),
.A2(n_485),
.B1(n_439),
.B2(n_442),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_450),
.B(n_46),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_524),
.B(n_48),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_471),
.A2(n_50),
.B1(n_52),
.B2(n_63),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_534),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_565),
.A2(n_83),
.B(n_89),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_524),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_513),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_528),
.B(n_143),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_528),
.B(n_98),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_475),
.B(n_142),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_484),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_453),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_533),
.B(n_106),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_470),
.B(n_108),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_526),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_574),
.B(n_116),
.Y(n_692)
);

O2A1O1Ixp5_ASAP7_75t_L g693 ( 
.A1(n_561),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_548),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_521),
.A2(n_553),
.B1(n_539),
.B2(n_551),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_453),
.Y(n_696)
);

XOR2xp5_ASAP7_75t_L g697 ( 
.A(n_509),
.B(n_120),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_515),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_548),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_546),
.A2(n_124),
.B1(n_133),
.B2(n_138),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_L g701 ( 
.A1(n_566),
.A2(n_569),
.B(n_568),
.C(n_481),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_454),
.B(n_472),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_557),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_548),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_454),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_462),
.B(n_506),
.Y(n_706)
);

INVx6_ASAP7_75t_L g707 ( 
.A(n_574),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_514),
.A2(n_531),
.B(n_512),
.C(n_506),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_481),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_502),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_505),
.B(n_512),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_505),
.B(n_563),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_558),
.A2(n_536),
.B1(n_550),
.B2(n_543),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_544),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_549),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_515),
.B(n_537),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_530),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_515),
.B(n_537),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_549),
.B(n_541),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_645),
.B(n_529),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_588),
.A2(n_663),
.B(n_615),
.C(n_662),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_708),
.A2(n_567),
.B(n_570),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_701),
.A2(n_567),
.B(n_573),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_585),
.B(n_498),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_661),
.B(n_667),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_615),
.B(n_503),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_672),
.A2(n_537),
.B(n_564),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_680),
.B(n_487),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_702),
.A2(n_572),
.B(n_564),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_605),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_585),
.B(n_664),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_584),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_582),
.B(n_717),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_592),
.B(n_498),
.Y(n_734)
);

AOI21x1_ASAP7_75t_L g735 ( 
.A1(n_633),
.A2(n_562),
.B(n_554),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_686),
.A2(n_571),
.B(n_572),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_588),
.A2(n_560),
.B1(n_564),
.B2(n_542),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_691),
.B(n_522),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_640),
.B(n_509),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_644),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_575),
.B(n_518),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_587),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_713),
.A2(n_435),
.B1(n_468),
.B2(n_504),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_594),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_623),
.B(n_468),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_707),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_596),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_597),
.A2(n_504),
.B1(n_552),
.B2(n_445),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_712),
.A2(n_445),
.B(n_501),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_631),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_716),
.A2(n_504),
.B(n_552),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_682),
.B(n_617),
.Y(n_752)
);

INVx3_ASAP7_75t_SL g753 ( 
.A(n_659),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_718),
.A2(n_504),
.B(n_552),
.Y(n_754)
);

AOI21x1_ASAP7_75t_L g755 ( 
.A1(n_633),
.A2(n_552),
.B(n_445),
.Y(n_755)
);

OAI21xp33_ASAP7_75t_L g756 ( 
.A1(n_621),
.A2(n_445),
.B(n_501),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_694),
.B(n_501),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_594),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_706),
.A2(n_501),
.B(n_711),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_660),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_631),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_621),
.A2(n_632),
.B(n_634),
.C(n_656),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_690),
.A2(n_576),
.B1(n_580),
.B2(n_634),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_699),
.B(n_704),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_687),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_577),
.B(n_579),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_711),
.A2(n_719),
.B(n_647),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_683),
.B(n_622),
.Y(n_768)
);

INVx11_ASAP7_75t_L g769 ( 
.A(n_622),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_707),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_644),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_632),
.A2(n_656),
.B(n_580),
.C(n_690),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_641),
.A2(n_696),
.B(n_647),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_641),
.A2(n_688),
.B(n_670),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_638),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_653),
.A2(n_583),
.B1(n_636),
.B2(n_610),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_684),
.A2(n_685),
.B(n_710),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_676),
.B(n_613),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_616),
.B(n_599),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_673),
.A2(n_655),
.B(n_695),
.C(n_586),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_673),
.B(n_581),
.C(n_655),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_705),
.A2(n_709),
.B(n_646),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_607),
.B(n_608),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_651),
.B(n_678),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_714),
.B(n_715),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_650),
.A2(n_654),
.B(n_705),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_689),
.A2(n_715),
.B(n_714),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_660),
.Y(n_788)
);

AND2x6_ASAP7_75t_L g789 ( 
.A(n_642),
.B(n_609),
.Y(n_789)
);

AOI21x1_ASAP7_75t_L g790 ( 
.A1(n_649),
.A2(n_657),
.B(n_591),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_671),
.A2(n_665),
.B(n_643),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_677),
.A2(n_674),
.B(n_601),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_593),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_598),
.A2(n_630),
.B(n_637),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_598),
.A2(n_630),
.B(n_624),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_628),
.B(n_589),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_601),
.A2(n_626),
.B(n_637),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_595),
.B(n_604),
.Y(n_798)
);

AOI22x1_ASAP7_75t_L g799 ( 
.A1(n_681),
.A2(n_624),
.B1(n_604),
.B2(n_626),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_658),
.B(n_603),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_669),
.A2(n_600),
.B(n_666),
.C(n_679),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_602),
.A2(n_635),
.B(n_698),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_590),
.B(n_594),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_606),
.A2(n_614),
.B1(n_612),
.B2(n_625),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_602),
.B(n_635),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_594),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_611),
.A2(n_693),
.B(n_627),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_648),
.A2(n_629),
.B(n_627),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_692),
.B(n_639),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_619),
.A2(n_675),
.B(n_700),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_692),
.A2(n_703),
.B(n_697),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_692),
.A2(n_620),
.B(n_618),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_652),
.A2(n_672),
.B(n_702),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_668),
.B(n_494),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_605),
.B(n_400),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_615),
.A2(n_588),
.B(n_585),
.C(n_664),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_605),
.Y(n_817)
);

AO22x1_ASAP7_75t_L g818 ( 
.A1(n_631),
.A2(n_432),
.B1(n_430),
.B2(n_298),
.Y(n_818)
);

OR2x4_ASAP7_75t_L g819 ( 
.A(n_588),
.B(n_530),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_578),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_585),
.B(n_295),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_L g822 ( 
.A(n_605),
.B(n_473),
.C(n_494),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_588),
.A2(n_663),
.B(n_615),
.C(n_494),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_615),
.B(n_478),
.Y(n_825)
);

INVx8_ASAP7_75t_L g826 ( 
.A(n_660),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_585),
.B(n_295),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_587),
.B(n_444),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_830)
);

CKINVDCx8_ASAP7_75t_R g831 ( 
.A(n_659),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_615),
.B(n_478),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_645),
.B(n_494),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_605),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_835)
);

CKINVDCx10_ASAP7_75t_R g836 ( 
.A(n_659),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_578),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_615),
.B(n_478),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_588),
.A2(n_663),
.B(n_615),
.C(n_494),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_585),
.B(n_295),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_585),
.B(n_410),
.C(n_408),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_645),
.B(n_494),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_645),
.B(n_494),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_713),
.A2(n_680),
.B1(n_596),
.B2(n_597),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_578),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_615),
.B(n_478),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_631),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_605),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_615),
.A2(n_588),
.B(n_585),
.C(n_664),
.Y(n_854)
);

NAND2x2_ASAP7_75t_L g855 ( 
.A(n_668),
.B(n_494),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_615),
.B(n_478),
.Y(n_857)
);

NAND2x1p5_ASAP7_75t_L g858 ( 
.A(n_645),
.B(n_661),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_708),
.A2(n_701),
.B(n_712),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_578),
.Y(n_860)
);

OAI21xp33_ASAP7_75t_L g861 ( 
.A1(n_588),
.A2(n_410),
.B(n_408),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_585),
.B(n_295),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_575),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_575),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_585),
.B(n_295),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_645),
.B(n_494),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_615),
.A2(n_588),
.B(n_585),
.C(n_664),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_585),
.A2(n_582),
.B1(n_588),
.B2(n_690),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_615),
.B(n_478),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_615),
.B(n_478),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_615),
.B(n_478),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_672),
.A2(n_702),
.B(n_716),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_731),
.B(n_848),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_816),
.B(n_854),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_826),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_825),
.A2(n_838),
.B(n_832),
.Y(n_878)
);

O2A1O1Ixp5_ASAP7_75t_L g879 ( 
.A1(n_762),
.A2(n_810),
.B(n_868),
.C(n_807),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_850),
.A2(n_871),
.B(n_857),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_724),
.B(n_778),
.Y(n_881)
);

BUFx2_ASAP7_75t_SL g882 ( 
.A(n_831),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_815),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_821),
.B(n_827),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_775),
.B(n_844),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_852),
.A2(n_863),
.B(n_856),
.Y(n_886)
);

INVx3_ASAP7_75t_SL g887 ( 
.A(n_753),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_822),
.B(n_843),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_864),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_872),
.B(n_873),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_787),
.A2(n_782),
.B(n_755),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_828),
.B(n_742),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_721),
.A2(n_823),
.B(n_841),
.C(n_772),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_869),
.B(n_766),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_782),
.A2(n_797),
.B(n_795),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_870),
.A2(n_874),
.B(n_829),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_870),
.A2(n_874),
.B(n_830),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_739),
.B(n_862),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_769),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_735),
.A2(n_835),
.B(n_824),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_SL g901 ( 
.A1(n_756),
.A2(n_801),
.B(n_763),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_765),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_839),
.A2(n_840),
.B(n_846),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_866),
.B(n_720),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_779),
.B(n_726),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_865),
.B(n_730),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_788),
.B(n_720),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_842),
.A2(n_781),
.B(n_767),
.Y(n_908)
);

AO21x2_ASAP7_75t_L g909 ( 
.A1(n_802),
.A2(n_808),
.B(n_723),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_744),
.B(n_758),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_826),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_861),
.A2(n_800),
.B1(n_733),
.B2(n_817),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_SL g913 ( 
.A(n_851),
.B(n_761),
.Y(n_913)
);

INVx5_ASAP7_75t_L g914 ( 
.A(n_826),
.Y(n_914)
);

AND2x2_ASAP7_75t_SL g915 ( 
.A(n_809),
.B(n_750),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_722),
.A2(n_727),
.B(n_729),
.Y(n_916)
);

AND2x6_ASAP7_75t_L g917 ( 
.A(n_744),
.B(n_758),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_773),
.A2(n_774),
.B(n_754),
.Y(n_918)
);

AOI21xp33_ASAP7_75t_L g919 ( 
.A1(n_783),
.A2(n_809),
.B(n_804),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_746),
.B(n_811),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_752),
.B(n_747),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_749),
.A2(n_751),
.B(n_759),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_734),
.B(n_819),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_820),
.B(n_837),
.Y(n_924)
);

BUFx4f_ASAP7_75t_L g925 ( 
.A(n_858),
.Y(n_925)
);

NAND3x1_ASAP7_75t_L g926 ( 
.A(n_811),
.B(n_812),
.C(n_741),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_776),
.A2(n_796),
.B(n_813),
.C(n_784),
.Y(n_927)
);

AOI21xp33_ASAP7_75t_L g928 ( 
.A1(n_737),
.A2(n_785),
.B(n_786),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_834),
.B(n_853),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_727),
.A2(n_794),
.B(n_729),
.Y(n_930)
);

OA22x2_ASAP7_75t_L g931 ( 
.A1(n_728),
.A2(n_814),
.B1(n_849),
.B2(n_860),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_818),
.B(n_812),
.Y(n_932)
);

NAND2x1_ASAP7_75t_SL g933 ( 
.A(n_740),
.B(n_771),
.Y(n_933)
);

INVxp33_ASAP7_75t_SL g934 ( 
.A(n_836),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_806),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_738),
.B(n_793),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_790),
.A2(n_748),
.B(n_805),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_725),
.B(n_858),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_L g939 ( 
.A(n_789),
.B(n_758),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_725),
.B(n_867),
.Y(n_940)
);

NAND2x1_ASAP7_75t_L g941 ( 
.A(n_806),
.B(n_744),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_743),
.A2(n_757),
.B(n_798),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_764),
.Y(n_943)
);

AOI21x1_ASAP7_75t_SL g944 ( 
.A1(n_819),
.A2(n_855),
.B(n_803),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_745),
.A2(n_740),
.B(n_771),
.Y(n_945)
);

OAI22x1_ASAP7_75t_L g946 ( 
.A1(n_833),
.A2(n_847),
.B1(n_845),
.B2(n_768),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_770),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_789),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_789),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_L g950 ( 
.A(n_789),
.B(n_762),
.C(n_816),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_736),
.A2(n_799),
.B(n_787),
.Y(n_951)
);

OA21x2_ASAP7_75t_L g952 ( 
.A1(n_736),
.A2(n_859),
.B(n_791),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_815),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_731),
.B(n_680),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_816),
.A2(n_868),
.B(n_854),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_732),
.Y(n_956)
);

NOR2x1_ASAP7_75t_L g957 ( 
.A(n_761),
.B(n_844),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_732),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_825),
.A2(n_838),
.B(n_832),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_777),
.A2(n_791),
.B(n_792),
.Y(n_960)
);

INVx4_ASAP7_75t_SL g961 ( 
.A(n_789),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_731),
.B(n_680),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_736),
.A2(n_799),
.B(n_787),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_821),
.B(n_827),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_816),
.A2(n_854),
.B1(n_868),
.B2(n_731),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_816),
.A2(n_868),
.B(n_854),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_739),
.B(n_400),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_816),
.A2(n_854),
.B1(n_868),
.B2(n_731),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_731),
.B(n_680),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_739),
.B(n_400),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_739),
.B(n_400),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_825),
.A2(n_838),
.B(n_832),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_731),
.B(n_680),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_826),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_825),
.A2(n_838),
.B(n_832),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_SL g976 ( 
.A1(n_772),
.A2(n_780),
.B(n_762),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_825),
.A2(n_838),
.B(n_832),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_828),
.B(n_587),
.Y(n_978)
);

OR2x6_ASAP7_75t_L g979 ( 
.A(n_826),
.B(n_660),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_731),
.B(n_680),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_731),
.B(n_680),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_731),
.B(n_680),
.Y(n_982)
);

HB1xp67_ASAP7_75t_SL g983 ( 
.A(n_831),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_731),
.B(n_680),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_760),
.B(n_775),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_731),
.B(n_680),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_877),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_884),
.B(n_964),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_898),
.A2(n_919),
.B1(n_904),
.B2(n_881),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_902),
.Y(n_990)
);

AND2x6_ASAP7_75t_L g991 ( 
.A(n_949),
.B(n_961),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_881),
.B(n_875),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_967),
.B(n_970),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_906),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_875),
.B(n_905),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_979),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_971),
.A2(n_888),
.B1(n_923),
.B2(n_912),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_983),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_878),
.A2(n_959),
.B(n_880),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_972),
.A2(n_977),
.B(n_975),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_SL g1001 ( 
.A1(n_950),
.A2(n_968),
.B1(n_965),
.B2(n_955),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_919),
.B(n_915),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_892),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_956),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_978),
.B(n_953),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_934),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_877),
.B(n_914),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_877),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_924),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_955),
.A2(n_966),
.B(n_876),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_924),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_R g1012 ( 
.A(n_887),
.B(n_899),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_929),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_894),
.A2(n_927),
.B(n_890),
.C(n_879),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_914),
.B(n_985),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_905),
.B(n_954),
.Y(n_1016)
);

BUFx4f_ASAP7_75t_L g1017 ( 
.A(n_974),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_954),
.B(n_962),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_SL g1019 ( 
.A1(n_965),
.A2(n_968),
.B1(n_966),
.B2(n_932),
.Y(n_1019)
);

NOR2x1_ASAP7_75t_R g1020 ( 
.A(n_882),
.B(n_914),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_SL g1021 ( 
.A1(n_876),
.A2(n_894),
.B1(n_957),
.B2(n_969),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_926),
.A2(n_920),
.B1(n_984),
.B2(n_962),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_958),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_969),
.B(n_973),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_SL g1025 ( 
.A1(n_886),
.A2(n_908),
.B(n_897),
.C(n_896),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_925),
.B(n_974),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_928),
.A2(n_986),
.B(n_982),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_883),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_907),
.B(n_889),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_973),
.B(n_980),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_907),
.B(n_901),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_938),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_943),
.B(n_980),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_925),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_981),
.B(n_982),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_981),
.B(n_921),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_921),
.B(n_885),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_936),
.B(n_976),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_896),
.A2(n_897),
.A3(n_903),
.B(n_922),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_893),
.A2(n_948),
.B1(n_936),
.B2(n_931),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_961),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_961),
.B(n_911),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_910),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_947),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_910),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_947),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_911),
.B(n_940),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_931),
.A2(n_886),
.B1(n_908),
.B2(n_916),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_947),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_913),
.B(n_946),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_910),
.Y(n_1051)
);

NOR2xp67_ASAP7_75t_L g1052 ( 
.A(n_935),
.B(n_945),
.Y(n_1052)
);

BUFx10_ASAP7_75t_L g1053 ( 
.A(n_910),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_933),
.Y(n_1054)
);

INVx5_ASAP7_75t_L g1055 ( 
.A(n_917),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_917),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_944),
.A2(n_960),
.B(n_952),
.C(n_900),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_941),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_942),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_937),
.A2(n_930),
.B(n_891),
.C(n_895),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_909),
.B(n_952),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_918),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_951),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_963),
.Y(n_1064)
);

OAI321xp33_ASAP7_75t_L g1065 ( 
.A1(n_884),
.A2(n_964),
.A3(n_763),
.B1(n_772),
.B2(n_968),
.C(n_965),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_939),
.Y(n_1066)
);

INVx3_ASAP7_75t_SL g1067 ( 
.A(n_983),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_878),
.A2(n_959),
.B(n_880),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_902),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_877),
.B(n_914),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_884),
.B(n_964),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_877),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_902),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_881),
.B(n_875),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_875),
.A2(n_884),
.B1(n_964),
.B2(n_731),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_961),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_983),
.B(n_831),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_875),
.A2(n_884),
.B1(n_964),
.B2(n_731),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_979),
.B(n_760),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_881),
.B(n_875),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_881),
.B(n_875),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_881),
.B(n_875),
.Y(n_1082)
);

AOI21xp33_ASAP7_75t_L g1083 ( 
.A1(n_884),
.A2(n_964),
.B(n_772),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_898),
.B(n_967),
.Y(n_1084)
);

AOI21xp33_ASAP7_75t_SL g1085 ( 
.A1(n_884),
.A2(n_964),
.B(n_753),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_887),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_979),
.B(n_826),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_892),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_902),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_979),
.B(n_760),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_881),
.B(n_875),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_898),
.B(n_967),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_898),
.B(n_967),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1017),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1019),
.B(n_1035),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1019),
.B(n_1001),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_988),
.A2(n_1071),
.B1(n_1078),
.B2(n_1075),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_990),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_SL g1099 ( 
.A(n_1006),
.Y(n_1099)
);

INVx5_ASAP7_75t_SL g1100 ( 
.A(n_1087),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1083),
.A2(n_1002),
.B1(n_1075),
.B2(n_1078),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1031),
.B(n_996),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_1003),
.Y(n_1103)
);

AND2x4_ASAP7_75t_SL g1104 ( 
.A(n_1053),
.B(n_1043),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_1077),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1083),
.A2(n_1002),
.B1(n_1021),
.B2(n_1030),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_1061),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1001),
.B(n_1033),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1018),
.A2(n_1037),
.B1(n_1031),
.B2(n_1022),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_999),
.A2(n_1068),
.B(n_1000),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1039),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1048),
.B(n_1036),
.Y(n_1112)
);

CKINVDCx6p67_ASAP7_75t_R g1113 ( 
.A(n_1067),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1009),
.B(n_1011),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1065),
.A2(n_997),
.B1(n_1081),
.B2(n_1082),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_1040),
.A2(n_1048),
.B1(n_1050),
.B2(n_1038),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1045),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_1039),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1040),
.A2(n_1038),
.B1(n_1024),
.B2(n_1080),
.Y(n_1119)
);

OAI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1065),
.A2(n_1080),
.B1(n_1074),
.B2(n_1082),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_SL g1121 ( 
.A1(n_1024),
.A2(n_1074),
.B1(n_1091),
.B2(n_1081),
.Y(n_1121)
);

INVx6_ASAP7_75t_L g1122 ( 
.A(n_1045),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_1084),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1091),
.A2(n_995),
.B1(n_1016),
.B2(n_1028),
.Y(n_1124)
);

CKINVDCx11_ASAP7_75t_R g1125 ( 
.A(n_998),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1069),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1013),
.Y(n_1127)
);

CKINVDCx11_ASAP7_75t_R g1128 ( 
.A(n_1086),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_1088),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1073),
.Y(n_1130)
);

CKINVDCx11_ASAP7_75t_R g1131 ( 
.A(n_1046),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1089),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1017),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1016),
.A2(n_1066),
.B1(n_991),
.B2(n_995),
.Y(n_1134)
);

BUFx2_ASAP7_75t_SL g1135 ( 
.A(n_1045),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1023),
.Y(n_1136)
);

BUFx2_ASAP7_75t_R g1137 ( 
.A(n_1056),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_996),
.B(n_1041),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1004),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_1092),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1013),
.B(n_994),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1010),
.A2(n_1093),
.B1(n_993),
.B2(n_989),
.Y(n_1142)
);

INVxp33_ASAP7_75t_L g1143 ( 
.A(n_1029),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_992),
.B(n_994),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1005),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_SL g1146 ( 
.A1(n_1066),
.A2(n_991),
.B1(n_1076),
.B2(n_1041),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1060),
.A2(n_1063),
.B(n_1027),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1059),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_1012),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1032),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1059),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1085),
.A2(n_1014),
.B1(n_1055),
.B2(n_1087),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1064),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1026),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1054),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1047),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1044),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_SL g1158 ( 
.A(n_1079),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1049),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1051),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1062),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1026),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1042),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1015),
.Y(n_1164)
);

BUFx4f_ASAP7_75t_SL g1165 ( 
.A(n_1034),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1042),
.A2(n_1090),
.B1(n_1079),
.B2(n_1053),
.Y(n_1166)
);

OA21x2_ASAP7_75t_L g1167 ( 
.A1(n_1052),
.A2(n_1025),
.B(n_1057),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1007),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1070),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1058),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_987),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1008),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1072),
.B(n_1020),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_988),
.A2(n_964),
.B1(n_884),
.B2(n_1071),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1019),
.B(n_1035),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_990),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1013),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_988),
.A2(n_964),
.B1(n_884),
.B2(n_1071),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_988),
.A2(n_964),
.B1(n_884),
.B2(n_1071),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1017),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_SL g1181 ( 
.A1(n_988),
.A2(n_1071),
.B1(n_884),
.B2(n_964),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_988),
.A2(n_1071),
.B1(n_1078),
.B2(n_1075),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1107),
.B(n_1111),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1153),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1153),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1138),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1111),
.Y(n_1187)
);

BUFx12f_ASAP7_75t_L g1188 ( 
.A(n_1125),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1118),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1107),
.B(n_1118),
.Y(n_1190)
);

NAND3xp33_ASAP7_75t_L g1191 ( 
.A(n_1178),
.B(n_1097),
.C(n_1174),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1096),
.A2(n_1181),
.B1(n_1182),
.B2(n_1101),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1110),
.A2(n_1152),
.B(n_1167),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1112),
.B(n_1095),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1147),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1151),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1147),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1096),
.B(n_1095),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1147),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1175),
.B(n_1108),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1167),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1098),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_1120),
.A2(n_1115),
.B(n_1124),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1175),
.B(n_1108),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1102),
.B(n_1161),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1148),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1121),
.B(n_1112),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1148),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1141),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1126),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1130),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1114),
.B(n_1132),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1171),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1176),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1141),
.B(n_1144),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1114),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1136),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1127),
.Y(n_1218)
);

AO21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1106),
.A2(n_1160),
.B(n_1109),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1135),
.B(n_1122),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1177),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1139),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1119),
.B(n_1116),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1125),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1142),
.B(n_1123),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1150),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1172),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1155),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1179),
.B(n_1103),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1140),
.B(n_1134),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1145),
.B(n_1163),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1156),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1146),
.B(n_1100),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1129),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1099),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1193),
.A2(n_1157),
.B(n_1159),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1195),
.B(n_1143),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1195),
.B(n_1143),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1185),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1195),
.B(n_1163),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1223),
.A2(n_1129),
.B1(n_1158),
.B2(n_1162),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1185),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1197),
.B(n_1168),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1207),
.B(n_1117),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1220),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1197),
.B(n_1168),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1206),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_R g1248 ( 
.A(n_1224),
.B(n_1149),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1202),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1196),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1223),
.A2(n_1158),
.B1(n_1154),
.B2(n_1162),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1199),
.B(n_1113),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1184),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1199),
.B(n_1113),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1199),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1199),
.B(n_1131),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1186),
.B(n_1104),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1216),
.B(n_1212),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1224),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1191),
.B(n_1131),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1216),
.B(n_1128),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1212),
.B(n_1128),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1201),
.B(n_1170),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1212),
.B(n_1169),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1184),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1213),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1207),
.B(n_1169),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1194),
.B(n_1173),
.Y(n_1268)
);

NAND2x1_ASAP7_75t_L g1269 ( 
.A(n_1220),
.B(n_1166),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1194),
.B(n_1164),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1184),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1258),
.B(n_1183),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1258),
.B(n_1183),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1239),
.B(n_1218),
.Y(n_1274)
);

AOI221xp5_ASAP7_75t_L g1275 ( 
.A1(n_1260),
.A2(n_1223),
.B1(n_1198),
.B2(n_1191),
.C(n_1200),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1239),
.B(n_1218),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_L g1277 ( 
.A(n_1260),
.B(n_1192),
.C(n_1229),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1244),
.B(n_1192),
.C(n_1229),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1241),
.A2(n_1198),
.B1(n_1188),
.B2(n_1200),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1242),
.B(n_1221),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1259),
.B(n_1188),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1242),
.B(n_1221),
.Y(n_1282)
);

AND2x2_ASAP7_75t_SL g1283 ( 
.A(n_1245),
.B(n_1187),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1237),
.B(n_1190),
.Y(n_1284)
);

NAND3xp33_ASAP7_75t_L g1285 ( 
.A(n_1244),
.B(n_1226),
.C(n_1210),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1253),
.B(n_1226),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1247),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1253),
.B(n_1209),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1253),
.B(n_1209),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1265),
.B(n_1210),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1248),
.B(n_1188),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1262),
.A2(n_1198),
.B(n_1204),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1247),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1267),
.A2(n_1203),
.B1(n_1219),
.B2(n_1225),
.Y(n_1294)
);

NAND3xp33_ASAP7_75t_L g1295 ( 
.A(n_1267),
.B(n_1228),
.C(n_1211),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1252),
.B(n_1228),
.C(n_1214),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1265),
.B(n_1204),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1248),
.B(n_1234),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1259),
.A2(n_1149),
.B1(n_1235),
.B2(n_1234),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1271),
.B(n_1204),
.Y(n_1300)
);

NAND3xp33_ASAP7_75t_L g1301 ( 
.A(n_1252),
.B(n_1208),
.C(n_1189),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1262),
.A2(n_1246),
.B(n_1243),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1257),
.A2(n_1203),
.B(n_1158),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1237),
.B(n_1238),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1238),
.B(n_1190),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1262),
.A2(n_1230),
.B(n_1234),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_L g1307 ( 
.A(n_1252),
.B(n_1214),
.C(n_1217),
.Y(n_1307)
);

OA211x2_ASAP7_75t_L g1308 ( 
.A1(n_1269),
.A2(n_1208),
.B(n_1233),
.C(n_1203),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1256),
.B(n_1230),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1240),
.B(n_1205),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1254),
.B(n_1217),
.C(n_1227),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1269),
.A2(n_1233),
.B1(n_1230),
.B2(n_1220),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1256),
.B(n_1235),
.Y(n_1313)
);

AOI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1270),
.A2(n_1203),
.B1(n_1225),
.B2(n_1232),
.C(n_1222),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1240),
.B(n_1205),
.Y(n_1315)
);

OAI221xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1241),
.A2(n_1187),
.B1(n_1203),
.B2(n_1231),
.C(n_1225),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1240),
.B(n_1205),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1287),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1304),
.B(n_1255),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1274),
.B(n_1270),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1281),
.B(n_1261),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1311),
.B(n_1245),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1293),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1276),
.B(n_1266),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1272),
.B(n_1256),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1280),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1293),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1284),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1282),
.B(n_1266),
.Y(n_1329)
);

AND2x2_ASAP7_75t_SL g1330 ( 
.A(n_1283),
.B(n_1245),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1284),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1272),
.B(n_1243),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1310),
.B(n_1245),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1273),
.B(n_1243),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1310),
.B(n_1245),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1311),
.B(n_1246),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1283),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1295),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1295),
.B(n_1250),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1273),
.B(n_1246),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1285),
.B(n_1250),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_SL g1342 ( 
.A(n_1316),
.B(n_1254),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1290),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1283),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1286),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1314),
.B(n_1250),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1296),
.B(n_1307),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1299),
.B(n_1291),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1296),
.B(n_1249),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1297),
.B(n_1300),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1315),
.B(n_1254),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1288),
.B(n_1215),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1289),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1305),
.B(n_1264),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1338),
.B(n_1278),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1338),
.B(n_1292),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1347),
.B(n_1326),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1347),
.B(n_1306),
.Y(n_1358)
);

AOI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1346),
.A2(n_1277),
.B1(n_1275),
.B2(n_1312),
.C(n_1294),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1328),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1339),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1348),
.B(n_1299),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1339),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1326),
.B(n_1307),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1349),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1344),
.B(n_1315),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1328),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1328),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1343),
.B(n_1277),
.Y(n_1369)
);

NOR2x1_ASAP7_75t_L g1370 ( 
.A(n_1337),
.B(n_1298),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1331),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1321),
.B(n_1302),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1349),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1353),
.B(n_1261),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1341),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1341),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1342),
.B(n_1301),
.C(n_1279),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1343),
.B(n_1249),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1352),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1331),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1344),
.B(n_1317),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1320),
.B(n_1309),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1318),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1318),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1346),
.Y(n_1385)
);

AOI21xp33_ASAP7_75t_L g1386 ( 
.A1(n_1342),
.A2(n_1236),
.B(n_1268),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1352),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1320),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1337),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1330),
.B(n_1269),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1337),
.B(n_1317),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1345),
.B(n_1236),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1364),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1355),
.B(n_1345),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1383),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1383),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1377),
.A2(n_1337),
.B1(n_1330),
.B2(n_1336),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1362),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1365),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1389),
.B(n_1336),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1391),
.B(n_1332),
.Y(n_1401)
);

NOR2x1_ASAP7_75t_L g1402 ( 
.A(n_1370),
.B(n_1336),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1391),
.B(n_1332),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1384),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1369),
.B(n_1323),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1384),
.Y(n_1406)
);

NAND4xp25_ASAP7_75t_L g1407 ( 
.A(n_1358),
.B(n_1261),
.C(n_1336),
.D(n_1308),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1378),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1379),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1366),
.B(n_1332),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1385),
.A2(n_1303),
.B(n_1322),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1364),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1365),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1366),
.B(n_1334),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1387),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1388),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1361),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1361),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1360),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1363),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1363),
.Y(n_1421)
);

OAI31xp33_ASAP7_75t_L g1422 ( 
.A1(n_1386),
.A2(n_1322),
.A3(n_1308),
.B(n_1353),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1357),
.B(n_1323),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1375),
.B(n_1323),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1373),
.B(n_1327),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1376),
.B(n_1327),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1381),
.B(n_1334),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1376),
.Y(n_1428)
);

OAI211xp5_ASAP7_75t_L g1429 ( 
.A1(n_1358),
.A2(n_1303),
.B(n_1327),
.C(n_1313),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1356),
.B(n_1359),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1382),
.B(n_1350),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1382),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1374),
.B(n_1319),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1360),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1389),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1410),
.B(n_1389),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1398),
.A2(n_1372),
.B(n_1390),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1432),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1430),
.B(n_1381),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1393),
.A2(n_1219),
.B1(n_1390),
.B2(n_1392),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1395),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1395),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1396),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1394),
.B(n_1367),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1402),
.B(n_1322),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1396),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1404),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1404),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1431),
.B(n_1367),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1394),
.B(n_1368),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1405),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1431),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1402),
.A2(n_1397),
.B1(n_1429),
.B2(n_1400),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1410),
.B(n_1334),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1406),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1405),
.B(n_1368),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1419),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1406),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1393),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1407),
.A2(n_1390),
.B(n_1392),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1416),
.B(n_1371),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1416),
.B(n_1371),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1409),
.B(n_1380),
.Y(n_1463)
);

NOR2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1435),
.B(n_1322),
.Y(n_1464)
);

AND2x4_ASAP7_75t_SL g1465 ( 
.A(n_1409),
.B(n_1333),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1414),
.B(n_1340),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1415),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1415),
.B(n_1380),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1399),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1413),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1412),
.A2(n_1434),
.B(n_1419),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_L g1472 ( 
.A(n_1439),
.B(n_1418),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1438),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1441),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1471),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1443),
.Y(n_1478)
);

AO21x1_ASAP7_75t_L g1479 ( 
.A1(n_1453),
.A2(n_1428),
.B(n_1420),
.Y(n_1479)
);

AOI222xp33_ASAP7_75t_L g1480 ( 
.A1(n_1459),
.A2(n_1412),
.B1(n_1411),
.B2(n_1428),
.C1(n_1420),
.C2(n_1421),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1440),
.A2(n_1422),
.B1(n_1434),
.B2(n_1219),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1446),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1450),
.B(n_1408),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1469),
.B(n_1433),
.Y(n_1485)
);

AOI21xp33_ASAP7_75t_L g1486 ( 
.A1(n_1444),
.A2(n_1421),
.B(n_1417),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1447),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1440),
.A2(n_1417),
.B1(n_1408),
.B2(n_1425),
.Y(n_1488)
);

OAI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1460),
.A2(n_1423),
.B1(n_1426),
.B2(n_1424),
.C(n_1251),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1436),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1454),
.B(n_1414),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1471),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1449),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1444),
.B(n_1427),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1456),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1437),
.A2(n_1423),
.B(n_1424),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1490),
.B(n_1470),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1475),
.B(n_1495),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1479),
.B(n_1467),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1495),
.B(n_1454),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1493),
.B(n_1466),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_R g1502 ( 
.A1(n_1479),
.A2(n_1457),
.B1(n_1448),
.B2(n_1455),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1472),
.A2(n_1457),
.B1(n_1445),
.B2(n_1462),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1493),
.B(n_1466),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1483),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1485),
.B(n_1427),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1472),
.A2(n_1445),
.B1(n_1461),
.B2(n_1456),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1476),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1491),
.Y(n_1509)
);

AND2x2_ASAP7_75t_SL g1510 ( 
.A(n_1481),
.B(n_1445),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1491),
.B(n_1436),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1476),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1473),
.Y(n_1513)
);

INVxp33_ASAP7_75t_L g1514 ( 
.A(n_1494),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1484),
.B(n_1458),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_L g1516 ( 
.A(n_1499),
.B(n_1486),
.C(n_1477),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1501),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1504),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1499),
.A2(n_1496),
.B(n_1480),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1508),
.A2(n_1492),
.B(n_1477),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1502),
.B(n_1488),
.C(n_1492),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_SL g1522 ( 
.A1(n_1512),
.A2(n_1474),
.B(n_1487),
.C(n_1478),
.Y(n_1522)
);

NOR4xp25_ASAP7_75t_L g1523 ( 
.A(n_1505),
.B(n_1482),
.C(n_1489),
.D(n_1484),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1500),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1498),
.A2(n_1468),
.B(n_1463),
.C(n_1464),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1509),
.B(n_1401),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_SL g1527 ( 
.A(n_1519),
.B(n_1523),
.C(n_1516),
.Y(n_1527)
);

NAND4xp25_ASAP7_75t_L g1528 ( 
.A(n_1522),
.B(n_1503),
.C(n_1507),
.D(n_1497),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1520),
.Y(n_1529)
);

AOI22x1_ASAP7_75t_L g1530 ( 
.A1(n_1517),
.A2(n_1513),
.B1(n_1514),
.B2(n_1403),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1520),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1521),
.B(n_1515),
.C(n_1506),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1518),
.B(n_1511),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1526),
.B(n_1510),
.Y(n_1534)
);

XOR2x2_ASAP7_75t_L g1535 ( 
.A(n_1524),
.B(n_1510),
.Y(n_1535)
);

NAND4xp25_ASAP7_75t_SL g1536 ( 
.A(n_1525),
.B(n_1403),
.C(n_1401),
.D(n_1463),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1534),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_L g1538 ( 
.A(n_1527),
.B(n_1468),
.Y(n_1538)
);

NOR3xp33_ASAP7_75t_L g1539 ( 
.A(n_1528),
.B(n_1105),
.C(n_1094),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1529),
.A2(n_1465),
.B1(n_1330),
.B2(n_1236),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1531),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1535),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1538),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1537),
.B(n_1533),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1542),
.B(n_1532),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1539),
.A2(n_1528),
.B1(n_1541),
.B2(n_1536),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1540),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1538),
.A2(n_1465),
.B1(n_1530),
.B2(n_1165),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1544),
.B(n_1354),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1543),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1545),
.B(n_1340),
.Y(n_1551)
);

NOR2xp67_ASAP7_75t_L g1552 ( 
.A(n_1548),
.B(n_1324),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1547),
.A2(n_1170),
.B1(n_1236),
.B2(n_1335),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1549),
.B(n_1546),
.Y(n_1554)
);

NAND3x1_ASAP7_75t_L g1555 ( 
.A(n_1550),
.B(n_1340),
.C(n_1325),
.Y(n_1555)
);

NOR3xp33_ASAP7_75t_L g1556 ( 
.A(n_1552),
.B(n_1133),
.C(n_1094),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1555),
.Y(n_1557)
);

NOR3xp33_ASAP7_75t_L g1558 ( 
.A(n_1557),
.B(n_1554),
.C(n_1556),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1558),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1558),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1559),
.A2(n_1557),
.B(n_1560),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1559),
.Y(n_1562)
);

XOR2xp5_ASAP7_75t_L g1563 ( 
.A(n_1562),
.B(n_1551),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1561),
.A2(n_1553),
.B(n_1180),
.Y(n_1564)
);

AOI21xp33_ASAP7_75t_L g1565 ( 
.A1(n_1563),
.A2(n_1180),
.B(n_1133),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1565),
.Y(n_1566)
);

AOI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1566),
.A2(n_1564),
.B1(n_1325),
.B2(n_1236),
.C(n_1351),
.Y(n_1567)
);

AOI211xp5_ASAP7_75t_L g1568 ( 
.A1(n_1567),
.A2(n_1263),
.B(n_1137),
.C(n_1329),
.Y(n_1568)
);


endmodule