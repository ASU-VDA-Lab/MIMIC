module real_jpeg_25700_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_0),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_0),
.A2(n_36),
.B1(n_69),
.B2(n_71),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_0),
.A2(n_22),
.B1(n_27),
.B2(n_36),
.Y(n_158)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_2),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_2),
.B(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_2),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_33),
.B1(n_37),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_22),
.B1(n_27),
.B2(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_3),
.A2(n_69),
.B1(n_71),
.B2(n_84),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_84),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_4),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_69),
.B1(n_71),
.B2(n_99),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_33),
.B1(n_43),
.B2(n_99),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_99),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_7),
.A2(n_32),
.B1(n_44),
.B2(n_68),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_178)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_31),
.B1(n_37),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_9),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_121),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_9),
.A2(n_69),
.B1(n_71),
.B2(n_121),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_121),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_11),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_11),
.B(n_21),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_69),
.C(n_95),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_11),
.B(n_136),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_11),
.A2(n_69),
.B1(n_71),
.B2(n_224),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_11),
.B(n_57),
.C(n_74),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_11),
.A2(n_56),
.B(n_284),
.Y(n_312)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_13),
.A2(n_38),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_13),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_13),
.A2(n_22),
.B1(n_27),
.B2(n_88),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_13),
.A2(n_69),
.B1(n_71),
.B2(n_88),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_88),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_15),
.A2(n_32),
.B1(n_38),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_15),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_15),
.A2(n_22),
.B1(n_27),
.B2(n_170),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_15),
.A2(n_69),
.B1(n_71),
.B2(n_170),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_170),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_16),
.A2(n_42),
.B1(n_69),
.B2(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_16),
.A2(n_42),
.B1(n_57),
.B2(n_58),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_16),
.A2(n_22),
.B1(n_27),
.B2(n_42),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_48),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_29),
.B(n_35),
.Y(n_20)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_21),
.A2(n_29),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_21),
.A2(n_29),
.B1(n_120),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_21),
.A2(n_29),
.B1(n_41),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_21)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_22),
.A2(n_27),
.B1(n_95),
.B2(n_96),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g196 ( 
.A(n_22),
.B(n_28),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_22),
.B(n_249),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_25),
.A2(n_27),
.A3(n_32),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_29),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_29),
.A2(n_124),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_32),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_34),
.A2(n_83),
.B(n_85),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_34),
.B(n_87),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_34),
.A2(n_83),
.B1(n_122),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_34),
.A2(n_122),
.B1(n_144),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_34),
.A2(n_85),
.B(n_187),
.Y(n_186)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_40),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_40),
.B(n_359),
.Y(n_360)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_358),
.B(n_360),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_346),
.B(n_357),
.Y(n_49)
);

OAI31xp33_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_146),
.A3(n_160),
.B(n_343),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_125),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_52),
.B(n_125),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_90),
.C(n_106),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_53),
.A2(n_90),
.B1(n_91),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_53),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_79),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_54),
.A2(n_55),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_55),
.A2(n_65),
.B1(n_66),
.B2(n_80),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_61),
.B(n_64),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_56),
.A2(n_61),
.B1(n_64),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_56),
.A2(n_111),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_56),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_56),
.A2(n_200),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_56),
.B(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_56),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_58),
.B(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_63),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_72),
.B1(n_78),
.B2(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_69),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_71),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_69),
.B(n_291),
.Y(n_290)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_72),
.A2(n_78),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_72),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_72),
.A2(n_78),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_76),
.A2(n_102),
.B1(n_115),
.B2(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_76),
.A2(n_182),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_76),
.A2(n_220),
.B(n_257),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_76),
.B(n_224),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_78),
.B(n_221),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_101),
.B(n_105),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_100),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_93),
.A2(n_94),
.B1(n_138),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_93),
.A2(n_189),
.B(n_191),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_93),
.A2(n_191),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_94),
.A2(n_117),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_94),
.A2(n_173),
.B(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_102),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_102),
.A2(n_272),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_106),
.A2(n_107),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.C(n_118),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_108),
.A2(n_109),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_116),
.B(n_118),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B(n_123),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_128),
.C(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_143),
.B2(n_145),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_140),
.C(n_143),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_135),
.A2(n_136),
.B1(n_190),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_135),
.A2(n_136),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_136),
.B(n_174),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_140),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_140),
.B(n_153),
.C(n_157),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_143),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_145),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_143),
.B(n_149),
.C(n_152),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_147),
.A2(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_159),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_148),
.B(n_159),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_154),
.Y(n_353)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_158),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_336),
.B(n_342),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_209),
.B(n_335),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_202),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_163),
.B(n_202),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_183),
.C(n_185),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_164),
.A2(n_165),
.B1(n_183),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_171),
.C(n_175),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_176),
.B(n_181),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_197)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_183),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_185),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_192),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_188),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_197),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_198),
.A2(n_295),
.B1(n_297),
.B2(n_299),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_204),
.B(n_205),
.C(n_208),
.Y(n_341)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_241),
.B(n_329),
.C(n_334),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_235),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_226),
.C(n_227),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_212),
.A2(n_213),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_218),
.C(n_222),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_224),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_226),
.B(n_227),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_234),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_323),
.B(n_328),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_273),
.B(n_322),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_262),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_246),
.B(n_262),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.C(n_259),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_250),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B(n_253),
.Y(n_250)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_255),
.A2(n_259),
.B1(n_260),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_269),
.C(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_316),
.B(n_321),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_292),
.B(n_315),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_286),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_290),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_302),
.B(n_314),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_300),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_300),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_308),
.B(n_313),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_341),
.Y(n_342)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_348),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_356),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_350),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_352),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_354),
.C(n_356),
.Y(n_359)
);


endmodule