module fake_netlist_5_1252_n_448 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_448);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_448;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_136;
wire n_315;
wire n_268;
wire n_408;
wire n_376;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_397;
wire n_155;
wire n_423;
wire n_284;
wire n_245;
wire n_139;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_417;
wire n_385;
wire n_212;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_209;
wire n_259;
wire n_375;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_325;
wire n_132;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_387;
wire n_374;
wire n_276;
wire n_163;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_344;
wire n_287;
wire n_422;
wire n_415;
wire n_141;
wire n_355;
wire n_336;
wire n_145;
wire n_337;
wire n_430;
wire n_313;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_213;
wire n_342;
wire n_361;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_277;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_239;
wire n_420;
wire n_310;
wire n_358;
wire n_362;
wire n_332;
wire n_170;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_441;
wire n_312;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_143;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_437;
wire n_177;
wire n_403;
wire n_421;
wire n_405;
wire n_359;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_410;
wire n_269;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_135;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_29),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_2),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_31),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_10),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_6),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g148 ( 
.A(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_48),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_19),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_56),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_55),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_102),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_17),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_40),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_25),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_3),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_39),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_65),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_90),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_38),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_42),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_73),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_87),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_16),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_51),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_28),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_24),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_4),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_15),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_59),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_71),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_62),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_74),
.B(n_107),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_43),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_13),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_11),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_37),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_7),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_49),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_81),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_0),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_61),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_86),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_111),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_85),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_100),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_124),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_58),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_130),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_115),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_20),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_41),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_126),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_97),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_12),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_69),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_121),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_32),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g236 ( 
.A(n_114),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_54),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_104),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_78),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_35),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_70),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_133),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_0),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_134),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_135),
.B(n_1),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

NAND2xp33_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_8),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_181),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_132),
.B(n_22),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_177),
.B(n_23),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_141),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_138),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_142),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_145),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_164),
.B(n_36),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_146),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_147),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_149),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_150),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_151),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_152),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_44),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_155),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_156),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_157),
.B(n_158),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_180),
.B(n_45),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_160),
.B(n_46),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_191),
.B(n_47),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_161),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_165),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_168),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_169),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_185),
.B(n_50),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_173),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g286 ( 
.A(n_144),
.B(n_52),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_213),
.A2(n_53),
.B(n_63),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_174),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_175),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_179),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_182),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_184),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_186),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_252),
.B(n_197),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_250),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_273),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_187),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_257),
.B(n_189),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_270),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_207),
.B1(n_237),
.B2(n_236),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_245),
.B(n_166),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_143),
.C(n_228),
.Y(n_310)
);

AO22x2_ASAP7_75t_L g311 ( 
.A1(n_255),
.A2(n_214),
.B1(n_239),
.B2(n_238),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_148),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_SL g313 ( 
.A(n_253),
.B(n_154),
.C(n_172),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_188),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

BUFx6f_ASAP7_75t_SL g317 ( 
.A(n_286),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_203),
.B1(n_218),
.B2(n_176),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_274),
.B(n_163),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_243),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_316),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_221),
.B1(n_171),
.B2(n_196),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_317),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_224),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_244),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_246),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_297),
.A2(n_249),
.B1(n_286),
.B2(n_194),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_295),
.B(n_294),
.C(n_291),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_283),
.B1(n_223),
.B2(n_226),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_140),
.B1(n_202),
.B2(n_136),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_248),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_251),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_306),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_288),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_333),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_328),
.A2(n_311),
.B1(n_193),
.B2(n_162),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_311),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_298),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_315),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_302),
.Y(n_355)
);

INVx6_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_344),
.A2(n_241),
.B(n_323),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_347),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_266),
.C(n_254),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_SL g360 ( 
.A1(n_340),
.A2(n_209),
.B(n_208),
.C(n_206),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_342),
.A2(n_195),
.B1(n_190),
.B2(n_178),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_319),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_336),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_346),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_329),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_363),
.A2(n_338),
.B(n_287),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_352),
.Y(n_369)
);

BUFx8_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_353),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_327),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_331),
.B1(n_345),
.B2(n_211),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_366),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_361),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_305),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

AND2x4_ASAP7_75t_SL g383 ( 
.A(n_369),
.B(n_367),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_371),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_348),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_350),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_359),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_377),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_375),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_357),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_378),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_324),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_368),
.B(n_234),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_384),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_394),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_387),
.A2(n_362),
.B1(n_381),
.B2(n_269),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_390),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_382),
.Y(n_400)
);

AOI21xp33_ASAP7_75t_SL g401 ( 
.A1(n_385),
.A2(n_170),
.B(n_284),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

AO21x2_ASAP7_75t_L g403 ( 
.A1(n_387),
.A2(n_360),
.B(n_200),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_388),
.A2(n_199),
.B1(n_233),
.B2(n_232),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

OAI221xp5_ASAP7_75t_L g407 ( 
.A1(n_389),
.A2(n_230),
.B1(n_201),
.B2(n_212),
.C(n_215),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_400),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_404),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_406),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_383),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_282),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_198),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_397),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_412),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_410),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_411),
.B(n_397),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_409),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_398),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_419),
.B(n_417),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_407),
.C(n_414),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_420),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_418),
.A2(n_395),
.B(n_403),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_418),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_415),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_413),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_217),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_426),
.B(n_401),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_427),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_219),
.Y(n_431)
);

AOI221xp5_ASAP7_75t_SL g432 ( 
.A1(n_431),
.A2(n_425),
.B1(n_220),
.B2(n_227),
.C(n_229),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_422),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_66),
.Y(n_434)
);

AOI211xp5_ASAP7_75t_L g435 ( 
.A1(n_433),
.A2(n_432),
.B(n_434),
.C(n_428),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_424),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_436),
.Y(n_437)
);

OAI22x1_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_281),
.B1(n_280),
.B2(n_271),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_436),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_SL g440 ( 
.A(n_437),
.B(n_439),
.C(n_438),
.Y(n_440)
);

AOI221x1_ASAP7_75t_L g441 ( 
.A1(n_437),
.A2(n_260),
.B1(n_267),
.B2(n_265),
.C(n_264),
.Y(n_441)
);

NOR3xp33_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_231),
.C(n_225),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

NAND5xp2_ASAP7_75t_L g444 ( 
.A(n_442),
.B(n_222),
.C(n_256),
.D(n_72),
.E(n_75),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_440),
.Y(n_445)
);

OAI221xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_262),
.B1(n_259),
.B2(n_76),
.C(n_84),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_447),
.A2(n_443),
.B(n_444),
.Y(n_448)
);


endmodule