module real_aes_4235_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_0), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g49 ( .A(n_1), .Y(n_49) );
CKINVDCx5p33_ASAP7_75t_R g47 ( .A(n_2), .Y(n_47) );
NOR2xp33_ASAP7_75t_R g27 ( .A(n_3), .B(n_7), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_3), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g23 ( .A(n_4), .B(n_24), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_5), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_6), .Y(n_22) );
NOR4xp25_ASAP7_75t_SL g30 ( .A(n_6), .B(n_21), .C(n_31), .D(n_33), .Y(n_30) );
NAND2xp33_ASAP7_75t_R g43 ( .A(n_6), .B(n_23), .Y(n_43) );
NAND2xp33_ASAP7_75t_R g29 ( .A(n_7), .B(n_30), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g38 ( .A(n_7), .Y(n_38) );
NOR2xp33_ASAP7_75t_R g40 ( .A(n_7), .B(n_41), .Y(n_40) );
NAND2xp33_ASAP7_75t_R g46 ( .A(n_7), .B(n_42), .Y(n_46) );
NAND3xp33_ASAP7_75t_SL g48 ( .A(n_7), .B(n_18), .C(n_33), .Y(n_48) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_8), .Y(n_34) );
NAND3xp33_ASAP7_75t_SL g24 ( .A(n_9), .B(n_25), .C(n_26), .Y(n_24) );
AOI221xp5_ASAP7_75t_R g35 ( .A1(n_10), .A2(n_15), .B1(n_36), .B2(n_39), .C(n_45), .Y(n_35) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_11), .B(n_19), .C(n_20), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_11), .B(n_12), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_12), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_13), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_14), .Y(n_26) );
OAI221xp5_ASAP7_75t_R g16 ( .A1(n_17), .A2(n_28), .B1(n_29), .B2(n_34), .C(n_35), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_18), .B(n_27), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g20 ( .A(n_21), .B(n_22), .C(n_23), .Y(n_20) );
NOR4xp25_ASAP7_75t_SL g42 ( .A(n_21), .B(n_33), .C(n_43), .D(n_44), .Y(n_42) );
NAND2xp33_ASAP7_75t_R g31 ( .A(n_23), .B(n_32), .Y(n_31) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_30), .B(n_38), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g44 ( .A(n_32), .Y(n_44) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
HB1xp67_ASAP7_75t_L g39 ( .A(n_40), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g41 ( .A(n_42), .Y(n_41) );
OAI22xp33_ASAP7_75t_L g45 ( .A1(n_46), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_45) );
endmodule