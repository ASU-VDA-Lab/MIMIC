module real_aes_6646_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g232 ( .A1(n_0), .A2(n_233), .B(n_234), .C(n_238), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_1), .B(n_174), .Y(n_239) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g457 ( .A(n_2), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_3), .B(n_146), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_4), .A2(n_132), .B(n_137), .C(n_501), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_5), .A2(n_127), .B(n_539), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_6), .A2(n_127), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_7), .B(n_174), .Y(n_545) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_8), .A2(n_162), .B(n_178), .Y(n_177) );
AND2x6_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_10), .A2(n_132), .B(n_137), .C(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g483 ( .A(n_11), .Y(n_483) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_12), .B(n_40), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_13), .B(n_237), .Y(n_503) );
INVx1_ASAP7_75t_L g156 ( .A(n_14), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_15), .B(n_146), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_16), .A2(n_147), .B(n_491), .C(n_493), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_17), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_18), .B(n_174), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_19), .B(n_211), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_20), .A2(n_137), .B(n_188), .C(n_207), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_21), .A2(n_186), .B(n_236), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_22), .B(n_237), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_23), .B(n_237), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_24), .Y(n_530) );
INVx1_ASAP7_75t_L g522 ( .A(n_25), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_26), .A2(n_137), .B(n_181), .C(n_188), .Y(n_180) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_27), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_28), .Y(n_499) );
INVx1_ASAP7_75t_L g579 ( .A(n_29), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_30), .A2(n_127), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g130 ( .A(n_31), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_32), .A2(n_135), .B(n_150), .C(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_33), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_34), .A2(n_236), .B(n_542), .C(n_544), .Y(n_541) );
INVxp67_ASAP7_75t_L g580 ( .A(n_35), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_36), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_37), .A2(n_137), .B(n_188), .C(n_521), .Y(n_520) );
CKINVDCx14_ASAP7_75t_R g540 ( .A(n_38), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_39), .A2(n_98), .B1(n_465), .B2(n_742), .C1(n_743), .C2(n_746), .Y(n_464) );
INVx1_ASAP7_75t_L g742 ( .A(n_39), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_40), .B(n_105), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_41), .A2(n_238), .B(n_481), .C(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_42), .B(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_43), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_44), .A2(n_119), .B1(n_120), .B2(n_450), .Y(n_118) );
INVx1_ASAP7_75t_L g450 ( .A(n_44), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_45), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_46), .B(n_127), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_47), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_48), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_49), .A2(n_135), .B(n_140), .C(n_150), .Y(n_134) );
INVx1_ASAP7_75t_L g235 ( .A(n_50), .Y(n_235) );
INVx1_ASAP7_75t_L g141 ( .A(n_51), .Y(n_141) );
INVx1_ASAP7_75t_L g511 ( .A(n_52), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_53), .B(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_54), .Y(n_214) );
CKINVDCx14_ASAP7_75t_R g479 ( .A(n_55), .Y(n_479) );
INVx1_ASAP7_75t_L g133 ( .A(n_56), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_57), .B(n_127), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_58), .B(n_174), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_59), .A2(n_168), .B(n_170), .C(n_172), .Y(n_167) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
INVx1_ASAP7_75t_SL g543 ( .A(n_61), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_62), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_63), .B(n_146), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_64), .B(n_174), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_65), .B(n_147), .Y(n_249) );
INVx1_ASAP7_75t_L g533 ( .A(n_66), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_67), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_68), .B(n_143), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_69), .A2(n_137), .B(n_150), .C(n_220), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g166 ( .A(n_70), .Y(n_166) );
INVx1_ASAP7_75t_L g111 ( .A(n_71), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_72), .A2(n_127), .B(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_73), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_74), .A2(n_127), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_75), .A2(n_205), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g489 ( .A(n_76), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_77), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_78), .B(n_142), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_79), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_80), .A2(n_127), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g492 ( .A(n_81), .Y(n_492) );
INVx2_ASAP7_75t_L g153 ( .A(n_82), .Y(n_153) );
INVx1_ASAP7_75t_L g502 ( .A(n_83), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_84), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_85), .B(n_237), .Y(n_250) );
INVx2_ASAP7_75t_L g108 ( .A(n_86), .Y(n_108) );
OR2x2_ASAP7_75t_L g454 ( .A(n_86), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g741 ( .A(n_86), .B(n_456), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_87), .A2(n_137), .B(n_150), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_88), .B(n_127), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_89), .Y(n_197) );
INVxp67_ASAP7_75t_L g171 ( .A(n_90), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_91), .B(n_162), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_92), .A2(n_100), .B1(n_112), .B2(n_750), .Y(n_99) );
INVx2_ASAP7_75t_L g514 ( .A(n_93), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_94), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g221 ( .A(n_95), .Y(n_221) );
INVx1_ASAP7_75t_L g245 ( .A(n_96), .Y(n_245) );
AND2x2_ASAP7_75t_L g157 ( .A(n_97), .B(n_152), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g750 ( .A(n_102), .Y(n_750) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g470 ( .A(n_108), .B(n_456), .Y(n_470) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_108), .B(n_455), .Y(n_745) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_463), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g749 ( .A(n_116), .Y(n_749) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_451), .B(n_459), .Y(n_117) );
AOI22x1_ASAP7_75t_SL g747 ( .A1(n_119), .A2(n_467), .B1(n_738), .B2(n_748), .Y(n_747) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_120), .A2(n_467), .B1(n_471), .B2(n_738), .Y(n_466) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR5x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_323), .C(n_401), .D(n_425), .E(n_442), .Y(n_121) );
OAI211xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_189), .B(n_240), .C(n_300), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_158), .Y(n_123) );
AND2x2_ASAP7_75t_L g254 ( .A(n_124), .B(n_160), .Y(n_254) );
INVx5_ASAP7_75t_SL g282 ( .A(n_124), .Y(n_282) );
AND2x2_ASAP7_75t_L g318 ( .A(n_124), .B(n_303), .Y(n_318) );
OR2x2_ASAP7_75t_L g357 ( .A(n_124), .B(n_159), .Y(n_357) );
OR2x2_ASAP7_75t_L g388 ( .A(n_124), .B(n_279), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_124), .B(n_292), .Y(n_424) );
AND2x2_ASAP7_75t_L g436 ( .A(n_124), .B(n_279), .Y(n_436) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_157), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_134), .B(n_152), .Y(n_125) );
BUFx2_ASAP7_75t_L g205 ( .A(n_127), .Y(n_205) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_128), .B(n_132), .Y(n_246) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
INVx1_ASAP7_75t_L g187 ( .A(n_130), .Y(n_187) );
INVx1_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
INVx3_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
INVx1_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_131), .Y(n_237) );
INVx4_ASAP7_75t_SL g151 ( .A(n_132), .Y(n_151) );
BUFx3_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_136), .A2(n_151), .B(n_166), .C(n_167), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g230 ( .A1(n_136), .A2(n_151), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_136), .A2(n_151), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_136), .A2(n_151), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_136), .A2(n_151), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_136), .A2(n_151), .B(n_540), .C(n_541), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_SL g575 ( .A1(n_136), .A2(n_151), .B(n_576), .C(n_577), .Y(n_575) );
INVx5_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx3_ASAP7_75t_L g149 ( .A(n_138), .Y(n_149) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_138), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_145), .C(n_148), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_142), .A2(n_148), .B(n_197), .C(n_198), .Y(n_196) );
O2A1O1Ixp5_ASAP7_75t_L g501 ( .A1(n_142), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_142), .A2(n_504), .B(n_533), .C(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_146), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g233 ( .A(n_146), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_146), .A2(n_210), .B(n_522), .C(n_523), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_146), .A2(n_169), .B1(n_579), .B2(n_580), .Y(n_578) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_147), .B(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g238 ( .A(n_149), .Y(n_238) );
INVx1_ASAP7_75t_L g493 ( .A(n_149), .Y(n_493) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_152), .A2(n_194), .B(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g212 ( .A(n_152), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_152), .Y(n_215) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_152), .A2(n_477), .B(n_484), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_152), .A2(n_246), .B(n_519), .C(n_520), .Y(n_518) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g163 ( .A(n_153), .B(n_154), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_L g435 ( .A(n_158), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
OR2x2_ASAP7_75t_L g298 ( .A(n_159), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_160), .B(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_160), .Y(n_291) );
INVx3_ASAP7_75t_L g306 ( .A(n_160), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_160), .B(n_176), .Y(n_330) );
OR2x2_ASAP7_75t_L g339 ( .A(n_160), .B(n_282), .Y(n_339) );
AND2x2_ASAP7_75t_L g343 ( .A(n_160), .B(n_303), .Y(n_343) );
AND2x2_ASAP7_75t_L g349 ( .A(n_160), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g386 ( .A(n_160), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_160), .B(n_243), .Y(n_400) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_164), .B(n_173), .Y(n_160) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_161), .A2(n_487), .B(n_494), .Y(n_486) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_161), .A2(n_509), .B(n_515), .Y(n_508) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_161), .A2(n_538), .B(n_545), .Y(n_537) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx4_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_162), .A2(n_179), .B(n_180), .Y(n_178) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g253 ( .A(n_163), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_168), .A2(n_221), .B(n_222), .C(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_169), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_169), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_172), .B(n_578), .Y(n_577) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_174), .A2(n_229), .B(n_239), .Y(n_228) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_175), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_175), .A2(n_218), .B(n_226), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_175), .B(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_175), .A2(n_244), .B(n_251), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_175), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_175), .B(n_525), .Y(n_524) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_175), .A2(n_529), .B(n_535), .Y(n_528) );
OR2x2_ASAP7_75t_L g292 ( .A(n_176), .B(n_243), .Y(n_292) );
AND2x2_ASAP7_75t_L g303 ( .A(n_176), .B(n_279), .Y(n_303) );
AND2x2_ASAP7_75t_L g315 ( .A(n_176), .B(n_306), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_176), .B(n_243), .Y(n_338) );
INVx1_ASAP7_75t_SL g350 ( .A(n_176), .Y(n_350) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g242 ( .A(n_177), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_177), .B(n_282), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_184), .B(n_185), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_185), .A2(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_201), .Y(n_190) );
AND2x2_ASAP7_75t_L g263 ( .A(n_191), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_191), .B(n_216), .Y(n_267) );
AND2x2_ASAP7_75t_L g270 ( .A(n_191), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_191), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g295 ( .A(n_191), .B(n_286), .Y(n_295) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_191), .Y(n_314) );
AND2x2_ASAP7_75t_L g335 ( .A(n_191), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g345 ( .A(n_191), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g391 ( .A(n_191), .B(n_274), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_191), .B(n_297), .Y(n_418) );
INVx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g288 ( .A(n_192), .Y(n_288) );
AND2x2_ASAP7_75t_L g354 ( .A(n_192), .B(n_286), .Y(n_354) );
AND2x2_ASAP7_75t_L g438 ( .A(n_192), .B(n_306), .Y(n_438) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_199), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_201), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_201), .Y(n_427) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_216), .Y(n_201) );
AND2x2_ASAP7_75t_L g257 ( .A(n_202), .B(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g266 ( .A(n_202), .B(n_264), .Y(n_266) );
INVx5_ASAP7_75t_L g274 ( .A(n_202), .Y(n_274) );
AND2x2_ASAP7_75t_L g297 ( .A(n_202), .B(n_228), .Y(n_297) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_202), .Y(n_334) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
AOI21xp5_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_206), .B(n_211), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_212), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_215), .A2(n_498), .B(n_505), .Y(n_497) );
INVx1_ASAP7_75t_L g375 ( .A(n_216), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_216), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g408 ( .A(n_216), .B(n_274), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_216), .A2(n_331), .B(n_438), .C(n_439), .Y(n_437) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_228), .Y(n_216) );
BUFx2_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
INVx2_ASAP7_75t_L g262 ( .A(n_217), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_225), .Y(n_218) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g544 ( .A(n_224), .Y(n_544) );
INVx2_ASAP7_75t_L g264 ( .A(n_228), .Y(n_264) );
AND2x2_ASAP7_75t_L g271 ( .A(n_228), .B(n_262), .Y(n_271) );
AND2x2_ASAP7_75t_L g362 ( .A(n_228), .B(n_274), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_236), .B(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g481 ( .A(n_237), .Y(n_481) );
INVx2_ASAP7_75t_L g504 ( .A(n_238), .Y(n_504) );
AOI211x1_ASAP7_75t_SL g240 ( .A1(n_241), .A2(n_255), .B(n_268), .C(n_293), .Y(n_240) );
INVx1_ASAP7_75t_L g359 ( .A(n_241), .Y(n_359) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_254), .Y(n_241) );
INVx5_ASAP7_75t_SL g279 ( .A(n_243), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_243), .B(n_349), .Y(n_348) );
AOI311xp33_ASAP7_75t_L g367 ( .A1(n_243), .A2(n_368), .A3(n_370), .B(n_371), .C(n_377), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g402 ( .A1(n_243), .A2(n_315), .B(n_403), .C(n_406), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_247), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_246), .A2(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_246), .A2(n_530), .B(n_531), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g572 ( .A(n_253), .Y(n_572) );
INVxp67_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
NAND4xp25_ASAP7_75t_SL g255 ( .A(n_256), .B(n_259), .C(n_265), .D(n_267), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_256), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g313 ( .A(n_257), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_260), .B(n_266), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_260), .B(n_273), .Y(n_393) );
BUFx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_261), .B(n_274), .Y(n_411) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g286 ( .A(n_262), .Y(n_286) );
INVxp67_ASAP7_75t_L g321 ( .A(n_263), .Y(n_321) );
AND2x4_ASAP7_75t_L g273 ( .A(n_264), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g347 ( .A(n_264), .B(n_286), .Y(n_347) );
INVx1_ASAP7_75t_L g374 ( .A(n_264), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_264), .B(n_361), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_265), .B(n_335), .Y(n_355) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_266), .B(n_288), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_266), .B(n_335), .Y(n_434) );
INVx1_ASAP7_75t_L g445 ( .A(n_267), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_275), .C(n_283), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g287 ( .A(n_271), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g325 ( .A(n_271), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g307 ( .A(n_272), .Y(n_307) );
AND2x2_ASAP7_75t_L g284 ( .A(n_273), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_273), .B(n_335), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_273), .B(n_354), .Y(n_378) );
OR2x2_ASAP7_75t_L g294 ( .A(n_274), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g326 ( .A(n_274), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_274), .B(n_286), .Y(n_341) );
AND2x2_ASAP7_75t_L g398 ( .A(n_274), .B(n_354), .Y(n_398) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_274), .Y(n_405) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_276), .A2(n_288), .B1(n_410), .B2(n_412), .C(n_415), .Y(n_409) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g299 ( .A(n_279), .B(n_282), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_279), .B(n_349), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_279), .B(n_306), .Y(n_414) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g399 ( .A(n_281), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g413 ( .A(n_281), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_282), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g310 ( .A(n_282), .B(n_303), .Y(n_310) );
AND2x2_ASAP7_75t_L g380 ( .A(n_282), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_282), .B(n_329), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_282), .B(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_287), .B(n_289), .Y(n_283) );
INVx2_ASAP7_75t_L g316 ( .A(n_284), .Y(n_316) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g336 ( .A(n_286), .Y(n_336) );
OR2x2_ASAP7_75t_L g340 ( .A(n_288), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g443 ( .A(n_288), .B(n_411), .Y(n_443) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AOI21xp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B(n_298), .Y(n_293) );
INVx1_ASAP7_75t_L g447 ( .A(n_294), .Y(n_447) );
INVx2_ASAP7_75t_SL g361 ( .A(n_295), .Y(n_361) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_298), .A2(n_379), .B(n_443), .C(n_444), .Y(n_442) );
OAI322xp33_ASAP7_75t_SL g311 ( .A1(n_299), .A2(n_312), .A3(n_315), .B1(n_316), .B2(n_317), .C1(n_319), .C2(n_322), .Y(n_311) );
INVx2_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B1(n_308), .B2(n_310), .C(n_311), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp33_ASAP7_75t_SL g377 ( .A1(n_302), .A2(n_378), .B1(n_379), .B2(n_382), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_303), .B(n_306), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_303), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g376 ( .A(n_305), .B(n_338), .Y(n_376) );
INVx1_ASAP7_75t_L g366 ( .A(n_306), .Y(n_366) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_310), .A2(n_420), .B(n_422), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g344 ( .A1(n_312), .A2(n_345), .B(n_348), .Y(n_344) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp67_ASAP7_75t_SL g373 ( .A(n_314), .B(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_314), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g430 ( .A(n_315), .Y(n_430) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND4xp25_ASAP7_75t_L g323 ( .A(n_324), .B(n_351), .C(n_367), .D(n_383), .Y(n_323) );
AOI211xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B(n_332), .C(n_344), .Y(n_324) );
INVx1_ASAP7_75t_L g416 ( .A(n_325), .Y(n_416) );
AND2x2_ASAP7_75t_L g364 ( .A(n_326), .B(n_347), .Y(n_364) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_331), .B(n_366), .Y(n_365) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_337), .B1(n_340), .B2(n_342), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_334), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g382 ( .A(n_335), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g396 ( .A1(n_335), .A2(n_374), .B(n_397), .C(n_399), .Y(n_396) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g381 ( .A(n_338), .Y(n_381) );
INVx1_ASAP7_75t_L g441 ( .A(n_339), .Y(n_441) );
NAND2xp33_ASAP7_75t_SL g431 ( .A(n_340), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g370 ( .A(n_349), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B(n_356), .C(n_358), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_363), .B2(n_365), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_361), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_366), .B(n_387), .Y(n_449) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI21xp33_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_375), .B(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_389), .B1(n_392), .B2(n_394), .C(n_396), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_399), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g401 ( .A(n_402), .B(n_409), .C(n_419), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B(n_428), .C(n_437), .Y(n_425) );
INVx1_ASAP7_75t_L g446 ( .A(n_426), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_433), .B2(n_435), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_447), .B2(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g462 ( .A(n_454), .Y(n_462) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_459), .B(n_464), .C(n_749), .Y(n_463) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g748 ( .A(n_471), .Y(n_748) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_668), .Y(n_471) );
NAND5xp2_ASAP7_75t_L g472 ( .A(n_473), .B(n_583), .C(n_615), .D(n_632), .E(n_655), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_516), .B1(n_546), .B2(n_550), .C(n_554), .Y(n_473) );
INVx1_ASAP7_75t_L g695 ( .A(n_474), .Y(n_695) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_495), .Y(n_474) );
AND3x2_ASAP7_75t_L g670 ( .A(n_475), .B(n_497), .C(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_476), .B(n_552), .Y(n_551) );
BUFx3_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
AND2x2_ASAP7_75t_L g565 ( .A(n_476), .B(n_507), .Y(n_565) );
INVx2_ASAP7_75t_L g592 ( .A(n_476), .Y(n_592) );
OR2x2_ASAP7_75t_L g603 ( .A(n_476), .B(n_508), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_476), .B(n_496), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_476), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g682 ( .A(n_476), .B(n_508), .Y(n_682) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
AND2x2_ASAP7_75t_L g623 ( .A(n_485), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_485), .B(n_496), .Y(n_642) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g553 ( .A(n_486), .B(n_496), .Y(n_553) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_486), .Y(n_560) );
AND2x2_ASAP7_75t_L g609 ( .A(n_486), .B(n_508), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_486), .B(n_495), .C(n_592), .Y(n_634) );
AND2x2_ASAP7_75t_L g699 ( .A(n_486), .B(n_497), .Y(n_699) );
AND2x2_ASAP7_75t_L g733 ( .A(n_486), .B(n_496), .Y(n_733) );
INVxp67_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_507), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_496), .B(n_592), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_496), .B(n_623), .Y(n_631) );
AND2x2_ASAP7_75t_L g681 ( .A(n_496), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g709 ( .A(n_496), .Y(n_709) );
INVx4_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g616 ( .A(n_497), .B(n_609), .Y(n_616) );
BUFx3_ASAP7_75t_L g648 ( .A(n_497), .Y(n_648) );
INVx2_ASAP7_75t_L g624 ( .A(n_507), .Y(n_624) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_516), .A2(n_684), .B1(n_686), .B2(n_687), .Y(n_683) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
AND2x2_ASAP7_75t_L g546 ( .A(n_517), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_SL g557 ( .A(n_517), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_517), .B(n_587), .Y(n_619) );
OR2x2_ASAP7_75t_L g638 ( .A(n_517), .B(n_527), .Y(n_638) );
AND2x2_ASAP7_75t_L g643 ( .A(n_517), .B(n_595), .Y(n_643) );
AND2x2_ASAP7_75t_L g646 ( .A(n_517), .B(n_588), .Y(n_646) );
AND2x2_ASAP7_75t_L g658 ( .A(n_517), .B(n_537), .Y(n_658) );
AND2x2_ASAP7_75t_L g674 ( .A(n_517), .B(n_528), .Y(n_674) );
AND2x4_ASAP7_75t_L g677 ( .A(n_517), .B(n_548), .Y(n_677) );
OR2x2_ASAP7_75t_L g694 ( .A(n_517), .B(n_630), .Y(n_694) );
OR2x2_ASAP7_75t_L g725 ( .A(n_517), .B(n_570), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_517), .B(n_653), .Y(n_727) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
AND2x2_ASAP7_75t_L g601 ( .A(n_526), .B(n_568), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_526), .B(n_588), .Y(n_720) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
AND2x2_ASAP7_75t_L g556 ( .A(n_527), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g587 ( .A(n_527), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g595 ( .A(n_527), .B(n_570), .Y(n_595) );
AND2x2_ASAP7_75t_L g613 ( .A(n_527), .B(n_548), .Y(n_613) );
OR2x2_ASAP7_75t_L g630 ( .A(n_527), .B(n_588), .Y(n_630) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g549 ( .A(n_528), .Y(n_549) );
AND2x2_ASAP7_75t_L g653 ( .A(n_528), .B(n_537), .Y(n_653) );
INVx2_ASAP7_75t_L g548 ( .A(n_537), .Y(n_548) );
INVx1_ASAP7_75t_L g665 ( .A(n_537), .Y(n_665) );
AND2x2_ASAP7_75t_L g715 ( .A(n_537), .B(n_557), .Y(n_715) );
AND2x2_ASAP7_75t_L g567 ( .A(n_547), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g599 ( .A(n_547), .B(n_557), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_547), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x2_ASAP7_75t_L g586 ( .A(n_548), .B(n_557), .Y(n_586) );
OR2x2_ASAP7_75t_L g702 ( .A(n_549), .B(n_676), .Y(n_702) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_552), .B(n_682), .Y(n_688) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OAI32xp33_ASAP7_75t_L g644 ( .A1(n_553), .A2(n_645), .A3(n_647), .B1(n_649), .B2(n_650), .Y(n_644) );
OR2x2_ASAP7_75t_L g661 ( .A(n_553), .B(n_603), .Y(n_661) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_553), .A2(n_563), .B(n_591), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B1(n_563), .B2(n_566), .Y(n_554) );
INVxp33_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_556), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_557), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g612 ( .A(n_557), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g712 ( .A(n_557), .B(n_653), .Y(n_712) );
OR2x2_ASAP7_75t_L g736 ( .A(n_557), .B(n_630), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_558), .A2(n_618), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_560), .B(n_565), .Y(n_614) );
AND2x2_ASAP7_75t_L g636 ( .A(n_561), .B(n_609), .Y(n_636) );
INVx1_ASAP7_75t_L g649 ( .A(n_561), .Y(n_649) );
OR2x2_ASAP7_75t_L g654 ( .A(n_561), .B(n_588), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_564), .B(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_565), .A2(n_585), .B1(n_590), .B2(n_594), .Y(n_584) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_568), .A2(n_627), .B1(n_634), .B2(n_635), .Y(n_633) );
AND2x2_ASAP7_75t_L g711 ( .A(n_568), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_570), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g730 ( .A(n_570), .B(n_613), .Y(n_730) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B(n_581), .Y(n_570) );
INVx1_ASAP7_75t_L g589 ( .A(n_571), .Y(n_589) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OA21x2_ASAP7_75t_L g588 ( .A1(n_574), .A2(n_582), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_596), .B1(n_597), .B2(n_602), .C(n_604), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_586), .B(n_588), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_586), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g605 ( .A(n_587), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_587), .A2(n_693), .B(n_694), .C(n_695), .Y(n_692) );
AND2x2_ASAP7_75t_L g697 ( .A(n_587), .B(n_677), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_SL g735 ( .A1(n_587), .A2(n_676), .B(n_736), .C(n_737), .Y(n_735) );
BUFx3_ASAP7_75t_L g627 ( .A(n_588), .Y(n_627) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_591), .B(n_648), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g710 ( .A1(n_591), .A2(n_711), .B(n_713), .C(n_719), .Y(n_710) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVxp67_ASAP7_75t_L g671 ( .A(n_593), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_595), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_599), .A2(n_616), .B(n_617), .C(n_625), .Y(n_615) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g700 ( .A(n_603), .Y(n_700) );
OR2x2_ASAP7_75t_L g717 ( .A(n_603), .B(n_647), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_611), .B2(n_614), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_606), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
OR2x2_ASAP7_75t_L g704 ( .A(n_608), .B(n_648), .Y(n_704) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g659 ( .A(n_609), .B(n_649), .Y(n_659) );
INVx1_ASAP7_75t_L g667 ( .A(n_610), .Y(n_667) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_613), .B(n_627), .Y(n_675) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_623), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g732 ( .A(n_624), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_631), .Y(n_625) );
INVx1_ASAP7_75t_L g662 ( .A(n_626), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_627), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_627), .B(n_658), .Y(n_657) );
NAND2x1p5_ASAP7_75t_L g678 ( .A(n_627), .B(n_653), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_627), .B(n_674), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_627), .A2(n_637), .B(n_677), .C(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_637), .B1(n_639), .B2(n_643), .C(n_644), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_641), .B(n_649), .Y(n_723) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_643), .A2(n_658), .B(n_660), .C(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_646), .B(n_653), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_647), .B(n_700), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g647 ( .A(n_648), .Y(n_647) );
INVxp33_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
AOI21xp33_ASAP7_75t_SL g663 ( .A1(n_652), .A2(n_664), .B(n_666), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_652), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_653), .B(n_707), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_660), .B2(n_662), .C(n_663), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_659), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g693 ( .A(n_665), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g668 ( .A(n_669), .B(n_696), .C(n_710), .D(n_721), .E(n_734), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B(n_679), .C(n_692), .Y(n_669) );
INVx2_ASAP7_75t_SL g716 ( .A(n_670), .Y(n_716) );
NAND4xp25_ASAP7_75t_SL g672 ( .A(n_673), .B(n_675), .C(n_676), .D(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_678), .A2(n_680), .B(n_683), .C(n_689), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_681), .A2(n_722), .B1(n_724), .B2(n_726), .C(n_728), .Y(n_721) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_698), .B1(n_701), .B2(n_703), .C(n_705), .Y(n_696) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_704), .A2(n_727), .B1(n_729), .B2(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
endmodule