module fake_jpeg_16957_n_28 (n_3, n_2, n_1, n_0, n_4, n_5, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

AND2x2_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_5),
.Y(n_6)
);

INVx5_ASAP7_75t_SL g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_6),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx12_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_16),
.B(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

NAND2x1p5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_7),
.Y(n_23)
);

OA21x2_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_20),
.B(n_6),
.Y(n_21)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_12),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_11),
.B2(n_0),
.Y(n_28)
);

AOI322xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_23),
.A3(n_22),
.B1(n_19),
.B2(n_7),
.C1(n_11),
.C2(n_10),
.Y(n_27)
);


endmodule