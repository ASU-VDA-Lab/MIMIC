module fake_jpeg_15300_n_375 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_38),
.B(n_50),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_41),
.B(n_43),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_44),
.B(n_59),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_53),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_32),
.B(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_56),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_32),
.B(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_23),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_37),
.B1(n_24),
.B2(n_19),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_76),
.B1(n_78),
.B2(n_86),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_15),
.B1(n_25),
.B2(n_24),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_72),
.A2(n_79),
.B1(n_118),
.B2(n_4),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_37),
.B1(n_24),
.B2(n_19),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_25),
.B1(n_15),
.B2(n_37),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_77),
.A2(n_88),
.B1(n_115),
.B2(n_53),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_25),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_42),
.B(n_25),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_102),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_31),
.B1(n_20),
.B2(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_38),
.A2(n_36),
.B1(n_30),
.B2(n_22),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_31),
.B1(n_30),
.B2(n_22),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_90),
.A2(n_101),
.B1(n_108),
.B2(n_4),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_20),
.C(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_96),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_14),
.B(n_34),
.C(n_29),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_14),
.B1(n_29),
.B2(n_6),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_105),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_61),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_47),
.A2(n_29),
.B1(n_5),
.B2(n_6),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_45),
.B(n_18),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_119),
.Y(n_154)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_18),
.B1(n_33),
.B2(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_33),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_116),
.B(n_11),
.Y(n_159)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_49),
.A2(n_33),
.B1(n_23),
.B2(n_7),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_123),
.Y(n_183)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_33),
.B1(n_23),
.B2(n_7),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_124),
.A2(n_157),
.B1(n_121),
.B2(n_170),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_125),
.B(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_23),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_126),
.B(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_4),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_139),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_80),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_133),
.Y(n_184)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_149),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_136),
.A2(n_122),
.B(n_152),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_138),
.A2(n_155),
.B1(n_164),
.B2(n_166),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_4),
.Y(n_139)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_71),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_73),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_151),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_70),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_157),
.B1(n_167),
.B2(n_84),
.Y(n_177)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_107),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_70),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_113),
.B(n_10),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_11),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_98),
.A2(n_97),
.B1(n_119),
.B2(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_98),
.A2(n_12),
.B1(n_111),
.B2(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_116),
.A2(n_12),
.B1(n_85),
.B2(n_94),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_137),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_96),
.B(n_12),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_81),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_73),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_171),
.A2(n_207),
.B(n_215),
.Y(n_244)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_176),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_178),
.B1(n_196),
.B2(n_198),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_74),
.B1(n_82),
.B2(n_99),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_182),
.B(n_151),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_193),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_103),
.C(n_114),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_140),
.C(n_145),
.Y(n_224)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_129),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_183),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_138),
.A2(n_131),
.B1(n_147),
.B2(n_167),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_199),
.A2(n_205),
.B1(n_191),
.B2(n_195),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_143),
.A2(n_144),
.B1(n_170),
.B2(n_153),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_206),
.B1(n_213),
.B2(n_187),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_147),
.A2(n_131),
.B1(n_127),
.B2(n_132),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_204),
.A2(n_191),
.B1(n_196),
.B2(n_207),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_125),
.A2(n_134),
.B1(n_161),
.B2(n_149),
.Y(n_205)
);

INVx4_ASAP7_75t_SL g206 ( 
.A(n_162),
.Y(n_206)
);

OR2x2_ASAP7_75t_SL g207 ( 
.A(n_169),
.B(n_159),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_143),
.A2(n_144),
.B1(n_135),
.B2(n_163),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_150),
.A2(n_120),
.B(n_130),
.Y(n_215)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_230),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_146),
.B(n_133),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_214),
.B(n_193),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_137),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_223),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_206),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_140),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_227),
.C(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_225),
.B(n_228),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_174),
.B(n_205),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_171),
.B(n_179),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_242),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_237),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_251),
.B1(n_211),
.B2(n_194),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_177),
.B(n_178),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_180),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_190),
.A2(n_188),
.B(n_209),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_248),
.B(n_200),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_181),
.Y(n_247)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_198),
.A2(n_206),
.B1(n_176),
.B2(n_185),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_185),
.C(n_201),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_214),
.B1(n_187),
.B2(n_180),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_186),
.B(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_257),
.A2(n_259),
.B(n_220),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_272),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_211),
.B(n_172),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_262),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_309)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_175),
.A3(n_194),
.B1(n_200),
.B2(n_223),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_264),
.B(n_259),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_265),
.A2(n_270),
.B(n_255),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_273),
.C(n_277),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_224),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_220),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_239),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_236),
.B1(n_218),
.B2(n_219),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_234),
.B1(n_249),
.B2(n_247),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_245),
.B1(n_253),
.B2(n_226),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_217),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_225),
.A2(n_226),
.B1(n_232),
.B2(n_251),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_238),
.A2(n_240),
.B1(n_254),
.B2(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_288),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_221),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_289),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_220),
.C(n_246),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_298),
.Y(n_326)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_294),
.B(n_306),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_257),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_308),
.C(n_312),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_299),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_280),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_283),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_304),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_270),
.A2(n_281),
.B1(n_276),
.B2(n_275),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_307),
.B1(n_311),
.B2(n_269),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_286),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_263),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_310),
.B1(n_269),
.B2(n_271),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_256),
.B(n_278),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_266),
.Y(n_308)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_277),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_325),
.B1(n_323),
.B2(n_331),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_258),
.C(n_265),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_332),
.C(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_309),
.B1(n_305),
.B2(n_294),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_323),
.B1(n_331),
.B2(n_313),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_309),
.A2(n_264),
.B1(n_271),
.B2(n_300),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_328),
.A2(n_330),
.B1(n_295),
.B2(n_290),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_301),
.B1(n_298),
.B2(n_296),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_312),
.C(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_333),
.B(n_338),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_291),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_335),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_310),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_336),
.B(n_317),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_293),
.C(n_288),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_344),
.C(n_345),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_318),
.A2(n_299),
.B(n_307),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_339),
.A2(n_340),
.B1(n_342),
.B2(n_347),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_315),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_326),
.A2(n_311),
.B1(n_325),
.B2(n_328),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_321),
.C(n_320),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_330),
.C(n_327),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_317),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_346),
.B(n_338),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_324),
.A2(n_314),
.B1(n_326),
.B2(n_329),
.Y(n_347)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_343),
.A2(n_347),
.B1(n_345),
.B2(n_340),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_356),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_319),
.C(n_329),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_353),
.C(n_354),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_342),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_339),
.C(n_343),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_334),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_355),
.A2(n_334),
.B1(n_353),
.B2(n_358),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_354),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_362),
.A2(n_358),
.B(n_357),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_355),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_365),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_367),
.C(n_368),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_349),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_359),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g372 ( 
.A1(n_371),
.A2(n_369),
.B(n_363),
.C(n_360),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_372),
.A2(n_363),
.B(n_349),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_367),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_374),
.Y(n_375)
);


endmodule