module fake_jpeg_25817_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_27),
.Y(n_52)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_44),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_79),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

OR2x4_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_40),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_22),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_72),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_78),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_81),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_87),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_37),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_47),
.B1(n_38),
.B2(n_42),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_54),
.B1(n_47),
.B2(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_92),
.Y(n_121)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_96),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_63),
.C(n_40),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_104),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_47),
.B1(n_46),
.B2(n_38),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_111),
.B1(n_120),
.B2(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_39),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_40),
.C(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_115),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_89),
.B1(n_73),
.B2(n_78),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_47),
.B1(n_42),
.B2(n_45),
.Y(n_111)
);

AO22x2_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_62),
.B1(n_64),
.B2(n_41),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_89),
.B1(n_73),
.B2(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_84),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_45),
.B1(n_41),
.B2(n_29),
.Y(n_120)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_130),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_31),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_152),
.B1(n_122),
.B2(n_17),
.Y(n_185)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_144),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_24),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_94),
.B1(n_45),
.B2(n_95),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_112),
.B1(n_117),
.B2(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_8),
.Y(n_145)
);

XOR2x2_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_29),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_30),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_25),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_111),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_95),
.B1(n_30),
.B2(n_36),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_25),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_154),
.A2(n_155),
.B(n_101),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_161),
.B1(n_171),
.B2(n_186),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_117),
.B(n_125),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_160),
.A2(n_164),
.B(n_169),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_113),
.B1(n_116),
.B2(n_100),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_149),
.B(n_148),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_113),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_184),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_101),
.B(n_115),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_170),
.B(n_175),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_100),
.B1(n_107),
.B2(n_108),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_109),
.B(n_108),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_173),
.B(n_176),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_118),
.C(n_125),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_140),
.C(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_135),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_123),
.B(n_76),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_181),
.B(n_22),
.Y(n_218)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_122),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_146),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_137),
.B1(n_129),
.B2(n_134),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_195),
.B1(n_197),
.B2(n_210),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_184),
.C(n_160),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_194),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_192),
.B(n_196),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_145),
.B1(n_130),
.B2(n_139),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_130),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_141),
.B1(n_138),
.B2(n_76),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_156),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_199),
.B(n_201),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_168),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_138),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_202),
.B(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_208),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_157),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_157),
.B1(n_167),
.B2(n_163),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_35),
.B1(n_31),
.B2(n_32),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_33),
.B1(n_28),
.B2(n_23),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_34),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_11),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_215),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_10),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_170),
.C(n_166),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_169),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_204),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_208),
.B1(n_206),
.B2(n_209),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_198),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_229),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_172),
.C(n_177),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_237),
.C(n_239),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_173),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_203),
.Y(n_262)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_181),
.C(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_201),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_186),
.C(n_159),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_158),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_182),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_217),
.C(n_191),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_193),
.C(n_212),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_220),
.B1(n_231),
.B2(n_232),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_254),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_205),
.B(n_226),
.C(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_188),
.B1(n_193),
.B2(n_195),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_252),
.A2(n_261),
.B1(n_23),
.B2(n_21),
.Y(n_284)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_257),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_191),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_215),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_234),
.B1(n_224),
.B2(n_220),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_266),
.B1(n_238),
.B2(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_241),
.B1(n_157),
.B2(n_163),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_210),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_243),
.C(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_230),
.CI(n_239),
.CON(n_268),
.SN(n_268)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_270),
.B(n_274),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_232),
.B1(n_214),
.B2(n_223),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_271),
.A2(n_273),
.B1(n_275),
.B2(n_21),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_241),
.B1(n_211),
.B2(n_180),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_249),
.B1(n_253),
.B2(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_263),
.C(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_281),
.C(n_283),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_252),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_221),
.C(n_162),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_34),
.C(n_28),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_20),
.B1(n_8),
.B2(n_9),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_280),
.B(n_265),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_285),
.B(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_291),
.B1(n_10),
.B2(n_16),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_291)
);

AOI21x1_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_0),
.B(n_3),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_291),
.B(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_8),
.C(n_15),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_283),
.C(n_278),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_7),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_272),
.B(n_282),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_299),
.B(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_270),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_301),
.B(n_305),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_296),
.B(n_292),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_290),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_278),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_0),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_268),
.B1(n_3),
.B2(n_4),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_312)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_287),
.B(n_294),
.C(n_286),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_312),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_320),
.A2(n_307),
.B1(n_303),
.B2(n_305),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_324),
.A3(n_321),
.B1(n_317),
.B2(n_326),
.C1(n_325),
.C2(n_316),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_301),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_328),
.B(n_12),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_309),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_9),
.C(n_15),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_331),
.A3(n_332),
.B1(n_15),
.B2(n_16),
.C1(n_5),
.C2(n_6),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_16),
.C(n_4),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_0),
.Y(n_337)
);

AOI221xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_5),
.B1(n_6),
.B2(n_229),
.C(n_203),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_5),
.Y(n_339)
);


endmodule