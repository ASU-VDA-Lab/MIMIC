module fake_jpeg_27021_n_412 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_412);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_412;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_6),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_20),
.A2(n_6),
.B(n_3),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_87),
.B(n_29),
.Y(n_128)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_6),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_64),
.A2(n_29),
.B1(n_41),
.B2(n_30),
.Y(n_135)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx8_ASAP7_75t_SL g71 ( 
.A(n_19),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_71),
.Y(n_98)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_19),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_13),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_28),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_77),
.Y(n_136)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_3),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_24),
.Y(n_80)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_36),
.Y(n_84)
);

CKINVDCx9p33_ASAP7_75t_R g125 ( 
.A(n_84),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_22),
.B(n_3),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_134),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_46),
.B1(n_34),
.B2(n_44),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_100),
.A2(n_85),
.B1(n_84),
.B2(n_77),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_46),
.B1(n_34),
.B2(n_38),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_115),
.B1(n_86),
.B2(n_81),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_54),
.A2(n_46),
.B1(n_34),
.B2(n_38),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_59),
.B1(n_51),
.B2(n_78),
.Y(n_165)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_22),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_47),
.Y(n_137)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_50),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_139),
.A2(n_164),
.B1(n_173),
.B2(n_115),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_41),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_140),
.B(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_145),
.Y(n_193)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

CKINVDCx12_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_148),
.Y(n_208)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_30),
.Y(n_153)
);

CKINVDCx6p67_ASAP7_75t_R g154 ( 
.A(n_90),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_157),
.Y(n_210)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_45),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_SL g216 ( 
.A(n_165),
.B(n_44),
.C(n_27),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_96),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_167),
.Y(n_192)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_95),
.B(n_43),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_43),
.Y(n_171)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_119),
.B(n_32),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_98),
.B(n_32),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_39),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_39),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_136),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_94),
.B1(n_124),
.B2(n_114),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_91),
.B1(n_109),
.B2(n_126),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_149),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_133),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_180),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_216),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_205),
.B1(n_160),
.B2(n_172),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_139),
.A2(n_130),
.B1(n_124),
.B2(n_114),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_49),
.C(n_123),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_170),
.C(n_168),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_72),
.A3(n_82),
.B1(n_69),
.B2(n_129),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_31),
.B(n_42),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_219),
.A2(n_215),
.B1(n_217),
.B2(n_198),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_175),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_221),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_229),
.Y(n_260)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_156),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_242),
.Y(n_270)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_233),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_149),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_231),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_26),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_197),
.B(n_45),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_235),
.A2(n_236),
.B1(n_241),
.B2(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_215),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_198),
.B1(n_217),
.B2(n_144),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_184),
.B(n_195),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_238),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_101),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_244),
.B(n_42),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_154),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_101),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_117),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_186),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_249),
.B1(n_150),
.B2(n_204),
.Y(n_276)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_192),
.C(n_188),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_252),
.C(n_259),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_189),
.C(n_154),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_185),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_258),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_185),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_189),
.C(n_187),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_196),
.B(n_31),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_271),
.B(n_273),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_187),
.C(n_208),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_26),
.B(n_25),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_237),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_239),
.A2(n_25),
.B(n_0),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_222),
.A2(n_0),
.B(n_4),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_0),
.B(n_222),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

AO22x1_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_94),
.B1(n_204),
.B2(n_117),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_279),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_234),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_281),
.B(n_282),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_294),
.Y(n_309)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_285),
.Y(n_325)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_286),
.B(n_296),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_269),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_291),
.Y(n_317)
);

AO22x1_ASAP7_75t_L g294 ( 
.A1(n_266),
.A2(n_228),
.B1(n_224),
.B2(n_245),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_303),
.B1(n_274),
.B2(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_297),
.B(n_299),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_255),
.B(n_249),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_301),
.B(n_302),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_243),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_270),
.C(n_254),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_314),
.C(n_322),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_259),
.Y(n_306)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_270),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_311),
.B(n_318),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_313),
.B1(n_280),
.B2(n_298),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_287),
.A2(n_265),
.B1(n_251),
.B2(n_263),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_254),
.C(n_275),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_271),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_284),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_321),
.B(n_327),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_256),
.C(n_227),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_227),
.B1(n_206),
.B2(n_147),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_326),
.A2(n_132),
.B1(n_118),
.B2(n_103),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_298),
.C(n_302),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_342),
.C(n_343),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_335),
.A2(n_338),
.B1(n_344),
.B2(n_345),
.Y(n_361)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

O2A1O1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_294),
.B(n_295),
.C(n_288),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_307),
.A2(n_280),
.B1(n_283),
.B2(n_293),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_317),
.B(n_290),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_341),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_290),
.C(n_206),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_158),
.C(n_162),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_300),
.B1(n_286),
.B2(n_158),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_313),
.Y(n_347)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g348 ( 
.A(n_331),
.B(n_322),
.CI(n_318),
.CON(n_348),
.SN(n_348)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_324),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_351),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_316),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_335),
.B(n_306),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_355),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_310),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_308),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_362),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_326),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_359),
.A2(n_332),
.B(n_310),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_364),
.A2(n_338),
.B(n_323),
.Y(n_376)
);

AO221x1_ASAP7_75t_L g368 ( 
.A1(n_357),
.A2(n_328),
.B1(n_319),
.B2(n_353),
.C(n_356),
.Y(n_368)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_361),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_371),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_344),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_375),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_342),
.C(n_352),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_374),
.C(n_350),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_329),
.C(n_334),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_323),
.Y(n_375)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_351),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_385),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_384),
.C(n_367),
.Y(n_390)
);

NOR2x1_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_348),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_386),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_370),
.B(n_345),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_381),
.B(n_363),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_161),
.C(n_146),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_151),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_365),
.A2(n_4),
.B(n_5),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_390),
.B(n_391),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_363),
.C(n_367),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_392),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_377),
.C(n_382),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_394),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_383),
.A2(n_371),
.B1(n_118),
.B2(n_83),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_151),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_395),
.A2(n_8),
.B1(n_12),
.B2(n_163),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_389),
.A2(n_386),
.B1(n_44),
.B2(n_12),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_400),
.Y(n_404)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_399),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_120),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_396),
.A2(n_395),
.B(n_387),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_387),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_405),
.A2(n_406),
.B(n_401),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_397),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_403),
.B(n_398),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_409),
.B(n_8),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_410),
.A2(n_12),
.B1(n_163),
.B2(n_120),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_411),
.A2(n_52),
.B(n_58),
.Y(n_412)
);


endmodule