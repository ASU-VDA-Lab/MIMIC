module fake_jpeg_30457_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_74),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_65),
.B1(n_57),
.B2(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_65),
.B1(n_57),
.B2(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_52),
.B1(n_53),
.B2(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_3),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_47),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_63),
.B1(n_62),
.B2(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_52),
.B1(n_55),
.B2(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_46),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_100),
.Y(n_119)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_80),
.B1(n_79),
.B2(n_47),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_2),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_104),
.Y(n_122)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_4),
.Y(n_127)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_90),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_23),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_97),
.B(n_105),
.C(n_95),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_116),
.B(n_118),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_8),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_127),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_25),
.B(n_40),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_30),
.B(n_37),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_9),
.B(n_10),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_128),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_27),
.C(n_38),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_133),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_147),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_5),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_136),
.B1(n_144),
.B2(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_6),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_29),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_7),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_143),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_114),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_31),
.B(n_36),
.C(n_13),
.D(n_15),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_113),
.C(n_111),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_130),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_122),
.B1(n_112),
.B2(n_9),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_145),
.B1(n_112),
.B2(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_160),
.B(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.C(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_148),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_153),
.B(n_158),
.C(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_148),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_138),
.B(n_147),
.C(n_21),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_35),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_32),
.Y(n_169)
);


endmodule