module fake_netlist_5_1008_n_2264 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2264);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2264;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_1070;
wire n_777;
wire n_422;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_2248;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_378;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2213;
wire n_2023;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_333;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2044;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_92),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_51),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_159),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_107),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_126),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_43),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_96),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_14),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_133),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_36),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_46),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_71),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_7),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_180),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_36),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_108),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_192),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_81),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_109),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_121),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_193),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_8),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_44),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_149),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_83),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_30),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_89),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_84),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_79),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_26),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_29),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_125),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_115),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_87),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_65),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_34),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_87),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_50),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_24),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_191),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_200),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_63),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_37),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_81),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_24),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_58),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_44),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_88),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_60),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_197),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_143),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_73),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_113),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_132),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_123),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_111),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_63),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_2),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_37),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_33),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_183),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_182),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_129),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_66),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_169),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_154),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_57),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_9),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_38),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_82),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_127),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_194),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_20),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_46),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_157),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_16),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_148),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_8),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_118),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_179),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_211),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_54),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_10),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_153),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_112),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_12),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_33),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_68),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_124),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_79),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_208),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_53),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_136),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_146),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_59),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_22),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_122),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_32),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_84),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_61),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_77),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_145),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_3),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_103),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_162),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_90),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_88),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_2),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_53),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_152),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_85),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_173),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_77),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_39),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_195),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_76),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_218),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_172),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_30),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_86),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_174),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_45),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_207),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_32),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_1),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_54),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_160),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_93),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_75),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_85),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_47),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_167),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_42),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_120),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_73),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_204),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_117),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_100),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_35),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_101),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_35),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_138),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_40),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_116),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_39),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_91),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_128),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_50),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_3),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_49),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_65),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_34),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_92),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_49),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_99),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_205),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_213),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_110),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_177),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_0),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_57),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_18),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_98),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_7),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_47),
.Y(n_401)
);

BUFx5_ASAP7_75t_L g402 ( 
.A(n_21),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_6),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_38),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_82),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_58),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_6),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_102),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_93),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_41),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_22),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_106),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_42),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_186),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_59),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_13),
.Y(n_416)
);

BUFx2_ASAP7_75t_SL g417 ( 
.A(n_1),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_184),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_105),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_141),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_151),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_0),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_48),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_13),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_217),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_168),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_165),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_27),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_104),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_163),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_70),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_265),
.B(n_4),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_4),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_291),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_291),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_308),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_221),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_308),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_325),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_308),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_224),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_308),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_308),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_222),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_308),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_263),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_308),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_308),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_308),
.B(n_5),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_325),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_275),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_225),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_402),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_230),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_227),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_260),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_266),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_271),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_229),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_367),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_231),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_236),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_240),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_402),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_245),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_252),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_402),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_275),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_420),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_223),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_269),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_234),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_297),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_254),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_306),
.B(n_5),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_267),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_254),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_265),
.B(n_9),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_254),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_284),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_254),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_370),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_254),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_329),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_270),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_285),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_294),
.B(n_11),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_276),
.Y(n_494)
);

INVxp33_ASAP7_75t_SL g495 ( 
.A(n_219),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_276),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_306),
.B(n_11),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_276),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_297),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_287),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_288),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_289),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_312),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_315),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_319),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_324),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_326),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_276),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_328),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_332),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_347),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_307),
.B(n_12),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_294),
.B(n_14),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_276),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_307),
.B(n_15),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_228),
.B(n_15),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_220),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_337),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_282),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_339),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_345),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_362),
.B(n_17),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_357),
.B(n_17),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_350),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_232),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_353),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_282),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_369),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_371),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_282),
.Y(n_530)
);

BUFx6f_ASAP7_75t_SL g531 ( 
.A(n_347),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_372),
.Y(n_532)
);

INVxp33_ASAP7_75t_SL g533 ( 
.A(n_247),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_282),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_375),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_282),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_397),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_397),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_377),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_379),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_382),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_405),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_405),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_233),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_233),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_478),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_523),
.B(n_357),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_480),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_480),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_461),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_523),
.B(n_383),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_471),
.B(n_391),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_479),
.B(n_393),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_483),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_444),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_437),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_499),
.B(n_383),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_475),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_485),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_452),
.B(n_384),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_452),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g563 ( 
.A(n_446),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_497),
.B(n_250),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_475),
.B(n_362),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_446),
.B(n_347),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_451),
.B(n_223),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_441),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_475),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_457),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_459),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_487),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_511),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_451),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_453),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_R g579 ( 
.A(n_490),
.B(n_394),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_452),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_456),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_489),
.Y(n_582)
);

BUFx8_ASAP7_75t_L g583 ( 
.A(n_531),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_489),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_494),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_494),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_496),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_460),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_496),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_436),
.B(n_395),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_498),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_463),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_451),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_498),
.B(n_384),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_464),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_436),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_465),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_467),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_469),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_495),
.B(n_347),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_508),
.B(n_228),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_476),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_486),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_525),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_497),
.B(n_512),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_492),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_502),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_505),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_438),
.Y(n_611)
);

BUFx8_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_519),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_R g616 ( 
.A(n_507),
.B(n_399),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_519),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_R g618 ( 
.A(n_500),
.B(n_412),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_527),
.B(n_408),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_438),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_440),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_530),
.B(n_408),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_530),
.B(n_238),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_509),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_534),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_518),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_534),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_481),
.B(n_414),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_520),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_440),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_488),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_442),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_434),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_536),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_607),
.B(n_511),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_607),
.B(n_533),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_611),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_569),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_553),
.B(n_521),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_550),
.B(n_524),
.Y(n_641)
);

NAND3x1_ASAP7_75t_L g642 ( 
.A(n_629),
.B(n_433),
.C(n_512),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_611),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_611),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_553),
.B(n_528),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_577),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_550),
.B(n_576),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_577),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_580),
.B(n_529),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_561),
.B(n_511),
.Y(n_650)
);

INVx6_ASAP7_75t_L g651 ( 
.A(n_559),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_620),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_620),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_562),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_559),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_557),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_546),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_620),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_559),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_580),
.B(n_238),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_634),
.B(n_455),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_570),
.Y(n_662)
);

BUFx4f_ASAP7_75t_L g663 ( 
.A(n_569),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_559),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_550),
.B(n_532),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_562),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_601),
.B(n_223),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_562),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_621),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_577),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_634),
.B(n_455),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_569),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_593),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_559),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_561),
.B(n_537),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_621),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_621),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_580),
.B(n_239),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_593),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_601),
.B(n_239),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_569),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_554),
.B(n_535),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_615),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_567),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_631),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_561),
.B(n_537),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_569),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_554),
.B(n_540),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_629),
.B(n_541),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_631),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_558),
.B(n_538),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_578),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_558),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_546),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_596),
.B(n_536),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_632),
.B(n_435),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_593),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_615),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_631),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_601),
.B(n_242),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_558),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_547),
.A2(n_515),
.B1(n_516),
.B2(n_522),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_624),
.B(n_242),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_550),
.B(n_501),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_596),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_563),
.B(n_581),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_547),
.B(n_538),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_596),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_596),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_633),
.B(n_442),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_633),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_567),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_633),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_633),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_548),
.Y(n_718)
);

BUFx10_ASAP7_75t_L g719 ( 
.A(n_588),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_547),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_548),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_590),
.B(n_443),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_549),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_549),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_551),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_551),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_576),
.B(n_503),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_555),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_567),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_603),
.B(n_504),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_555),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_616),
.B(n_506),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_590),
.B(n_443),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_567),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_560),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_560),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_568),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_567),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_568),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_571),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_552),
.A2(n_522),
.B1(n_458),
.B2(n_449),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_552),
.B(n_542),
.Y(n_742)
);

INVx6_ASAP7_75t_L g743 ( 
.A(n_613),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_552),
.B(n_542),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_571),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_556),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_575),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_575),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_592),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_624),
.B(n_445),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_624),
.B(n_445),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_613),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_573),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_613),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_582),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_569),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_594),
.B(n_543),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_595),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_594),
.B(n_543),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_582),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_584),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_616),
.B(n_510),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_585),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_585),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_564),
.B(n_447),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_594),
.B(n_586),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_613),
.Y(n_768)
);

BUFx10_ASAP7_75t_L g769 ( 
.A(n_597),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_586),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_587),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_565),
.B(n_243),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_587),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_589),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_589),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_603),
.B(n_526),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_619),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_632),
.B(n_439),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_591),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_619),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_591),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_605),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_606),
.B(n_539),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_569),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_613),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_606),
.B(n_439),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_566),
.B(n_449),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_565),
.B(n_243),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_600),
.B(n_531),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_613),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_637),
.B(n_598),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_777),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_640),
.B(n_599),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_777),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_695),
.A2(n_703),
.B1(n_706),
.B2(n_681),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_695),
.B(n_417),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_712),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_691),
.B(n_602),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_645),
.B(n_604),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_777),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_661),
.B(n_563),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_690),
.B(n_608),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_636),
.B(n_609),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_636),
.B(n_610),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_681),
.A2(n_565),
.B1(n_623),
.B2(n_619),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_683),
.B(n_625),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_720),
.B(n_450),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_720),
.B(n_627),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_704),
.B(n_630),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_661),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_780),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_663),
.B(n_618),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_721),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_756),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_702),
.B(n_565),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_702),
.B(n_619),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_756),
.Y(n_817)
);

AND2x6_ASAP7_75t_L g818 ( 
.A(n_789),
.B(n_244),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_663),
.B(n_223),
.Y(n_819)
);

NAND2x1_ASAP7_75t_L g820 ( 
.A(n_673),
.B(n_569),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_650),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_787),
.B(n_417),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_660),
.B(n_623),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_750),
.A2(n_572),
.B(n_623),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_780),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_654),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_663),
.B(n_223),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_673),
.B(n_682),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_780),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_787),
.A2(n_474),
.B1(n_295),
.B2(n_246),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_673),
.B(n_248),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_721),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_710),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_786),
.B(n_482),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_660),
.B(n_623),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_710),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_742),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_L g838 ( 
.A1(n_705),
.A2(n_482),
.B1(n_432),
.B2(n_513),
.C(n_493),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_660),
.B(n_605),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_660),
.B(n_679),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_742),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_724),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_744),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_744),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_679),
.B(n_614),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_676),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_679),
.B(n_614),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_681),
.A2(n_249),
.B1(n_261),
.B2(n_244),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_712),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_676),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_679),
.B(n_617),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_673),
.B(n_248),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_787),
.A2(n_249),
.B1(n_262),
.B2(n_261),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_767),
.B(n_617),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_746),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_786),
.B(n_574),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_SL g857 ( 
.A(n_647),
.B(n_257),
.C(n_251),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_712),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_724),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_672),
.B(n_778),
.Y(n_860)
);

AOI22x1_ASAP7_75t_L g861 ( 
.A1(n_708),
.A2(n_262),
.B1(n_296),
.B2(n_278),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_650),
.B(n_626),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_654),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_787),
.A2(n_278),
.B1(n_299),
.B2(n_296),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_681),
.A2(n_706),
.B1(n_703),
.B2(n_787),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_728),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_693),
.B(n_626),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_657),
.B(n_531),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_693),
.B(n_628),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_703),
.B(n_706),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_756),
.B(n_299),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_728),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_642),
.A2(n_421),
.B1(n_425),
.B2(n_418),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_656),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_703),
.B(n_628),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_688),
.B(n_544),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_SL g877 ( 
.A(n_694),
.B(n_749),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_706),
.B(n_718),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_688),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_718),
.B(n_635),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_723),
.B(n_635),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_745),
.Y(n_882)
);

NOR2x1p5_ASAP7_75t_L g883 ( 
.A(n_778),
.B(n_264),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_642),
.A2(n_741),
.B1(n_766),
.B2(n_649),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_723),
.B(n_622),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_682),
.B(n_248),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_725),
.B(n_622),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_698),
.B(n_268),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_757),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_684),
.Y(n_890)
);

INVx5_ASAP7_75t_L g891 ( 
.A(n_756),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_745),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_682),
.B(n_248),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_696),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_725),
.B(n_726),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_772),
.A2(n_310),
.B1(n_314),
.B2(n_301),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_748),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_757),
.A2(n_484),
.B(n_493),
.C(n_432),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_772),
.A2(n_310),
.B1(n_314),
.B2(n_301),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_759),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_698),
.B(n_272),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_759),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_726),
.B(n_622),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_731),
.B(n_622),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_731),
.Y(n_905)
);

BUFx6f_ASAP7_75t_SL g906 ( 
.A(n_662),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_748),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_622),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_735),
.B(n_622),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_772),
.A2(n_320),
.B1(n_340),
.B2(n_316),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_751),
.A2(n_448),
.B(n_447),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_736),
.B(n_583),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_756),
.B(n_316),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_730),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_654),
.B(n_320),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_736),
.B(n_583),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_641),
.B(n_665),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_772),
.B(n_544),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_737),
.B(n_583),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_737),
.B(n_583),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_739),
.B(n_612),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_L g922 ( 
.A(n_667),
.B(n_270),
.Y(n_922)
);

AND2x6_ASAP7_75t_SL g923 ( 
.A(n_727),
.B(n_235),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_682),
.B(n_248),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_SL g925 ( 
.A(n_776),
.B(n_258),
.C(n_226),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_689),
.B(n_784),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_788),
.A2(n_430),
.B1(n_427),
.B2(n_290),
.Y(n_927)
);

AND2x6_ASAP7_75t_SL g928 ( 
.A(n_753),
.B(n_235),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_788),
.B(n_545),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_739),
.B(n_612),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_740),
.B(n_612),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_788),
.A2(n_747),
.B1(n_760),
.B2(n_740),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_747),
.B(n_612),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_788),
.A2(n_373),
.B1(n_429),
.B2(n_358),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_760),
.B(n_545),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_761),
.B(n_340),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_758),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_761),
.B(n_352),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_762),
.B(n_352),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_762),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_722),
.A2(n_572),
.B(n_454),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_713),
.A2(n_354),
.B(n_335),
.C(n_349),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_755),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_689),
.B(n_579),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_666),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_783),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_764),
.B(n_356),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_764),
.B(n_356),
.Y(n_948)
);

AND2x6_ASAP7_75t_SL g949 ( 
.A(n_707),
.B(n_253),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_732),
.B(n_273),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_666),
.A2(n_429),
.B1(n_358),
.B2(n_419),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_765),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_765),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_763),
.B(n_274),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_770),
.B(n_419),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_770),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_689),
.B(n_270),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_771),
.B(n_426),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_709),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_771),
.B(n_426),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_773),
.A2(n_569),
.B1(n_473),
.B2(n_472),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_914),
.B(n_662),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_874),
.B(n_662),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_891),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_799),
.B(n_773),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_791),
.B(n_662),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_793),
.B(n_774),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_802),
.B(n_774),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_858),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_813),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_821),
.B(n_781),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_803),
.B(n_719),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_821),
.B(n_781),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_905),
.B(n_940),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_952),
.B(n_666),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_813),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_884),
.A2(n_668),
.B1(n_700),
.B2(n_684),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_858),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_894),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_832),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_855),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_832),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_SL g983 ( 
.A(n_925),
.B(n_280),
.C(n_277),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_842),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_858),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_855),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_826),
.B(n_668),
.Y(n_987)
);

NAND3xp33_ASAP7_75t_SL g988 ( 
.A(n_830),
.B(n_334),
.C(n_302),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_810),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_874),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_826),
.B(n_668),
.Y(n_991)
);

NAND3xp33_ASAP7_75t_SL g992 ( 
.A(n_946),
.B(n_348),
.C(n_341),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_842),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_870),
.A2(n_711),
.B(n_714),
.C(n_708),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_953),
.B(n_684),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_937),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_859),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_866),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_SL g999 ( 
.A(n_857),
.B(n_689),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_866),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_956),
.B(n_700),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_889),
.B(n_900),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_860),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_801),
.Y(n_1004)
);

AND3x1_ASAP7_75t_SL g1005 ( 
.A(n_883),
.B(n_368),
.C(n_363),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_937),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_872),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_902),
.B(n_700),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_876),
.B(n_719),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_833),
.B(n_836),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_877),
.B(n_719),
.Y(n_1011)
);

NAND2x1p5_ASAP7_75t_L g1012 ( 
.A(n_814),
.B(n_784),
.Y(n_1012)
);

OAI221xp5_ASAP7_75t_L g1013 ( 
.A1(n_838),
.A2(n_901),
.B1(n_888),
.B2(n_834),
.C(n_917),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_863),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_890),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_822),
.B(n_784),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_872),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_882),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_804),
.B(n_719),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_882),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_849),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_892),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_892),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_795),
.B(n_711),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_897),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_801),
.Y(n_1026)
);

CKINVDCx16_ASAP7_75t_R g1027 ( 
.A(n_906),
.Y(n_1027)
);

HAxp5_ASAP7_75t_L g1028 ( 
.A(n_923),
.B(n_361),
.CON(n_1028),
.SN(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_890),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_897),
.Y(n_1030)
);

CKINVDCx11_ASAP7_75t_R g1031 ( 
.A(n_928),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_907),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_907),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_906),
.B(n_769),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_943),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_943),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_890),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_792),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_876),
.B(n_769),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_794),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_895),
.B(n_714),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_SL g1042 ( 
.A1(n_853),
.A2(n_716),
.B(n_717),
.C(n_697),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_906),
.B(n_769),
.Y(n_1043)
);

INVx3_ASAP7_75t_SL g1044 ( 
.A(n_822),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_SL g1045 ( 
.A1(n_856),
.A2(n_374),
.B1(n_404),
.B2(n_364),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_806),
.B(n_716),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_918),
.B(n_769),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_800),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_811),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_822),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_796),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_949),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_796),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_854),
.B(n_717),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_864),
.A2(n_733),
.B1(n_775),
.B2(n_755),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_796),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_918),
.B(n_775),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_849),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_825),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_808),
.B(n_784),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_829),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_837),
.B(n_779),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_841),
.B(n_779),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_840),
.B(n_782),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_935),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_935),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_959),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_878),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_875),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_815),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_807),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_816),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_809),
.B(n_639),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_843),
.B(n_782),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_807),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_891),
.B(n_639),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_844),
.B(n_655),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_849),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_891),
.B(n_639),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_929),
.B(n_638),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_929),
.B(n_638),
.Y(n_1081)
);

AO22x1_ASAP7_75t_L g1082 ( 
.A1(n_818),
.A2(n_667),
.B1(n_256),
.B2(n_259),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_950),
.B(n_283),
.C(n_281),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_954),
.B(n_655),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_846),
.B(n_655),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_932),
.B(n_643),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_863),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_850),
.B(n_655),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_867),
.B(n_643),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_849),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_822),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_879),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_839),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_880),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_915),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_881),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_863),
.B(n_945),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_891),
.Y(n_1098)
);

INVx5_ASAP7_75t_L g1099 ( 
.A(n_891),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_863),
.B(n_945),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_814),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_865),
.B(n_701),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_845),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_847),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_915),
.B(n_664),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_915),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_798),
.B(n_873),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_869),
.B(n_644),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_862),
.A2(n_653),
.B(n_644),
.C(n_652),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_851),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_871),
.B(n_913),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_797),
.B(n_652),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_871),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_823),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_835),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_871),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_911),
.B(n_653),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_885),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_871),
.B(n_664),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_798),
.B(n_868),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_SL g1121 ( 
.A(n_898),
.B(n_292),
.C(n_286),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_887),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_814),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_912),
.B(n_664),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_818),
.B(n_658),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_903),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_L g1127 ( 
.A(n_913),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_936),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_818),
.B(n_658),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_904),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_908),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_938),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_913),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_909),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_927),
.B(n_293),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_939),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_947),
.Y(n_1137)
);

BUFx12f_ASAP7_75t_SL g1138 ( 
.A(n_913),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_916),
.B(n_664),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_948),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_958),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_919),
.B(n_669),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_818),
.B(n_805),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_960),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_820),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_818),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_957),
.Y(n_1148)
);

INVx3_ASAP7_75t_SL g1149 ( 
.A(n_812),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_861),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_818),
.B(n_670),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1012),
.A2(n_824),
.B(n_957),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1117),
.A2(n_827),
.B(n_819),
.Y(n_1153)
);

NAND2x1p5_ASAP7_75t_L g1154 ( 
.A(n_1101),
.B(n_817),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1012),
.A2(n_827),
.B(n_819),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1013),
.B(n_1003),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1058),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1065),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_965),
.B(n_1071),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1065),
.Y(n_1160)
);

AO22x2_ASAP7_75t_L g1161 ( 
.A1(n_988),
.A2(n_256),
.B1(n_259),
.B2(n_253),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1125),
.A2(n_852),
.B(n_831),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1009),
.B(n_1039),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1123),
.A2(n_817),
.B(n_828),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_981),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1009),
.A2(n_920),
.B1(n_930),
.B2(n_921),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1069),
.A2(n_994),
.B(n_1093),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1026),
.B(n_931),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1039),
.B(n_817),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1066),
.A2(n_898),
.B(n_848),
.C(n_942),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_SL g1171 ( 
.A1(n_1107),
.A2(n_933),
.B(n_311),
.C(n_321),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1094),
.B(n_812),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1109),
.A2(n_941),
.B(n_893),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_979),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1075),
.B(n_237),
.Y(n_1175)
);

OAI21xp33_ASAP7_75t_L g1176 ( 
.A1(n_1135),
.A2(n_951),
.B(n_899),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1002),
.B(n_944),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1047),
.A2(n_944),
.B1(n_934),
.B2(n_886),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1096),
.B(n_896),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1066),
.Y(n_1180)
);

NAND2x1_ASAP7_75t_L g1181 ( 
.A(n_1101),
.B(n_651),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_976),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1016),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1129),
.A2(n_893),
.B(n_886),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1151),
.A2(n_924),
.B(n_687),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1123),
.A2(n_926),
.B(n_828),
.Y(n_1186)
);

AOI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_966),
.A2(n_910),
.B(n_924),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1073),
.A2(n_1064),
.B(n_1070),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_979),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1150),
.A2(n_670),
.A3(n_677),
.B(n_678),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_967),
.A2(n_926),
.B1(n_961),
.B2(n_651),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_981),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1123),
.A2(n_639),
.B(n_922),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1047),
.B(n_237),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1015),
.A2(n_1029),
.B(n_978),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1072),
.A2(n_677),
.A3(n_678),
.B(n_692),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1101),
.B(n_1123),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_968),
.B(n_686),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1069),
.A2(n_692),
.B(n_686),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1015),
.A2(n_687),
.B(n_669),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_986),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1015),
.A2(n_687),
.B(n_669),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_984),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1123),
.A2(n_639),
.B(n_922),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1057),
.B(n_701),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1057),
.B(n_646),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1120),
.A2(n_484),
.B(n_513),
.C(n_311),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_980),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1099),
.A2(n_639),
.B(n_659),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1128),
.B(n_646),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1099),
.A2(n_675),
.B(n_659),
.Y(n_1211)
);

AO21x1_ASAP7_75t_L g1212 ( 
.A1(n_999),
.A2(n_321),
.B(n_279),
.Y(n_1212)
);

AOI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1070),
.A2(n_671),
.B(n_648),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_SL g1214 ( 
.A(n_1011),
.B(n_300),
.C(n_298),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_SL g1215 ( 
.A1(n_1144),
.A2(n_667),
.B(n_743),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_984),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1004),
.B(n_303),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1068),
.B(n_648),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1099),
.A2(n_1098),
.B(n_964),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1068),
.B(n_671),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1140),
.B(n_674),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1093),
.B(n_1104),
.Y(n_1222)
);

NAND3x1_ASAP7_75t_L g1223 ( 
.A(n_962),
.B(n_322),
.C(n_279),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1104),
.A2(n_680),
.B(n_674),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_964),
.A2(n_675),
.B(n_659),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1101),
.B(n_669),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1101),
.B(n_687),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1136),
.A2(n_390),
.B(n_322),
.C(n_327),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_964),
.A2(n_715),
.B(n_675),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1058),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1098),
.A2(n_734),
.B(n_715),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1098),
.A2(n_1060),
.B(n_1148),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1058),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1004),
.B(n_237),
.Y(n_1234)
);

NOR2xp67_ASAP7_75t_SL g1235 ( 
.A(n_1147),
.B(n_327),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1072),
.A2(n_416),
.A3(n_331),
.B(n_343),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1024),
.A2(n_699),
.B(n_680),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1148),
.A2(n_734),
.B(n_715),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1058),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1029),
.A2(n_738),
.B(n_729),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1136),
.B(n_1137),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1137),
.B(n_699),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1142),
.A2(n_413),
.A3(n_331),
.B(n_343),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1142),
.B(n_729),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1114),
.A2(n_734),
.B(n_715),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1029),
.A2(n_738),
.B(n_729),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1114),
.A2(n_734),
.B(n_715),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_986),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_969),
.A2(n_738),
.B(n_729),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1102),
.A2(n_738),
.B(n_768),
.Y(n_1250)
);

NAND2x1_ASAP7_75t_L g1251 ( 
.A(n_969),
.B(n_651),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1141),
.B(n_768),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_997),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_990),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1126),
.A2(n_416),
.A3(n_335),
.B(n_346),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1103),
.B(n_768),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1103),
.B(n_768),
.Y(n_1257)
);

AOI21x1_ASAP7_75t_SL g1258 ( 
.A1(n_974),
.A2(n_1001),
.B(n_995),
.Y(n_1258)
);

AO21x1_ASAP7_75t_L g1259 ( 
.A1(n_999),
.A2(n_346),
.B(n_344),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_980),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_972),
.A2(n_390),
.B(n_344),
.C(n_349),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_990),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_997),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1110),
.B(n_790),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_977),
.A2(n_651),
.B1(n_685),
.B2(n_734),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1002),
.B(n_1010),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_969),
.A2(n_985),
.B(n_978),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_996),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1006),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_978),
.A2(n_790),
.B(n_491),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_985),
.A2(n_790),
.B(n_491),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1102),
.A2(n_790),
.B(n_667),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_998),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_993),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_L g1275 ( 
.A(n_983),
.B(n_305),
.C(n_304),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1046),
.A2(n_685),
.B(n_752),
.Y(n_1276)
);

AOI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1019),
.A2(n_313),
.B(n_309),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_985),
.A2(n_491),
.B(n_572),
.Y(n_1278)
);

AOI221x1_ASAP7_75t_L g1279 ( 
.A1(n_1130),
.A2(n_385),
.B1(n_422),
.B2(n_413),
.C(n_354),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1131),
.A2(n_431),
.A3(n_360),
.B(n_422),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1002),
.B(n_237),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1041),
.A2(n_685),
.B(n_754),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1110),
.B(n_667),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1149),
.A2(n_685),
.B1(n_743),
.B2(n_752),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1149),
.A2(n_685),
.B1(n_743),
.B2(n_752),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1145),
.B(n_685),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_993),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1010),
.B(n_241),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1089),
.A2(n_754),
.B(n_752),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1037),
.A2(n_462),
.B(n_448),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_989),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_996),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1145),
.A2(n_431),
.A3(n_360),
.B(n_410),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1132),
.A2(n_743),
.B1(n_754),
.B2(n_752),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1037),
.A2(n_462),
.B(n_454),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1095),
.Y(n_1296)
);

AOI21xp33_ASAP7_75t_L g1297 ( 
.A1(n_1115),
.A2(n_342),
.B(n_338),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1010),
.B(n_241),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1115),
.A2(n_667),
.B(n_473),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1058),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1118),
.A2(n_410),
.A3(n_409),
.B(n_400),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1086),
.A2(n_470),
.B(n_466),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_992),
.A2(n_385),
.B(n_409),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1092),
.B(n_241),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1054),
.A2(n_1132),
.B(n_1062),
.C(n_1127),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1146),
.A2(n_468),
.B(n_466),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1108),
.A2(n_470),
.B(n_468),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1127),
.A2(n_754),
.B1(n_785),
.B2(n_388),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1062),
.B(n_667),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1067),
.B(n_317),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1067),
.B(n_318),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1080),
.A2(n_477),
.B(n_472),
.Y(n_1312)
);

BUFx4_ASAP7_75t_SL g1313 ( 
.A(n_1254),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1174),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1172),
.A2(n_1081),
.B(n_975),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1207),
.A2(n_1055),
.B(n_1112),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1208),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1254),
.Y(n_1318)
);

AOI211xp5_ASAP7_75t_L g1319 ( 
.A1(n_1156),
.A2(n_1045),
.B(n_1052),
.C(n_963),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1305),
.A2(n_1122),
.B(n_1118),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1159),
.B(n_1063),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1215),
.A2(n_1134),
.B(n_1122),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1187),
.A2(n_973),
.B(n_971),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1174),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1159),
.B(n_1063),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1222),
.A2(n_1127),
.B1(n_1106),
.B2(n_1116),
.Y(n_1326)
);

BUFx4f_ASAP7_75t_SL g1327 ( 
.A(n_1268),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1195),
.A2(n_1134),
.B(n_1025),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1241),
.B(n_1063),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1266),
.B(n_987),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1183),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1168),
.A2(n_1052),
.B1(n_1027),
.B2(n_1006),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_SL g1333 ( 
.A(n_1176),
.B(n_1138),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1195),
.A2(n_1025),
.B(n_1018),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1156),
.B(n_1074),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1267),
.A2(n_1033),
.B(n_1018),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1267),
.A2(n_1036),
.B(n_1033),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_SL g1338 ( 
.A(n_1183),
.B(n_1147),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1163),
.B(n_1051),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1163),
.B(n_1050),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_1197),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1213),
.A2(n_1036),
.B(n_1000),
.Y(n_1342)
);

OAI221xp5_ASAP7_75t_L g1343 ( 
.A1(n_1303),
.A2(n_1277),
.B1(n_1311),
.B2(n_1310),
.C(n_1297),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1208),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1161),
.A2(n_1053),
.B1(n_1056),
.B2(n_1050),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1189),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1192),
.B(n_1091),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1305),
.A2(n_1259),
.B(n_1212),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_L g1349 ( 
.A(n_1261),
.B(n_1083),
.C(n_1121),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1210),
.B(n_1074),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1158),
.B(n_1160),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1183),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1260),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1165),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1177),
.B(n_987),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1200),
.A2(n_1240),
.B(n_1202),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1201),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1260),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1274),
.Y(n_1359)
);

CKINVDCx12_ASAP7_75t_R g1360 ( 
.A(n_1234),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1180),
.B(n_1074),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1161),
.A2(n_1008),
.B1(n_1113),
.B2(n_1116),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1200),
.A2(n_1240),
.B(n_1202),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1291),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1207),
.A2(n_1000),
.B(n_998),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1167),
.A2(n_1199),
.B(n_1153),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1279),
.A2(n_1007),
.A3(n_1048),
.B(n_1059),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1274),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1246),
.A2(n_1007),
.B(n_1146),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1161),
.A2(n_1194),
.B1(n_1223),
.B2(n_1177),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1246),
.A2(n_1146),
.B(n_982),
.Y(n_1371)
);

AOI222xp33_ASAP7_75t_L g1372 ( 
.A1(n_1217),
.A2(n_400),
.B1(n_255),
.B2(n_323),
.C1(n_241),
.C2(n_380),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1249),
.A2(n_1017),
.B(n_970),
.Y(n_1373)
);

AO31x2_ASAP7_75t_L g1374 ( 
.A1(n_1261),
.A2(n_1048),
.A3(n_1059),
.B(n_1032),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1287),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1166),
.A2(n_1061),
.B(n_1049),
.C(n_1038),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1223),
.A2(n_1008),
.B1(n_1040),
.B2(n_1044),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_SL g1378 ( 
.A1(n_1169),
.A2(n_1022),
.B(n_1035),
.C(n_1030),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1228),
.A2(n_1028),
.B(n_1044),
.C(n_1042),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1198),
.B(n_1008),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1287),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1248),
.B(n_1310),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1185),
.A2(n_1023),
.B(n_1020),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1179),
.B(n_1113),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1182),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1250),
.A2(n_1139),
.B(n_1124),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1177),
.B(n_987),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1307),
.A2(n_1143),
.B(n_1084),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1249),
.A2(n_1090),
.B(n_1079),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1306),
.A2(n_1090),
.B(n_1076),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1203),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1183),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1296),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1157),
.Y(n_1394)
);

CKINVDCx6p67_ASAP7_75t_R g1395 ( 
.A(n_1262),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1281),
.B(n_1077),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1188),
.A2(n_1021),
.B(n_1078),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1306),
.A2(n_477),
.B(n_378),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1216),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1214),
.A2(n_1298),
.B1(n_1288),
.B2(n_1296),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1217),
.A2(n_1133),
.B1(n_1085),
.B2(n_1077),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1270),
.A2(n_1016),
.B(n_1082),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1262),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1311),
.A2(n_1133),
.B1(n_1085),
.B2(n_1077),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1228),
.A2(n_415),
.B1(n_355),
.B2(n_359),
.C(n_365),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1178),
.A2(n_1088),
.B(n_1085),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1197),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1270),
.A2(n_1016),
.B(n_1082),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1271),
.A2(n_1016),
.B(n_1111),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1271),
.A2(n_1278),
.B(n_1185),
.Y(n_1410)
);

INVx8_ASAP7_75t_L g1411 ( 
.A(n_1157),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1205),
.B(n_1088),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1230),
.B(n_991),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1206),
.B(n_1088),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1253),
.B(n_1105),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1292),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1278),
.A2(n_1111),
.B(n_1078),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1237),
.A2(n_1100),
.B(n_1097),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1275),
.B(n_411),
.C(n_333),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1230),
.Y(n_1420)
);

NOR2xp67_ASAP7_75t_L g1421 ( 
.A(n_1239),
.B(n_1021),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1154),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1269),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1263),
.B(n_1105),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1175),
.A2(n_1138),
.B1(n_1105),
.B2(n_991),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1239),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1154),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1155),
.A2(n_1111),
.B(n_1005),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1273),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1290),
.A2(n_1111),
.B(n_1100),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1295),
.A2(n_1100),
.B(n_1097),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1269),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1218),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1272),
.A2(n_1097),
.B(n_1119),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1191),
.A2(n_991),
.B(n_1119),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1220),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1299),
.A2(n_1119),
.B(n_1043),
.Y(n_1437)
);

AO31x2_ASAP7_75t_L g1438 ( 
.A1(n_1170),
.A2(n_1028),
.A3(n_270),
.B(n_1087),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1196),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1169),
.B(n_1014),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1164),
.B(n_1232),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1221),
.A2(n_1087),
.B1(n_1014),
.B2(n_398),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1196),
.Y(n_1443)
);

AOI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1304),
.A2(n_389),
.B(n_428),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_SL g1445 ( 
.A1(n_1170),
.A2(n_1034),
.B(n_270),
.C(n_135),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1152),
.A2(n_785),
.B(n_754),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1242),
.B(n_330),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1244),
.B(n_336),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1152),
.A2(n_785),
.B(n_270),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1196),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1196),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1309),
.A2(n_396),
.B1(n_351),
.B2(n_424),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1312),
.A2(n_387),
.B(n_366),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1258),
.A2(n_785),
.B(n_270),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1162),
.A2(n_401),
.B(n_376),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1256),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1243),
.B(n_255),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1252),
.B(n_381),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1162),
.A2(n_215),
.B(n_210),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1184),
.A2(n_202),
.B(n_201),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1235),
.A2(n_255),
.B1(n_323),
.B2(n_1031),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1302),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1184),
.A2(n_199),
.B(n_198),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1224),
.A2(n_423),
.B(n_407),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1243),
.B(n_255),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1257),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1233),
.Y(n_1467)
);

AOI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1302),
.A2(n_155),
.B(n_196),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1219),
.A2(n_190),
.B(n_188),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1186),
.A2(n_187),
.B(n_178),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1233),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1190),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1226),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1302),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1300),
.B(n_176),
.Y(n_1475)
);

AO21x2_ASAP7_75t_L g1476 ( 
.A1(n_1286),
.A2(n_171),
.B(n_170),
.Y(n_1476)
);

OR2x6_ASAP7_75t_L g1477 ( 
.A(n_1300),
.B(n_166),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1283),
.A2(n_406),
.B1(n_403),
.B2(n_386),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1282),
.A2(n_161),
.B(n_158),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1264),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1286),
.B(n_323),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1308),
.A2(n_323),
.B1(n_1031),
.B2(n_20),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1289),
.A2(n_150),
.B(n_147),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1357),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1343),
.A2(n_1265),
.B1(n_1251),
.B2(n_1276),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1372),
.A2(n_1173),
.B1(n_1245),
.B2(n_1247),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1335),
.B(n_1255),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1382),
.A2(n_1285),
.B1(n_1284),
.B2(n_1294),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1357),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1400),
.A2(n_1226),
.B1(n_1227),
.B2(n_1238),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1372),
.A2(n_1173),
.B1(n_1227),
.B2(n_1181),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1330),
.B(n_1243),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1327),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1321),
.B(n_1325),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1330),
.B(n_1301),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1333),
.A2(n_1173),
.B1(n_19),
.B2(n_21),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1333),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1482),
.A2(n_1243),
.B1(n_1236),
.B2(n_1255),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1423),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1329),
.B(n_1280),
.Y(n_1500)
);

CKINVDCx16_ASAP7_75t_R g1501 ( 
.A(n_1318),
.Y(n_1501)
);

INVx4_ASAP7_75t_SL g1502 ( 
.A(n_1331),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1330),
.B(n_1236),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1384),
.B(n_23),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1397),
.A2(n_1231),
.B(n_1225),
.Y(n_1505)
);

INVx3_ASAP7_75t_SL g1506 ( 
.A(n_1403),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1347),
.B(n_1384),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1350),
.B(n_1280),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1444),
.A2(n_1229),
.B1(n_1193),
.B2(n_1204),
.C(n_1255),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1477),
.B(n_1211),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1347),
.B(n_1280),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1385),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1339),
.B(n_1280),
.Y(n_1513)
);

OR2x6_ASAP7_75t_SL g1514 ( 
.A(n_1403),
.B(n_1255),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1441),
.A2(n_1209),
.B(n_1171),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1457),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1516)
);

AOI21xp33_ASAP7_75t_L g1517 ( 
.A1(n_1453),
.A2(n_1236),
.B(n_1293),
.Y(n_1517)
);

A2O1A1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1379),
.A2(n_1236),
.B(n_1293),
.C(n_1301),
.Y(n_1518)
);

CKINVDCx11_ASAP7_75t_R g1519 ( 
.A(n_1395),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1404),
.A2(n_1293),
.B1(n_1301),
.B2(n_1190),
.Y(n_1520)
);

AND2x6_ASAP7_75t_L g1521 ( 
.A(n_1392),
.B(n_1301),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1446),
.A2(n_1190),
.B(n_1293),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1370),
.B(n_1190),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1324),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1423),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1396),
.B(n_25),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1385),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1392),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1392),
.Y(n_1529)
);

CKINVDCx6p67_ASAP7_75t_R g1530 ( 
.A(n_1360),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1349),
.A2(n_28),
.B1(n_31),
.B2(n_40),
.Y(n_1531)
);

INVxp33_ASAP7_75t_L g1532 ( 
.A(n_1314),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1330),
.B(n_144),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1349),
.A2(n_1465),
.B1(n_1457),
.B2(n_1370),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1393),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1324),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1461),
.A2(n_28),
.B1(n_31),
.B2(n_41),
.C(n_48),
.Y(n_1537)
);

CKINVDCx8_ASAP7_75t_R g1538 ( 
.A(n_1346),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1405),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.C(n_56),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1391),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1401),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_1541)
);

NAND4xp25_ASAP7_75t_L g1542 ( 
.A(n_1319),
.B(n_60),
.C(n_61),
.D(n_62),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1391),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1441),
.A2(n_142),
.B(n_140),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1416),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1377),
.A2(n_1380),
.B1(n_1447),
.B2(n_1477),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1377),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1416),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1446),
.A2(n_139),
.B(n_134),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1360),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1477),
.B(n_131),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1425),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_1552)
);

OAI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1319),
.A2(n_69),
.B(n_71),
.C(n_72),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1465),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1346),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1396),
.B(n_74),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1392),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1472),
.A2(n_76),
.B(n_78),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1313),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_SL g1560 ( 
.A1(n_1406),
.A2(n_78),
.B(n_80),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1361),
.B(n_80),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1413),
.B(n_130),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1445),
.A2(n_83),
.B1(n_86),
.B2(n_89),
.C(n_90),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1399),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1441),
.A2(n_97),
.B(n_114),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1429),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1340),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1429),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1361),
.B(n_94),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1399),
.Y(n_1570)
);

AOI21xp33_ASAP7_75t_L g1571 ( 
.A1(n_1452),
.A2(n_95),
.B(n_119),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1441),
.A2(n_1366),
.B(n_1435),
.Y(n_1572)
);

CKINVDCx16_ASAP7_75t_R g1573 ( 
.A(n_1432),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1392),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1352),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_R g1576 ( 
.A(n_1418),
.B(n_1316),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1353),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1351),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1354),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1351),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1364),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1331),
.Y(n_1582)
);

INVx6_ASAP7_75t_L g1583 ( 
.A(n_1331),
.Y(n_1583)
);

AO31x2_ASAP7_75t_L g1584 ( 
.A1(n_1472),
.A2(n_1451),
.A3(n_1450),
.B(n_1439),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1413),
.B(n_1355),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1317),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1364),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1317),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1344),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1340),
.A2(n_1323),
.B1(n_1419),
.B2(n_1316),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1419),
.A2(n_1316),
.B1(n_1345),
.B2(n_1362),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1432),
.A2(n_1332),
.B1(n_1326),
.B2(n_1447),
.Y(n_1592)
);

INVx5_ASAP7_75t_L g1593 ( 
.A(n_1331),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1433),
.B(n_1436),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1418),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1462),
.A2(n_1474),
.B(n_1451),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1462),
.A2(n_1474),
.B(n_1439),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1413),
.B(n_1355),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1355),
.B(n_1387),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1344),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1358),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1433),
.B(n_1436),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1315),
.B(n_1376),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1413),
.B(n_1355),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1358),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1477),
.A2(n_1437),
.B1(n_1316),
.B2(n_1455),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1353),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1359),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1359),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1394),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1381),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1458),
.B(n_1448),
.Y(n_1612)
);

OR2x6_ASAP7_75t_L g1613 ( 
.A(n_1477),
.B(n_1352),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1478),
.A2(n_1481),
.B1(n_1442),
.B2(n_1320),
.C(n_1480),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1368),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1387),
.A2(n_1352),
.B1(n_1440),
.B2(n_1422),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1467),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1381),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1412),
.B(n_1414),
.Y(n_1619)
);

AOI222xp33_ASAP7_75t_L g1620 ( 
.A1(n_1412),
.A2(n_1414),
.B1(n_1387),
.B2(n_1424),
.C1(n_1415),
.C2(n_1456),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1387),
.A2(n_1466),
.B1(n_1456),
.B2(n_1415),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1622)
);

AOI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1320),
.A2(n_1466),
.B1(n_1378),
.B2(n_1368),
.C(n_1375),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1411),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1475),
.A2(n_1437),
.B1(n_1338),
.B2(n_1434),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1375),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1438),
.B(n_1475),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1322),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_SL g1629 ( 
.A(n_1440),
.B(n_1450),
.C(n_1443),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1464),
.A2(n_1348),
.B1(n_1366),
.B2(n_1434),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1394),
.Y(n_1631)
);

AOI31xp67_ASAP7_75t_L g1632 ( 
.A1(n_1443),
.A2(n_1475),
.A3(n_1348),
.B(n_1388),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1438),
.B(n_1475),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1418),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1438),
.B(n_1420),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1464),
.A2(n_1440),
.B1(n_1341),
.B2(n_1338),
.C(n_1365),
.Y(n_1636)
);

NOR2xp67_ASAP7_75t_L g1637 ( 
.A(n_1407),
.B(n_1473),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1426),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1418),
.A2(n_1407),
.B1(n_1421),
.B2(n_1427),
.Y(n_1639)
);

OAI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1464),
.A2(n_1365),
.B1(n_1427),
.B2(n_1407),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1322),
.Y(n_1641)
);

AND2x2_ASAP7_75t_SL g1642 ( 
.A(n_1464),
.B(n_1365),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1426),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1348),
.A2(n_1366),
.B1(n_1434),
.B2(n_1365),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1421),
.A2(n_1427),
.B1(n_1473),
.B2(n_1426),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1473),
.A2(n_1426),
.B1(n_1420),
.B2(n_1471),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1374),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1397),
.A2(n_1437),
.B1(n_1386),
.B2(n_1476),
.C(n_1438),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1374),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1470),
.A2(n_1479),
.B(n_1428),
.C(n_1483),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1386),
.A2(n_1428),
.B1(n_1476),
.B2(n_1388),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1438),
.B(n_1420),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1476),
.A2(n_1386),
.B1(n_1388),
.B2(n_1470),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1426),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1479),
.A2(n_1483),
.B1(n_1471),
.B2(n_1383),
.Y(n_1655)
);

AO21x2_ASAP7_75t_L g1656 ( 
.A1(n_1410),
.A2(n_1449),
.B(n_1363),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1374),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_SL g1658 ( 
.A(n_1471),
.B(n_1383),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1374),
.B(n_1411),
.Y(n_1659)
);

AOI22x1_ASAP7_75t_L g1660 ( 
.A1(n_1374),
.A2(n_1367),
.B1(n_1469),
.B2(n_1463),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1411),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1542),
.A2(n_1411),
.B1(n_1468),
.B2(n_1383),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1635),
.B(n_1367),
.Y(n_1663)
);

INVx11_ASAP7_75t_L g1664 ( 
.A(n_1521),
.Y(n_1664)
);

AOI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1537),
.A2(n_1547),
.B(n_1553),
.C(n_1592),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1539),
.A2(n_1411),
.B1(n_1430),
.B2(n_1469),
.Y(n_1666)
);

OAI222xp33_ASAP7_75t_L g1667 ( 
.A1(n_1531),
.A2(n_1468),
.B1(n_1367),
.B2(n_1430),
.C1(n_1459),
.C2(n_1463),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1494),
.B(n_1367),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1531),
.A2(n_1409),
.B1(n_1459),
.B2(n_1460),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1612),
.A2(n_1383),
.B1(n_1460),
.B2(n_1409),
.C(n_1367),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1603),
.A2(n_1408),
.B(n_1402),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1513),
.B(n_1454),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1573),
.B(n_1501),
.Y(n_1673)
);

CKINVDCx11_ASAP7_75t_R g1674 ( 
.A(n_1519),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1524),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1538),
.A2(n_1431),
.B1(n_1408),
.B2(n_1402),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1563),
.A2(n_1547),
.B1(n_1571),
.B2(n_1554),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1554),
.A2(n_1431),
.B1(n_1417),
.B2(n_1454),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1614),
.A2(n_1398),
.B(n_1417),
.Y(n_1679)
);

A2O1A1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1496),
.A2(n_1328),
.B(n_1373),
.C(n_1342),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1560),
.A2(n_1390),
.B1(n_1371),
.B2(n_1369),
.Y(n_1681)
);

OA21x2_ASAP7_75t_L g1682 ( 
.A1(n_1518),
.A2(n_1410),
.B(n_1363),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1497),
.A2(n_1371),
.B1(n_1389),
.B2(n_1369),
.C(n_1337),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1545),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1567),
.A2(n_1389),
.B1(n_1336),
.B2(n_1337),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1540),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1627),
.B(n_1633),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_SL g1688 ( 
.A1(n_1594),
.A2(n_1356),
.B(n_1334),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1567),
.A2(n_1516),
.B1(n_1497),
.B2(n_1534),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1534),
.A2(n_1334),
.B1(n_1336),
.B2(n_1356),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1546),
.B(n_1620),
.Y(n_1691)
);

AOI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1658),
.A2(n_1520),
.B(n_1515),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1652),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1617),
.A2(n_1621),
.B1(n_1530),
.B2(n_1551),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1621),
.A2(n_1551),
.B1(n_1506),
.B2(n_1550),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1516),
.A2(n_1496),
.B1(n_1504),
.B2(n_1541),
.C(n_1591),
.Y(n_1696)
);

NOR2x1p5_ASAP7_75t_L g1697 ( 
.A(n_1582),
.B(n_1559),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1546),
.A2(n_1552),
.B1(n_1551),
.B2(n_1504),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1533),
.A2(n_1599),
.B1(n_1613),
.B2(n_1562),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1492),
.A2(n_1503),
.B1(n_1495),
.B2(n_1533),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1619),
.B(n_1523),
.Y(n_1701)
);

OAI332xp33_ASAP7_75t_L g1702 ( 
.A1(n_1507),
.A2(n_1569),
.A3(n_1561),
.B1(n_1556),
.B2(n_1526),
.B3(n_1511),
.C1(n_1487),
.C2(n_1488),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1543),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1544),
.A2(n_1565),
.B1(n_1613),
.B2(n_1593),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1517),
.A2(n_1498),
.B1(n_1591),
.B2(n_1532),
.C(n_1485),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1498),
.A2(n_1532),
.B1(n_1485),
.B2(n_1590),
.C(n_1535),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1508),
.B(n_1500),
.Y(n_1707)
);

OAI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1613),
.A2(n_1506),
.B1(n_1625),
.B2(n_1514),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1495),
.B(n_1585),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1606),
.A2(n_1590),
.B1(n_1486),
.B2(n_1491),
.C(n_1535),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1548),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1599),
.A2(n_1585),
.B1(n_1598),
.B2(n_1604),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1587),
.A2(n_1525),
.B1(n_1499),
.B2(n_1555),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1606),
.A2(n_1636),
.B(n_1650),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1523),
.B(n_1578),
.Y(n_1715)
);

CKINVDCx6p67_ASAP7_75t_R g1716 ( 
.A(n_1493),
.Y(n_1716)
);

BUFx4f_ASAP7_75t_SL g1717 ( 
.A(n_1484),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1524),
.A2(n_1536),
.B(n_1486),
.C(n_1630),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1593),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1598),
.A2(n_1604),
.B1(n_1562),
.B2(n_1579),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1489),
.Y(n_1721)
);

A2O1A1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1518),
.A2(n_1623),
.B(n_1648),
.C(n_1491),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1536),
.A2(n_1640),
.B1(n_1630),
.B2(n_1490),
.C(n_1644),
.Y(n_1723)
);

OAI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1581),
.A2(n_1510),
.B1(n_1593),
.B2(n_1602),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1510),
.A2(n_1624),
.B1(n_1616),
.B2(n_1582),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_SL g1726 ( 
.A1(n_1558),
.A2(n_1642),
.B1(n_1583),
.B2(n_1510),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1584),
.B(n_1647),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1640),
.A2(n_1644),
.B1(n_1653),
.B2(n_1580),
.C(n_1509),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1622),
.A2(n_1521),
.B1(n_1583),
.B2(n_1659),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1622),
.A2(n_1521),
.B1(n_1583),
.B2(n_1575),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_SL g1731 ( 
.A1(n_1558),
.A2(n_1642),
.B1(n_1521),
.B2(n_1575),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1595),
.B(n_1634),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1502),
.B(n_1529),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1595),
.B(n_1634),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1653),
.A2(n_1657),
.B1(n_1649),
.B2(n_1639),
.C(n_1570),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1522),
.A2(n_1650),
.B(n_1660),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1521),
.A2(n_1575),
.B1(n_1629),
.B2(n_1610),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1575),
.A2(n_1629),
.B1(n_1564),
.B2(n_1512),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1527),
.A2(n_1566),
.B1(n_1568),
.B2(n_1529),
.Y(n_1739)
);

OA21x2_ASAP7_75t_L g1740 ( 
.A1(n_1651),
.A2(n_1655),
.B(n_1641),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1631),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1528),
.A2(n_1557),
.B1(n_1574),
.B2(n_1558),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1577),
.B(n_1607),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1528),
.A2(n_1557),
.B1(n_1574),
.B2(n_1654),
.Y(n_1744)
);

AO21x1_ASAP7_75t_SL g1745 ( 
.A1(n_1657),
.A2(n_1655),
.B(n_1589),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1637),
.A2(n_1661),
.B1(n_1646),
.B2(n_1645),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1654),
.A2(n_1626),
.B1(n_1588),
.B2(n_1615),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1586),
.B(n_1608),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1600),
.A2(n_1609),
.B1(n_1605),
.B2(n_1601),
.Y(n_1749)
);

AOI222xp33_ASAP7_75t_L g1750 ( 
.A1(n_1502),
.A2(n_1618),
.B1(n_1611),
.B2(n_1661),
.C1(n_1643),
.C2(n_1638),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1576),
.A2(n_1643),
.B1(n_1638),
.B2(n_1628),
.C(n_1596),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1505),
.A2(n_1638),
.B1(n_1576),
.B2(n_1656),
.C(n_1632),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1505),
.A2(n_1638),
.B1(n_1656),
.B2(n_1502),
.C(n_1549),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1597),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1597),
.A2(n_1013),
.B1(n_637),
.B2(n_1343),
.C(n_1547),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1597),
.A2(n_799),
.B(n_1013),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1542),
.A2(n_1343),
.B1(n_1013),
.B2(n_1537),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1513),
.B(n_1652),
.Y(n_1761)
);

OAI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1531),
.A2(n_1343),
.B1(n_1013),
.B2(n_799),
.C(n_802),
.Y(n_1762)
);

AO21x2_ASAP7_75t_L g1763 ( 
.A1(n_1650),
.A2(n_1640),
.B(n_1517),
.Y(n_1763)
);

BUFx4f_ASAP7_75t_SL g1764 ( 
.A(n_1617),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1765)
);

A2O1A1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1563),
.A2(n_1013),
.B(n_1176),
.C(n_799),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1545),
.Y(n_1767)
);

AOI222xp33_ASAP7_75t_L g1768 ( 
.A1(n_1539),
.A2(n_988),
.B1(n_1045),
.B2(n_925),
.C1(n_1013),
.C2(n_1531),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1635),
.B(n_1627),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1538),
.A2(n_1343),
.B1(n_799),
.B2(n_1013),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1524),
.Y(n_1771)
);

AO221x2_ASAP7_75t_L g1772 ( 
.A1(n_1547),
.A2(n_1546),
.B1(n_1592),
.B2(n_1541),
.C(n_1045),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1603),
.A2(n_799),
.B(n_1572),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1495),
.B(n_1613),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1539),
.B(n_799),
.C(n_1013),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_SL g1777 ( 
.A1(n_1553),
.A2(n_1343),
.B1(n_799),
.B2(n_1013),
.Y(n_1777)
);

AOI22x1_ASAP7_75t_L g1778 ( 
.A1(n_1560),
.A2(n_1372),
.B1(n_914),
.B2(n_1161),
.Y(n_1778)
);

OAI221xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1531),
.A2(n_1372),
.B1(n_1343),
.B2(n_1482),
.C(n_1013),
.Y(n_1779)
);

OR2x6_ASAP7_75t_L g1780 ( 
.A(n_1613),
.B(n_1572),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1539),
.B(n_799),
.C(n_1013),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1538),
.A2(n_1343),
.B1(n_799),
.B2(n_1013),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1542),
.A2(n_1343),
.B1(n_1013),
.B2(n_1537),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1635),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1635),
.B(n_1627),
.Y(n_1785)
);

OAI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1531),
.A2(n_1343),
.B1(n_1013),
.B2(n_799),
.C(n_802),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1787)
);

AO21x1_ASAP7_75t_L g1788 ( 
.A1(n_1603),
.A2(n_1547),
.B(n_1546),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1538),
.A2(n_1343),
.B1(n_799),
.B2(n_1013),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1792)
);

OA21x2_ASAP7_75t_L g1793 ( 
.A1(n_1518),
.A2(n_1648),
.B(n_1522),
.Y(n_1793)
);

OAI21xp33_ASAP7_75t_L g1794 ( 
.A1(n_1531),
.A2(n_637),
.B(n_799),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1795)
);

AOI222xp33_ASAP7_75t_L g1796 ( 
.A1(n_1539),
.A2(n_988),
.B1(n_1045),
.B2(n_925),
.C1(n_1013),
.C2(n_1531),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1539),
.A2(n_1343),
.B1(n_1013),
.B2(n_988),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1538),
.A2(n_1343),
.B1(n_799),
.B2(n_1013),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1504),
.B(n_1372),
.C(n_637),
.D(n_1156),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1547),
.A2(n_1013),
.B1(n_637),
.B2(n_1343),
.C(n_1537),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1635),
.B(n_1627),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1531),
.A2(n_1343),
.B1(n_1013),
.B2(n_799),
.C(n_802),
.Y(n_1803)
);

AOI222xp33_ASAP7_75t_L g1804 ( 
.A1(n_1539),
.A2(n_988),
.B1(n_1045),
.B2(n_925),
.C1(n_1013),
.C2(n_1531),
.Y(n_1804)
);

OAI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1542),
.A2(n_1343),
.B1(n_1013),
.B2(n_1537),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1559),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1547),
.A2(n_1013),
.B1(n_637),
.B2(n_1343),
.C(n_1537),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1772),
.A2(n_1794),
.B1(n_1800),
.B2(n_1796),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1663),
.B(n_1687),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1780),
.B(n_1774),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1754),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1663),
.B(n_1687),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1761),
.B(n_1732),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1769),
.B(n_1785),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1769),
.B(n_1785),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1727),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1727),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1732),
.Y(n_1818)
);

AOI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1779),
.A2(n_1801),
.B1(n_1807),
.B2(n_1803),
.C(n_1786),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1664),
.Y(n_1820)
);

NOR4xp25_ASAP7_75t_SL g1821 ( 
.A(n_1762),
.B(n_1755),
.C(n_1791),
.D(n_1766),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1664),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1675),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1780),
.B(n_1774),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1802),
.B(n_1734),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1707),
.B(n_1668),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1707),
.B(n_1761),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1772),
.A2(n_1804),
.B1(n_1768),
.B2(n_1775),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1771),
.B(n_1701),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1770),
.B(n_1782),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1684),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1802),
.B(n_1734),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1715),
.B(n_1784),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1688),
.Y(n_1834)
);

AOI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1781),
.A2(n_1783),
.B(n_1757),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1684),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1780),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1688),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1764),
.B(n_1673),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1693),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1686),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1703),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1701),
.B(n_1773),
.Y(n_1843)
);

AO21x2_ASAP7_75t_L g1844 ( 
.A1(n_1722),
.A2(n_1714),
.B(n_1679),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1674),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1793),
.B(n_1740),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1672),
.B(n_1793),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1672),
.B(n_1740),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1731),
.B(n_1745),
.Y(n_1849)
);

OAI211xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1777),
.A2(n_1789),
.B(n_1795),
.C(n_1758),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1745),
.B(n_1763),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1748),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1763),
.B(n_1726),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1763),
.B(n_1752),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1670),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1728),
.B(n_1682),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1671),
.B(n_1709),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1682),
.B(n_1692),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1682),
.B(n_1723),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1735),
.B(n_1736),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1751),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1690),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1724),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1743),
.Y(n_1864)
);

AOI21xp33_ASAP7_75t_L g1865 ( 
.A1(n_1805),
.A2(n_1790),
.B(n_1799),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1736),
.B(n_1722),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1736),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1683),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1766),
.A2(n_1756),
.B(n_1791),
.Y(n_1869)
);

OR2x6_ASAP7_75t_L g1870 ( 
.A(n_1788),
.B(n_1676),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1709),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1749),
.Y(n_1872)
);

OR2x6_ASAP7_75t_L g1873 ( 
.A(n_1788),
.B(n_1691),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1680),
.B(n_1705),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1710),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1680),
.B(n_1685),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1681),
.B(n_1691),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1706),
.B(n_1702),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1772),
.A2(n_1677),
.B1(n_1689),
.B2(n_1696),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1828),
.A2(n_1765),
.B1(n_1792),
.B2(n_1760),
.C(n_1798),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1819),
.A2(n_1759),
.B1(n_1797),
.B2(n_1787),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1841),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1829),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1829),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1865),
.A2(n_1776),
.B(n_1698),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1819),
.A2(n_1778),
.B1(n_1694),
.B2(n_1695),
.Y(n_1886)
);

OAI31xp33_ASAP7_75t_L g1887 ( 
.A1(n_1828),
.A2(n_1708),
.A3(n_1662),
.B(n_1718),
.Y(n_1887)
);

BUFx3_ASAP7_75t_L g1888 ( 
.A(n_1831),
.Y(n_1888)
);

OAI31xp33_ASAP7_75t_L g1889 ( 
.A1(n_1850),
.A2(n_1725),
.A3(n_1713),
.B(n_1746),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1841),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1831),
.Y(n_1891)
);

AOI222xp33_ASAP7_75t_L g1892 ( 
.A1(n_1808),
.A2(n_1711),
.B1(n_1665),
.B2(n_1721),
.C1(n_1767),
.C2(n_1717),
.Y(n_1892)
);

NAND4xp25_ASAP7_75t_L g1893 ( 
.A(n_1808),
.B(n_1767),
.C(n_1739),
.D(n_1747),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1830),
.A2(n_1719),
.B1(n_1741),
.B2(n_1733),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1841),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1842),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1830),
.A2(n_1704),
.B1(n_1699),
.B2(n_1720),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1809),
.B(n_1729),
.Y(n_1898)
);

OAI31xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1865),
.A2(n_1733),
.A3(n_1753),
.B(n_1750),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1879),
.A2(n_1700),
.B1(n_1712),
.B2(n_1730),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1809),
.B(n_1737),
.Y(n_1901)
);

INVxp67_ASAP7_75t_SL g1902 ( 
.A(n_1811),
.Y(n_1902)
);

AOI31xp33_ASAP7_75t_L g1903 ( 
.A1(n_1879),
.A2(n_1806),
.A3(n_1738),
.B(n_1666),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1835),
.A2(n_1697),
.B1(n_1716),
.B2(n_1674),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1835),
.A2(n_1716),
.B1(n_1669),
.B2(n_1733),
.Y(n_1905)
);

OAI21xp33_ASAP7_75t_L g1906 ( 
.A1(n_1873),
.A2(n_1742),
.B(n_1678),
.Y(n_1906)
);

CKINVDCx16_ASAP7_75t_R g1907 ( 
.A(n_1839),
.Y(n_1907)
);

AOI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1867),
.A2(n_1667),
.B(n_1744),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_R g1909 ( 
.A(n_1845),
.B(n_1806),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_R g1910 ( 
.A(n_1836),
.B(n_1820),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1827),
.B(n_1826),
.Y(n_1911)
);

OAI33xp33_ASAP7_75t_L g1912 ( 
.A1(n_1878),
.A2(n_1850),
.A3(n_1843),
.B1(n_1823),
.B2(n_1816),
.B3(n_1817),
.Y(n_1912)
);

OAI221xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1873),
.A2(n_1878),
.B1(n_1869),
.B2(n_1870),
.C(n_1875),
.Y(n_1913)
);

OA21x2_ASAP7_75t_L g1914 ( 
.A1(n_1867),
.A2(n_1858),
.B(n_1846),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1840),
.Y(n_1915)
);

AO21x2_ASAP7_75t_L g1916 ( 
.A1(n_1867),
.A2(n_1854),
.B(n_1858),
.Y(n_1916)
);

AOI31xp33_ASAP7_75t_L g1917 ( 
.A1(n_1869),
.A2(n_1875),
.A3(n_1877),
.B(n_1874),
.Y(n_1917)
);

OAI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1858),
.A2(n_1834),
.B(n_1838),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1840),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1836),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1827),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1818),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1816),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1813),
.Y(n_1924)
);

NAND3xp33_ASAP7_75t_L g1925 ( 
.A(n_1821),
.B(n_1873),
.C(n_1855),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1846),
.A2(n_1854),
.B(n_1851),
.Y(n_1926)
);

AOI222xp33_ASAP7_75t_L g1927 ( 
.A1(n_1874),
.A2(n_1877),
.B1(n_1821),
.B2(n_1876),
.C1(n_1843),
.C2(n_1856),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1826),
.B(n_1864),
.Y(n_1928)
);

AO21x2_ASAP7_75t_L g1929 ( 
.A1(n_1854),
.A2(n_1846),
.B(n_1844),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_R g1930 ( 
.A(n_1853),
.B(n_1849),
.Y(n_1930)
);

AND4x1_ASAP7_75t_L g1931 ( 
.A(n_1874),
.B(n_1877),
.C(n_1853),
.D(n_1876),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1817),
.Y(n_1932)
);

BUFx2_ASAP7_75t_L g1933 ( 
.A(n_1810),
.Y(n_1933)
);

AOI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1855),
.A2(n_1861),
.B1(n_1868),
.B2(n_1844),
.C(n_1856),
.Y(n_1934)
);

NAND4xp25_ASAP7_75t_SL g1935 ( 
.A(n_1853),
.B(n_1876),
.C(n_1849),
.D(n_1856),
.Y(n_1935)
);

AOI221xp5_ASAP7_75t_L g1936 ( 
.A1(n_1861),
.A2(n_1868),
.B1(n_1844),
.B2(n_1862),
.C(n_1859),
.Y(n_1936)
);

OA21x2_ASAP7_75t_L g1937 ( 
.A1(n_1851),
.A2(n_1866),
.B(n_1868),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1873),
.A2(n_1844),
.B1(n_1870),
.B2(n_1872),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1818),
.Y(n_1939)
);

OAI21x1_ASAP7_75t_L g1940 ( 
.A1(n_1834),
.A2(n_1838),
.B(n_1866),
.Y(n_1940)
);

OAI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1873),
.A2(n_1870),
.B1(n_1863),
.B2(n_1872),
.C(n_1862),
.Y(n_1941)
);

NAND3xp33_ASAP7_75t_L g1942 ( 
.A(n_1870),
.B(n_1863),
.C(n_1866),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1924),
.B(n_1813),
.Y(n_1943)
);

AOI33xp33_ASAP7_75t_L g1944 ( 
.A1(n_1938),
.A2(n_1934),
.A3(n_1881),
.B1(n_1936),
.B2(n_1886),
.B3(n_1859),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1929),
.B(n_1813),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1929),
.B(n_1847),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1882),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1914),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1933),
.B(n_1809),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1914),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1933),
.B(n_1812),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1926),
.B(n_1812),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1929),
.B(n_1926),
.Y(n_1953)
);

INVxp67_ASAP7_75t_SL g1954 ( 
.A(n_1937),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1921),
.B(n_1883),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1884),
.B(n_1823),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1914),
.Y(n_1957)
);

INVxp67_ASAP7_75t_SL g1958 ( 
.A(n_1937),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1928),
.B(n_1811),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1882),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1890),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1940),
.B(n_1857),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1890),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1895),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1915),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1940),
.B(n_1857),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1914),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1926),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1907),
.B(n_1871),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1919),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1926),
.B(n_1812),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1922),
.B(n_1849),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1895),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1896),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1939),
.B(n_1825),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1937),
.B(n_1825),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1902),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1911),
.B(n_1871),
.Y(n_1978)
);

NAND2x1_ASAP7_75t_L g1979 ( 
.A(n_1937),
.B(n_1857),
.Y(n_1979)
);

AND2x4_ASAP7_75t_SL g1980 ( 
.A(n_1897),
.B(n_1820),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1901),
.B(n_1825),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1901),
.B(n_1832),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1918),
.B(n_1857),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1888),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1923),
.B(n_1832),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1880),
.B(n_1917),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1893),
.B(n_1871),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1898),
.B(n_1832),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1898),
.B(n_1833),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1923),
.B(n_1852),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1918),
.B(n_1857),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1916),
.B(n_1847),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1888),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1916),
.B(n_1833),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1942),
.B(n_1810),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1932),
.B(n_1852),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1916),
.B(n_1847),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1945),
.B(n_1943),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1948),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1987),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1947),
.Y(n_2001)
);

AO21x1_ASAP7_75t_L g2002 ( 
.A1(n_1986),
.A2(n_1930),
.B(n_1887),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1948),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1978),
.B(n_1927),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1952),
.B(n_1931),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1947),
.Y(n_2006)
);

NOR2x1_ASAP7_75t_SL g2007 ( 
.A(n_1953),
.B(n_1870),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1960),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1948),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1950),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1952),
.B(n_1971),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1960),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1971),
.B(n_1851),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1961),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1976),
.B(n_1837),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1961),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1945),
.B(n_1935),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1963),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1976),
.B(n_1837),
.Y(n_2019)
);

INVxp67_ASAP7_75t_L g2020 ( 
.A(n_1956),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1943),
.B(n_1932),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1963),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1964),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1955),
.B(n_1814),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_1984),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1980),
.A2(n_1925),
.B1(n_1885),
.B2(n_1870),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1950),
.Y(n_2027)
);

INVx4_ASAP7_75t_L g2028 ( 
.A(n_1980),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1964),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1973),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1955),
.B(n_1814),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1994),
.B(n_1949),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1973),
.Y(n_2033)
);

INVx1_ASAP7_75t_SL g2034 ( 
.A(n_1965),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1946),
.B(n_1848),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1974),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1994),
.B(n_1920),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1946),
.B(n_1848),
.Y(n_2038)
);

INVx1_ASAP7_75t_SL g2039 ( 
.A(n_1970),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1949),
.B(n_1920),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1977),
.B(n_1848),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1956),
.B(n_1814),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1981),
.B(n_1815),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1951),
.B(n_1891),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1974),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1980),
.A2(n_1913),
.B(n_1903),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1981),
.B(n_1815),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1950),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1985),
.B(n_1959),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1951),
.B(n_1815),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1999),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2001),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_2004),
.B(n_1912),
.C(n_1944),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2000),
.B(n_1982),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2001),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2005),
.B(n_1995),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1999),
.Y(n_2057)
);

NAND4xp25_ASAP7_75t_L g2058 ( 
.A(n_2046),
.B(n_1892),
.C(n_2026),
.D(n_1889),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1999),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_2028),
.B(n_1995),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2006),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2006),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2008),
.Y(n_2063)
);

INVx4_ASAP7_75t_L g2064 ( 
.A(n_2025),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_2028),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2003),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2049),
.B(n_1992),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2020),
.B(n_1982),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_2034),
.Y(n_2069)
);

INVx4_ASAP7_75t_L g2070 ( 
.A(n_2025),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2008),
.Y(n_2071)
);

NOR3xp33_ASAP7_75t_SL g2072 ( 
.A(n_2002),
.B(n_1941),
.C(n_1906),
.Y(n_2072)
);

AOI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_2002),
.A2(n_1958),
.B1(n_1954),
.B2(n_1953),
.C(n_1968),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2003),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2012),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2034),
.B(n_1988),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2003),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2009),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2009),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2039),
.B(n_1988),
.Y(n_2080)
);

OAI31xp33_ASAP7_75t_L g2081 ( 
.A1(n_2005),
.A2(n_1900),
.A3(n_1904),
.B(n_1905),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2012),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2039),
.B(n_2042),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2014),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2024),
.B(n_1989),
.Y(n_2085)
);

AND2x4_ASAP7_75t_SL g2086 ( 
.A(n_2028),
.B(n_1995),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2014),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2016),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2032),
.B(n_1995),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2032),
.B(n_1972),
.Y(n_2090)
);

AOI221xp5_ASAP7_75t_L g2091 ( 
.A1(n_2017),
.A2(n_1958),
.B1(n_1954),
.B2(n_1968),
.C(n_1959),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_2028),
.Y(n_2092)
);

INVxp33_ASAP7_75t_L g2093 ( 
.A(n_2031),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2049),
.B(n_2017),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2043),
.B(n_1989),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2007),
.B(n_1972),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_1998),
.B(n_1992),
.Y(n_2097)
);

INVxp67_ASAP7_75t_SL g2098 ( 
.A(n_2007),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_1998),
.B(n_1997),
.Y(n_2099)
);

OAI32xp33_ASAP7_75t_L g2100 ( 
.A1(n_2053),
.A2(n_1968),
.A3(n_1997),
.B1(n_2025),
.B2(n_2041),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2056),
.B(n_2013),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2069),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2072),
.A2(n_2026),
.B1(n_1894),
.B2(n_2047),
.Y(n_2103)
);

OAI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_2058),
.A2(n_1899),
.B(n_1859),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_2058),
.A2(n_1979),
.B(n_1969),
.Y(n_2105)
);

OAI221xp5_ASAP7_75t_L g2106 ( 
.A1(n_2081),
.A2(n_1979),
.B1(n_2041),
.B2(n_2038),
.C(n_2035),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_2054),
.B(n_2050),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2052),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2081),
.B(n_2050),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2076),
.B(n_2044),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2052),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_2080),
.B(n_1909),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2051),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2064),
.B(n_2044),
.Y(n_2114)
);

AOI21xp33_ASAP7_75t_L g2115 ( 
.A1(n_2092),
.A2(n_2038),
.B(n_2035),
.Y(n_2115)
);

OAI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_2073),
.A2(n_1966),
.B(n_1962),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2055),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2064),
.B(n_2015),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2055),
.Y(n_2119)
);

NOR3xp33_ASAP7_75t_L g2120 ( 
.A(n_2064),
.B(n_1968),
.C(n_2009),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2061),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_2093),
.B(n_1984),
.Y(n_2122)
);

OAI22xp5_ASAP7_75t_SL g2123 ( 
.A1(n_2092),
.A2(n_1822),
.B1(n_1820),
.B2(n_1984),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2051),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2061),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2056),
.B(n_2086),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2064),
.B(n_2015),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2070),
.B(n_2019),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2051),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2070),
.B(n_2019),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2086),
.B(n_2013),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2094),
.A2(n_1824),
.B1(n_1810),
.B2(n_1860),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2062),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2086),
.B(n_2037),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2094),
.A2(n_2098),
.B1(n_2060),
.B2(n_2083),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2060),
.A2(n_1824),
.B1(n_1810),
.B2(n_1860),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2062),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2063),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2126),
.B(n_2065),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2126),
.Y(n_2140)
);

OAI321xp33_ASAP7_75t_L g2141 ( 
.A1(n_2135),
.A2(n_2091),
.A3(n_2096),
.B1(n_2068),
.B2(n_2097),
.C(n_2099),
.Y(n_2141)
);

XOR2x2_ASAP7_75t_L g2142 ( 
.A(n_2103),
.B(n_2070),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2134),
.B(n_2065),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2102),
.B(n_2068),
.Y(n_2144)
);

NAND2x1_ASAP7_75t_L g2145 ( 
.A(n_2134),
.B(n_2065),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2108),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_2131),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2108),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2131),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2104),
.B(n_2070),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2101),
.B(n_2065),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2110),
.B(n_2067),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2109),
.A2(n_2060),
.B1(n_2090),
.B2(n_2096),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2111),
.Y(n_2154)
);

AOI221xp5_ASAP7_75t_L g2155 ( 
.A1(n_2100),
.A2(n_2060),
.B1(n_2071),
.B2(n_2084),
.C(n_2075),
.Y(n_2155)
);

OAI222xp33_ASAP7_75t_L g2156 ( 
.A1(n_2106),
.A2(n_2105),
.B1(n_2114),
.B2(n_2128),
.C1(n_2127),
.C2(n_2118),
.Y(n_2156)
);

OAI22xp5_ASAP7_75t_SL g2157 ( 
.A1(n_2123),
.A2(n_2116),
.B1(n_2122),
.B2(n_2130),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2111),
.Y(n_2158)
);

OAI31xp33_ASAP7_75t_L g2159 ( 
.A1(n_2112),
.A2(n_2115),
.A3(n_2136),
.B(n_2132),
.Y(n_2159)
);

AOI221xp5_ASAP7_75t_L g2160 ( 
.A1(n_2100),
.A2(n_2087),
.B1(n_2082),
.B2(n_2075),
.C(n_2084),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_2107),
.A2(n_2088),
.B(n_2082),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2117),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2117),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2121),
.B(n_2067),
.Y(n_2164)
);

OAI321xp33_ASAP7_75t_L g2165 ( 
.A1(n_2101),
.A2(n_2138),
.A3(n_2137),
.B1(n_2119),
.B2(n_2125),
.C(n_2133),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_2119),
.Y(n_2166)
);

O2A1O1Ixp33_ASAP7_75t_L g2167 ( 
.A1(n_2120),
.A2(n_2063),
.B(n_2071),
.C(n_2087),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2146),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2148),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2140),
.B(n_2090),
.Y(n_2170)
);

CKINVDCx20_ASAP7_75t_R g2171 ( 
.A(n_2142),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2139),
.B(n_2089),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2139),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2150),
.B(n_2125),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2154),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2158),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2162),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_2156),
.B(n_2141),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2163),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_2165),
.B(n_2144),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2144),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2143),
.B(n_2089),
.Y(n_2182)
);

NAND3xp33_ASAP7_75t_L g2183 ( 
.A(n_2155),
.B(n_2138),
.C(n_2137),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2164),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2149),
.B(n_2095),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2143),
.B(n_2113),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2164),
.Y(n_2187)
);

NAND2x1_ASAP7_75t_L g2188 ( 
.A(n_2147),
.B(n_2113),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2166),
.Y(n_2189)
);

NOR3xp33_ASAP7_75t_SL g2190 ( 
.A(n_2157),
.B(n_2088),
.C(n_2085),
.Y(n_2190)
);

AOI31xp33_ASAP7_75t_L g2191 ( 
.A1(n_2153),
.A2(n_2129),
.A3(n_2124),
.B(n_2097),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2173),
.B(n_2182),
.Y(n_2192)
);

XOR2x2_ASAP7_75t_L g2193 ( 
.A(n_2178),
.B(n_2142),
.Y(n_2193)
);

AND4x1_ASAP7_75t_L g2194 ( 
.A(n_2190),
.B(n_2159),
.C(n_2161),
.D(n_2167),
.Y(n_2194)
);

OR3x1_ASAP7_75t_L g2195 ( 
.A(n_2178),
.B(n_2180),
.C(n_2174),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2184),
.Y(n_2196)
);

NAND3xp33_ASAP7_75t_L g2197 ( 
.A(n_2180),
.B(n_2160),
.C(n_2149),
.Y(n_2197)
);

NAND2xp33_ASAP7_75t_SL g2198 ( 
.A(n_2171),
.B(n_2145),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2187),
.B(n_2147),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_2171),
.B(n_2152),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2181),
.B(n_2147),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2186),
.Y(n_2202)
);

NAND4xp75_ASAP7_75t_L g2203 ( 
.A(n_2189),
.B(n_2151),
.C(n_2145),
.D(n_2124),
.Y(n_2203)
);

INVxp67_ASAP7_75t_SL g2204 ( 
.A(n_2188),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_2183),
.B(n_2151),
.C(n_2152),
.Y(n_2205)
);

O2A1O1Ixp33_ASAP7_75t_L g2206 ( 
.A1(n_2191),
.A2(n_2129),
.B(n_2099),
.C(n_2079),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2174),
.B(n_2011),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2200),
.B(n_2186),
.Y(n_2208)
);

OAI22xp33_ASAP7_75t_SL g2209 ( 
.A1(n_2204),
.A2(n_2201),
.B1(n_2196),
.B2(n_2199),
.Y(n_2209)
);

NAND4xp25_ASAP7_75t_L g2210 ( 
.A(n_2197),
.B(n_2170),
.C(n_2168),
.D(n_2179),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2192),
.B(n_2182),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2203),
.Y(n_2212)
);

OAI211xp5_ASAP7_75t_SL g2213 ( 
.A1(n_2201),
.A2(n_2177),
.B(n_2176),
.C(n_2175),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2202),
.B(n_2172),
.Y(n_2214)
);

OAI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2195),
.A2(n_2185),
.B1(n_2169),
.B2(n_2037),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2205),
.B(n_2011),
.Y(n_2216)
);

NAND5xp2_ASAP7_75t_L g2217 ( 
.A(n_2206),
.B(n_2040),
.C(n_1908),
.D(n_1860),
.E(n_1975),
.Y(n_2217)
);

AOI222xp33_ASAP7_75t_L g2218 ( 
.A1(n_2193),
.A2(n_2079),
.B1(n_2057),
.B2(n_2059),
.C1(n_2066),
.C2(n_2078),
.Y(n_2218)
);

AOI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2198),
.A2(n_2207),
.B(n_2194),
.Y(n_2219)
);

A2O1A1Ixp33_ASAP7_75t_L g2220 ( 
.A1(n_2207),
.A2(n_1993),
.B(n_1957),
.C(n_1967),
.Y(n_2220)
);

AOI221xp5_ASAP7_75t_L g2221 ( 
.A1(n_2197),
.A2(n_2079),
.B1(n_2057),
.B2(n_2078),
.C(n_2059),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2212),
.B(n_2040),
.Y(n_2222)
);

NOR3xp33_ASAP7_75t_L g2223 ( 
.A(n_2208),
.B(n_2219),
.C(n_2209),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2215),
.A2(n_1993),
.B1(n_1991),
.B2(n_1983),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2211),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2214),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_2216),
.Y(n_2227)
);

NAND4xp75_ASAP7_75t_L g2228 ( 
.A(n_2221),
.B(n_2078),
.C(n_2077),
.D(n_2074),
.Y(n_2228)
);

HB1xp67_ASAP7_75t_L g2229 ( 
.A(n_2210),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2213),
.Y(n_2230)
);

BUFx2_ASAP7_75t_L g2231 ( 
.A(n_2227),
.Y(n_2231)
);

NAND4xp75_ASAP7_75t_L g2232 ( 
.A(n_2230),
.B(n_2218),
.C(n_2217),
.D(n_2220),
.Y(n_2232)
);

OAI211xp5_ASAP7_75t_SL g2233 ( 
.A1(n_2223),
.A2(n_2077),
.B(n_2074),
.C(n_2057),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2228),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2222),
.B(n_2226),
.Y(n_2235)
);

NOR2x1_ASAP7_75t_L g2236 ( 
.A(n_2225),
.B(n_2059),
.Y(n_2236)
);

AOI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2229),
.A2(n_2077),
.B1(n_2066),
.B2(n_2074),
.C(n_2027),
.Y(n_2237)
);

OAI311xp33_ASAP7_75t_L g2238 ( 
.A1(n_2224),
.A2(n_2021),
.A3(n_1990),
.B1(n_1996),
.C1(n_1985),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_2231),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2235),
.Y(n_2240)
);

OAI311xp33_ASAP7_75t_L g2241 ( 
.A1(n_2237),
.A2(n_2224),
.A3(n_2021),
.B1(n_1990),
.C1(n_1996),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2234),
.B(n_2066),
.Y(n_2242)
);

AND3x2_ASAP7_75t_L g2243 ( 
.A(n_2233),
.B(n_2022),
.C(n_2018),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2232),
.B(n_2016),
.Y(n_2244)
);

OAI221xp5_ASAP7_75t_L g2245 ( 
.A1(n_2236),
.A2(n_2048),
.B1(n_2010),
.B2(n_2027),
.C(n_1957),
.Y(n_2245)
);

OAI322xp33_ASAP7_75t_L g2246 ( 
.A1(n_2238),
.A2(n_2048),
.A3(n_2010),
.B1(n_2027),
.B2(n_1967),
.C1(n_1957),
.C2(n_2030),
.Y(n_2246)
);

AOI21xp33_ASAP7_75t_L g2247 ( 
.A1(n_2239),
.A2(n_2048),
.B(n_2010),
.Y(n_2247)
);

INVx1_ASAP7_75t_SL g2248 ( 
.A(n_2240),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2242),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2244),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2250),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2248),
.A2(n_2243),
.B1(n_2245),
.B2(n_2241),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2252),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2251),
.Y(n_2254)
);

NOR2xp67_ASAP7_75t_L g2255 ( 
.A(n_2254),
.B(n_2249),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2253),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2253),
.A2(n_2247),
.B1(n_2246),
.B2(n_2033),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2256),
.Y(n_2258)
);

AOI21xp33_ASAP7_75t_SL g2259 ( 
.A1(n_2257),
.A2(n_2045),
.B(n_2018),
.Y(n_2259)
);

OAI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2258),
.A2(n_2255),
.B1(n_2033),
.B2(n_2045),
.Y(n_2260)
);

AOI21xp33_ASAP7_75t_L g2261 ( 
.A1(n_2259),
.A2(n_2036),
.B(n_2030),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_2260),
.A2(n_2036),
.B1(n_2029),
.B2(n_2023),
.Y(n_2262)
);

OAI221xp5_ASAP7_75t_R g2263 ( 
.A1(n_2262),
.A2(n_2261),
.B1(n_2029),
.B2(n_2023),
.C(n_2022),
.Y(n_2263)
);

AOI211xp5_ASAP7_75t_L g2264 ( 
.A1(n_2263),
.A2(n_1910),
.B(n_1967),
.C(n_1991),
.Y(n_2264)
);


endmodule