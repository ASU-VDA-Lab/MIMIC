module fake_jpeg_17983_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.C(n_34),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_45),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_22),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_36),
.B1(n_52),
.B2(n_41),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_75),
.B1(n_76),
.B2(n_80),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_74),
.Y(n_105)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_21),
.B1(n_17),
.B2(n_36),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_32),
.B1(n_37),
.B2(n_35),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_21),
.B1(n_28),
.B2(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_21),
.B1(n_28),
.B2(n_27),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_46),
.B(n_44),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_88),
.B(n_25),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_89),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_44),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_45),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_82),
.C(n_73),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_106),
.B1(n_110),
.B2(n_18),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_31),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_37),
.B1(n_32),
.B2(n_34),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_78),
.B1(n_55),
.B2(n_53),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_49),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_0),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_31),
.B1(n_25),
.B2(n_18),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_65),
.A2(n_22),
.B1(n_15),
.B2(n_49),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_23),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_134),
.B1(n_107),
.B2(n_92),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_123),
.C(n_126),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_119),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_131),
.CI(n_122),
.CON(n_141),
.SN(n_141)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_131),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_61),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_107),
.B1(n_93),
.B2(n_96),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_78),
.C(n_24),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_15),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_109),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_83),
.B(n_74),
.C(n_72),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_58),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_54),
.B1(n_58),
.B2(n_35),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_112),
.B1(n_128),
.B2(n_95),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_146),
.B1(n_148),
.B2(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_107),
.B1(n_86),
.B2(n_93),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_158),
.B1(n_126),
.B2(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_98),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_156),
.C(n_115),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_115),
.B(n_134),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_98),
.B1(n_112),
.B2(n_109),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_100),
.B(n_104),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_25),
.B(n_20),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_24),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_168),
.A2(n_175),
.B1(n_186),
.B2(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_130),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_171),
.C(n_174),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_125),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_185),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_173),
.B(n_0),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_92),
.B1(n_94),
.B2(n_91),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_54),
.C(n_79),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_179),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_97),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_196),
.B(n_137),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_54),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_182),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_70),
.C(n_58),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_91),
.B1(n_58),
.B2(n_30),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_91),
.Y(n_191)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_144),
.B(n_137),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_26),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_137),
.Y(n_216)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_26),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_148),
.A2(n_30),
.B1(n_29),
.B2(n_20),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_159),
.CI(n_155),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_202),
.B(n_213),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_210),
.C(n_219),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_160),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_142),
.B1(n_158),
.B2(n_140),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_220),
.B(n_227),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_224),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_141),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_141),
.B(n_151),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_151),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_222),
.C(n_189),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_26),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_173),
.A2(n_26),
.B(n_9),
.Y(n_225)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_200),
.B1(n_13),
.B2(n_14),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_180),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_232),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_184),
.B1(n_178),
.B2(n_198),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_190),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_232),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_198),
.B1(n_183),
.B2(n_186),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_9),
.C(n_14),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_209),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_1),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_1),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_221),
.C(n_201),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_262),
.C(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_254),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_208),
.B(n_210),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_243),
.B(n_246),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_244),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_202),
.B1(n_204),
.B2(n_206),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_248),
.B1(n_245),
.B2(n_231),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_201),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_1),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_206),
.C(n_209),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_216),
.C(n_30),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_275),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_235),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_281),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_265),
.B(n_230),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_274),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_240),
.C(n_248),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_258),
.B1(n_259),
.B2(n_255),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_277),
.B1(n_2),
.B2(n_3),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_229),
.B1(n_237),
.B2(n_3),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_257),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_12),
.B(n_11),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_254),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_286),
.B1(n_294),
.B2(n_269),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_291),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_250),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_277),
.Y(n_296)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_2),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_262),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_2),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_268),
.A2(n_266),
.B1(n_251),
.B2(n_10),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_269),
.C(n_267),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_301),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_299),
.Y(n_312)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_281),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_29),
.B1(n_20),
.B2(n_11),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_29),
.B1(n_5),
.B2(n_6),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_3),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_SL g304 ( 
.A(n_284),
.B(n_4),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_304),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_296),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_311),
.B1(n_7),
.B2(n_4),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_289),
.B1(n_288),
.B2(n_292),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_4),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_297),
.B(n_288),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_312),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_318),
.C(n_313),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_312),
.B(n_305),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_316),
.C(n_6),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_6),
.B(n_7),
.Y(n_325)
);


endmodule