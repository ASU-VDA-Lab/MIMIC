module fake_aes_12094_n_660 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_660);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_660;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_74), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_3), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_39), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_2), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_48), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_71), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_4), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_46), .B(n_24), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_16), .Y(n_87) );
BUFx2_ASAP7_75t_SL g88 ( .A(n_20), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_43), .Y(n_89) );
INVx2_ASAP7_75t_SL g90 ( .A(n_64), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_22), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_66), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_67), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_63), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_61), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_1), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_16), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_37), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_75), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_9), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_30), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_38), .B(n_28), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g104 ( .A(n_15), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_47), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_29), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_7), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_18), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_11), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_68), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_60), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_31), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_32), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_23), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_1), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_11), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_44), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_42), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_107), .Y(n_122) );
OR2x2_ASAP7_75t_L g123 ( .A(n_82), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_107), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_89), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_90), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_104), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_89), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_94), .B(n_2), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_121), .B(n_4), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_113), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_90), .B(n_5), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_113), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_113), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_79), .B(n_98), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_108), .B(n_5), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_105), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_80), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_82), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_95), .B(n_8), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_115), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_78), .B(n_9), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_96), .B(n_10), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_99), .B(n_10), .Y(n_156) );
NAND2xp33_ASAP7_75t_SL g157 ( .A(n_84), .B(n_12), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
INVx1_ASAP7_75t_SL g159 ( .A(n_149), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_124), .B(n_120), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_132), .B(n_101), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_124), .B(n_83), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_152), .A2(n_120), .B(n_116), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_132), .B(n_87), .Y(n_168) );
INVx1_ASAP7_75t_SL g169 ( .A(n_145), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_122), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_127), .B(n_101), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_127), .B(n_111), .Y(n_172) );
INVx11_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_122), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_129), .B(n_102), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_122), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_133), .B(n_118), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_129), .B(n_102), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_122), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_139), .B(n_87), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_123), .B(n_119), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_139), .B(n_83), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_145), .B(n_109), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_140), .B(n_109), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_125), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_125), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_125), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
AND2x6_ASAP7_75t_L g195 ( .A(n_140), .B(n_119), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_126), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_134), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_126), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_141), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_134), .Y(n_201) );
OR2x6_ASAP7_75t_L g202 ( .A(n_123), .B(n_88), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_180), .B(n_142), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_187), .Y(n_208) );
AND2x6_ASAP7_75t_L g209 ( .A(n_185), .B(n_141), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_195), .A2(n_158), .B1(n_144), .B2(n_146), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_200), .B(n_144), .Y(n_211) );
NAND2xp33_ASAP7_75t_L g212 ( .A(n_195), .B(n_158), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_159), .B(n_135), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g214 ( .A1(n_159), .A2(n_97), .B1(n_147), .B2(n_148), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_180), .B(n_150), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
NAND3xp33_ASAP7_75t_SL g217 ( .A(n_169), .B(n_106), .C(n_100), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_200), .B(n_146), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_182), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_202), .A2(n_150), .B1(n_153), .B2(n_128), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_184), .B(n_153), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_182), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_162), .B(n_157), .Y(n_223) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_169), .B(n_100), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_175), .B(n_154), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_202), .B(n_85), .Y(n_226) );
NOR2x1p5_ASAP7_75t_L g227 ( .A(n_183), .B(n_85), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_202), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_182), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_175), .B(n_155), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_202), .B(n_110), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_164), .B(n_156), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_187), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_172), .B(n_131), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_176), .B(n_137), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_172), .B(n_131), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_163), .B(n_137), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_183), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_182), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g240 ( .A1(n_202), .A2(n_117), .B1(n_110), .B2(n_118), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_163), .B(n_112), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_168), .B(n_91), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_168), .B(n_117), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_186), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_179), .B(n_88), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_186), .Y(n_247) );
BUFx4f_ASAP7_75t_SL g248 ( .A(n_195), .Y(n_248) );
CKINVDCx11_ASAP7_75t_R g249 ( .A(n_173), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_187), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_186), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_179), .B(n_134), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_185), .B(n_86), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_166), .A2(n_103), .B1(n_138), .B2(n_136), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_192), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_196), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_238), .A2(n_160), .B(n_196), .C(n_199), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_249), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_238), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_223), .B(n_173), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_207), .B(n_166), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_207), .B(n_166), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_257), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_209), .B(n_166), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_225), .B(n_192), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_209), .B(n_195), .Y(n_267) );
NOR2x1_ASAP7_75t_L g268 ( .A(n_217), .B(n_160), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_240), .A2(n_199), .B(n_181), .C(n_188), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_211), .A2(n_188), .B(n_189), .Y(n_270) );
AND2x6_ASAP7_75t_L g271 ( .A(n_226), .B(n_181), .Y(n_271) );
BUFx12f_ASAP7_75t_L g272 ( .A(n_226), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_209), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_246), .A2(n_189), .B(n_174), .C(n_170), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
INVx4_ASAP7_75t_L g277 ( .A(n_209), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_228), .Y(n_278) );
BUFx5_ASAP7_75t_L g279 ( .A(n_204), .Y(n_279) );
OAI22x1_ASAP7_75t_L g280 ( .A1(n_227), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_219), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_219), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_205), .Y(n_283) );
NOR2x1_ASAP7_75t_L g284 ( .A(n_240), .B(n_174), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_231), .A2(n_192), .B1(n_170), .B2(n_177), .Y(n_285) );
CKINVDCx11_ASAP7_75t_R g286 ( .A(n_231), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_248), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_248), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_208), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_211), .A2(n_177), .B(n_192), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_206), .Y(n_291) );
AO21x1_ASAP7_75t_L g292 ( .A1(n_255), .A2(n_167), .B(n_161), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_215), .B(n_195), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_214), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_233), .Y(n_295) );
NOR2xp67_ASAP7_75t_SL g296 ( .A(n_224), .B(n_195), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_218), .A2(n_165), .B(n_201), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_246), .A2(n_195), .B1(n_201), .B2(n_198), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_230), .B(n_201), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_218), .A2(n_165), .B(n_201), .Y(n_301) );
BUFx12f_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_250), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_216), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_277), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_262), .A2(n_220), .B1(n_210), .B2(n_251), .Y(n_307) );
NOR2x1_ASAP7_75t_SL g308 ( .A(n_277), .B(n_221), .Y(n_308) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_292), .A2(n_244), .B(n_252), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_265), .A2(n_210), .B(n_213), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_262), .A2(n_237), .B(n_247), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_286), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_265), .A2(n_229), .B(n_245), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_260), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_276), .B(n_239), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_274), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_283), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_272), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_291), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_279), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_263), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_271), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_294), .A2(n_232), .B1(n_222), .B2(n_195), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_279), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_289), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_263), .A2(n_242), .B(n_241), .C(n_254), .Y(n_329) );
AO21x1_ASAP7_75t_L g330 ( .A1(n_258), .A2(n_237), .B(n_232), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_278), .A2(n_236), .B1(n_234), .B2(n_235), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_296), .B(n_235), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_268), .A2(n_203), .B(n_194), .Y(n_334) );
NOR2x1_ASAP7_75t_SL g335 ( .A(n_267), .B(n_212), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_270), .A2(n_203), .B(n_178), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_275), .A2(n_198), .B(n_165), .C(n_138), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g338 ( .A(n_288), .B(n_165), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_329), .A2(n_293), .B(n_269), .C(n_284), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_324), .A2(n_317), .B1(n_314), .B2(n_325), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_329), .A2(n_293), .B(n_266), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_324), .A2(n_273), .B1(n_267), .B2(n_264), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_319), .B(n_261), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_332), .A2(n_302), .B1(n_280), .B2(n_305), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_319), .Y(n_346) );
AOI222xp33_ASAP7_75t_L g347 ( .A1(n_314), .A2(n_300), .B1(n_259), .B2(n_282), .C1(n_281), .C2(n_271), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
BUFx4f_ASAP7_75t_SL g349 ( .A(n_315), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_337), .A2(n_270), .B(n_290), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_321), .Y(n_352) );
OAI21xp5_ASAP7_75t_SL g353 ( .A1(n_326), .A2(n_298), .B(n_287), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_313), .A2(n_279), .B1(n_281), .B2(n_271), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_315), .A2(n_285), .B1(n_303), .B2(n_288), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_303), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g357 ( .A1(n_313), .A2(n_290), .B1(n_299), .B2(n_301), .C(n_297), .Y(n_357) );
AOI222xp33_ASAP7_75t_L g358 ( .A1(n_322), .A2(n_271), .B1(n_299), .B2(n_295), .C1(n_304), .C2(n_289), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_289), .Y(n_359) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_316), .A2(n_301), .B(n_297), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_325), .A2(n_198), .B1(n_151), .B2(n_138), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_316), .Y(n_362) );
BUFx10_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_316), .B(n_13), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_325), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_359), .B(n_311), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_362), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_348), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_360), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_364), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_359), .B(n_311), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_346), .B(n_311), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_350), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_360), .Y(n_374) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_364), .B(n_309), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_360), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_356), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_356), .B(n_309), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_344), .B(n_318), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_345), .B(n_318), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_363), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_352), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_347), .B(n_318), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_363), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_363), .B(n_309), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_357), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_365), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_309), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_349), .A2(n_307), .B1(n_306), .B2(n_331), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_339), .B(n_323), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_352), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_339), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_343), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_341), .B(n_323), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_342), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_381), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_378), .B(n_310), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_367), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_381), .B(n_310), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_366), .B(n_334), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_382), .Y(n_403) );
AO31x2_ASAP7_75t_L g404 ( .A1(n_386), .A2(n_330), .A3(n_351), .B(n_307), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_370), .B(n_330), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_366), .B(n_334), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_367), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_384), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_387), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_392), .B(n_353), .Y(n_410) );
AOI322xp5_ASAP7_75t_L g411 ( .A1(n_368), .A2(n_354), .A3(n_15), .B1(n_14), .B2(n_318), .C1(n_306), .C2(n_312), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_369), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_370), .B(n_334), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_369), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_369), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_380), .A2(n_358), .B1(n_355), .B2(n_333), .C(n_361), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
OAI321xp33_ASAP7_75t_L g418 ( .A1(n_389), .A2(n_393), .A3(n_383), .B1(n_388), .B2(n_386), .C(n_385), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_371), .B(n_336), .Y(n_419) );
AO21x2_ASAP7_75t_L g420 ( .A1(n_386), .A2(n_336), .B(n_308), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_372), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_378), .B(n_323), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
OR2x6_ASAP7_75t_L g424 ( .A(n_396), .B(n_310), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_371), .B(n_312), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_384), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_374), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_372), .B(n_312), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_368), .B(n_395), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_377), .B(n_308), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_385), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_374), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_395), .B(n_327), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_379), .A2(n_333), .B1(n_338), .B2(n_328), .C(n_327), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_377), .A2(n_327), .B1(n_333), .B2(n_328), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_376), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_394), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_376), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_376), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_399), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_421), .B(n_375), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_421), .B(n_375), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_399), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_410), .B(n_394), .C(n_393), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_400), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_429), .B(n_391), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_412), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_400), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_403), .B(n_390), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_419), .B(n_391), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_432), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_429), .B(n_388), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_387), .Y(n_454) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_409), .B(n_387), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_417), .B(n_390), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_422), .B(n_396), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_398), .B(n_396), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_432), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_425), .B(n_151), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_411), .B(n_136), .C(n_138), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_437), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_437), .B(n_328), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_407), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_425), .B(n_151), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_419), .B(n_336), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_428), .B(n_151), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_428), .B(n_151), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_408), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_419), .B(n_151), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_407), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_414), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_408), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_419), .B(n_138), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_407), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_402), .B(n_406), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_422), .B(n_138), .Y(n_477) );
NOR2xp67_ASAP7_75t_L g478 ( .A(n_426), .B(n_328), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_402), .B(n_17), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_405), .B(n_335), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_414), .Y(n_481) );
NOR2xp67_ASAP7_75t_L g482 ( .A(n_426), .B(n_19), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_402), .B(n_21), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_415), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_397), .B(n_26), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_402), .B(n_27), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_415), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_406), .B(n_33), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_406), .B(n_34), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_409), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_411), .A2(n_338), .B1(n_193), .B2(n_161), .C(n_167), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_406), .B(n_35), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_423), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_431), .B(n_36), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_433), .B(n_335), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_431), .A2(n_338), .B1(n_45), .B2(n_49), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_447), .B(n_438), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_462), .B(n_438), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_453), .B(n_405), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_440), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_469), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_462), .B(n_431), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_440), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_450), .B(n_397), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_456), .B(n_397), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_453), .B(n_431), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_454), .B(n_439), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_454), .B(n_439), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_441), .B(n_433), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_441), .B(n_430), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_473), .B(n_423), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_455), .Y(n_513) );
OAI21xp33_ASAP7_75t_SL g514 ( .A1(n_455), .A2(n_435), .B(n_413), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_451), .B(n_431), .Y(n_515) );
OAI21xp33_ASAP7_75t_L g516 ( .A1(n_461), .A2(n_401), .B(n_435), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_451), .B(n_431), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_442), .B(n_413), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_490), .B(n_427), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_451), .B(n_401), .Y(n_520) );
OR2x6_ASAP7_75t_L g521 ( .A(n_482), .B(n_401), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_490), .B(n_436), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_444), .Y(n_523) );
AOI31xp33_ASAP7_75t_L g524 ( .A1(n_461), .A2(n_436), .A3(n_427), .B(n_416), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_442), .B(n_404), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_446), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_446), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_451), .B(n_424), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_457), .B(n_424), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_476), .B(n_424), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_482), .A2(n_418), .B(n_434), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_485), .A2(n_424), .B(n_404), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_457), .B(n_424), .Y(n_533) );
NOR2x1p5_ASAP7_75t_L g534 ( .A(n_476), .B(n_404), .Y(n_534) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_455), .A2(n_193), .B(n_167), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_445), .B(n_41), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_460), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_449), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_458), .B(n_404), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_458), .B(n_404), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_467), .B(n_420), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_443), .Y(n_542) );
NAND2x1_ASAP7_75t_L g543 ( .A(n_478), .B(n_476), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_449), .B(n_420), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_476), .B(n_420), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_452), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_452), .B(n_50), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_467), .B(n_51), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_470), .B(n_474), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_468), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_494), .B(n_52), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_470), .B(n_53), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_479), .B(n_54), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_499), .B(n_468), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_500), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_501), .B(n_474), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_507), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_524), .A2(n_478), .B1(n_479), .B2(n_488), .Y(n_559) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_524), .B(n_494), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_506), .B(n_466), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_537), .B(n_466), .Y(n_562) );
NOR2xp33_ASAP7_75t_SL g563 ( .A(n_516), .B(n_483), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_497), .B(n_460), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_503), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_516), .A2(n_496), .B(n_492), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_544), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_531), .A2(n_489), .B(n_483), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_514), .B(n_464), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_511), .Y(n_570) );
AO22x2_ASAP7_75t_L g571 ( .A1(n_513), .A2(n_459), .B1(n_471), .B2(n_475), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_543), .A2(n_486), .B(n_492), .C(n_488), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_531), .A2(n_489), .B(n_486), .Y(n_573) );
OAI32xp33_ASAP7_75t_L g574 ( .A1(n_551), .A2(n_459), .A3(n_464), .B1(n_477), .B2(n_480), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_521), .A2(n_466), .B1(n_495), .B2(n_464), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_523), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_512), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_532), .A2(n_480), .B1(n_463), .B2(n_475), .C(n_471), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_544), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_508), .B(n_481), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_526), .B(n_527), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_SL g582 ( .A1(n_504), .A2(n_481), .B(n_477), .C(n_464), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_538), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_535), .A2(n_466), .B(n_448), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_546), .B(n_465), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_518), .B(n_493), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_522), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_549), .Y(n_588) );
OAI31xp33_ASAP7_75t_L g589 ( .A1(n_534), .A2(n_465), .A3(n_491), .B(n_487), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_532), .A2(n_493), .B1(n_487), .B2(n_484), .C(n_472), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_498), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_540), .B(n_493), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_530), .B(n_487), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_550), .B(n_484), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_536), .A2(n_484), .B1(n_472), .B2(n_448), .C(n_443), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_573), .A2(n_505), .B1(n_545), .B2(n_528), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_555), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_581), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_588), .B(n_520), .Y(n_599) );
OAI222xp33_ASAP7_75t_L g600 ( .A1(n_560), .A2(n_521), .B1(n_539), .B2(n_529), .C1(n_533), .C2(n_525), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_567), .B(n_542), .Y(n_601) );
OAI221xp5_ASAP7_75t_SL g602 ( .A1(n_589), .A2(n_509), .B1(n_510), .B2(n_517), .C(n_515), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_556), .Y(n_603) );
XOR2x2_ASAP7_75t_L g604 ( .A(n_568), .B(n_551), .Y(n_604) );
XNOR2xp5_ASAP7_75t_L g605 ( .A(n_558), .B(n_552), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_561), .B(n_502), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_563), .B(n_535), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_555), .Y(n_608) );
OAI322xp33_ASAP7_75t_SL g609 ( .A1(n_569), .A2(n_578), .A3(n_590), .B1(n_554), .B2(n_564), .C1(n_557), .C2(n_592), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_580), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_565), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_559), .A2(n_553), .B1(n_541), .B2(n_521), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_566), .A2(n_547), .B1(n_548), .B2(n_472), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_570), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_569), .A2(n_547), .B(n_448), .C(n_443), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_572), .B(n_191), .Y(n_616) );
OAI322xp33_ASAP7_75t_L g617 ( .A1(n_567), .A2(n_161), .A3(n_178), .B1(n_194), .B2(n_193), .C1(n_203), .C2(n_190), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_595), .B(n_194), .C(n_178), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_562), .A2(n_197), .B1(n_191), .B2(n_190), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_577), .B(n_55), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_579), .B(n_56), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_596), .A2(n_575), .B1(n_571), .B2(n_579), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_597), .B(n_594), .Y(n_623) );
AOI322xp5_ASAP7_75t_L g624 ( .A1(n_613), .A2(n_594), .A3(n_587), .B1(n_593), .B2(n_591), .C1(n_583), .C2(n_576), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_604), .A2(n_571), .B1(n_585), .B2(n_582), .Y(n_625) );
OAI22xp33_ASAP7_75t_SL g626 ( .A1(n_602), .A2(n_584), .B1(n_586), .B2(n_571), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_603), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_612), .A2(n_584), .B1(n_574), .B2(n_197), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_608), .B(n_57), .Y(n_629) );
OAI21xp33_ASAP7_75t_SL g630 ( .A1(n_607), .A2(n_58), .B(n_59), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_615), .B(n_197), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_609), .A2(n_197), .B1(n_191), .B2(n_190), .C(n_198), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_610), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_SL g634 ( .A1(n_599), .A2(n_62), .B(n_65), .C(n_69), .Y(n_634) );
OAI21xp33_ASAP7_75t_SL g635 ( .A1(n_616), .A2(n_70), .B(n_73), .Y(n_635) );
AO22x2_ASAP7_75t_L g636 ( .A1(n_598), .A2(n_76), .B1(n_77), .B2(n_190), .Y(n_636) );
NOR4xp25_ASAP7_75t_L g637 ( .A(n_622), .B(n_600), .C(n_621), .D(n_611), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_624), .B(n_614), .Y(n_638) );
AOI21x1_ASAP7_75t_L g639 ( .A1(n_631), .A2(n_605), .B(n_621), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_626), .B(n_618), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_633), .B(n_606), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_627), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_625), .A2(n_601), .B1(n_617), .B2(n_620), .C(n_619), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_628), .A2(n_601), .B(n_191), .Y(n_644) );
AO22x2_ASAP7_75t_L g645 ( .A1(n_623), .A2(n_190), .B1(n_191), .B2(n_197), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_640), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_638), .Y(n_647) );
CKINVDCx16_ASAP7_75t_R g648 ( .A(n_637), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_642), .Y(n_649) );
NOR4xp25_ASAP7_75t_SL g650 ( .A(n_644), .B(n_634), .C(n_632), .D(n_630), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_648), .B(n_643), .Y(n_651) );
OR4x2_ASAP7_75t_L g652 ( .A(n_647), .B(n_639), .C(n_641), .D(n_645), .Y(n_652) );
NAND2x1p5_ASAP7_75t_L g653 ( .A(n_646), .B(n_629), .Y(n_653) );
OAI222xp33_ASAP7_75t_L g654 ( .A1(n_651), .A2(n_649), .B1(n_650), .B2(n_645), .C1(n_635), .C2(n_636), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_652), .Y(n_655) );
AO22x2_ASAP7_75t_SL g656 ( .A1(n_655), .A2(n_649), .B1(n_653), .B2(n_636), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_656), .B(n_655), .Y(n_657) );
OR2x6_ASAP7_75t_L g658 ( .A(n_657), .B(n_654), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_658), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_659), .A2(n_190), .B(n_191), .Y(n_660) );
endmodule