module fake_jpeg_18187_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_40),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_36),
.B1(n_31),
.B2(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_32),
.B1(n_26),
.B2(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_25),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_23),
.B(n_29),
.C(n_34),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_21),
.B(n_1),
.C(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_57),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_26),
.B1(n_18),
.B2(n_29),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_68),
.B1(n_3),
.B2(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_20),
.B1(n_17),
.B2(n_37),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_64),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_22),
.C(n_14),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_66),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_43),
.B1(n_49),
.B2(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_7),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_21),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_77),
.Y(n_86)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_7),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_68),
.B1(n_63),
.B2(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

XNOR2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_72),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_63),
.B(n_66),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_70),
.B(n_73),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_88),
.B(n_89),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_81),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_105),
.C(n_94),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_77),
.CI(n_82),
.CON(n_106),
.SN(n_106)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_106),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_74),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_108),
.B(n_113),
.Y(n_115)
);

AO221x1_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_93),
.B1(n_80),
.B2(n_71),
.C(n_78),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_105),
.C(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_74),
.B1(n_86),
.B2(n_95),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_98),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_117),
.B(n_118),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_119),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_92),
.C(n_86),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_106),
.B(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_71),
.B(n_11),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_124),
.Y(n_129)
);


endmodule