module fake_netlist_6_1092_n_145 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_61, n_39, n_63, n_60, n_59, n_32, n_4, n_66, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_20, n_50, n_49, n_7, n_30, n_64, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_62, n_31, n_65, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_145);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_61;
input n_39;
input n_63;
input n_60;
input n_59;
input n_32;
input n_4;
input n_66;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_64;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_62;
input n_31;
input n_65;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_145;

wire n_91;
wire n_119;
wire n_88;
wire n_98;
wire n_113;
wire n_73;
wire n_138;
wire n_68;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_132;
wire n_102;
wire n_87;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_75;
wire n_109;
wire n_122;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_112;
wire n_81;
wire n_76;
wire n_124;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_116;
wire n_117;
wire n_118;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_115;
wire n_69;
wire n_128;
wire n_79;

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_64),
.B1(n_46),
.B2(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_28),
.A2(n_58),
.B1(n_20),
.B2(n_29),
.Y(n_68)
);

OAI21x1_ASAP7_75t_L g69 ( 
.A1(n_30),
.A2(n_34),
.B(n_57),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_0),
.A2(n_63),
.B1(n_14),
.B2(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx8_ASAP7_75t_SL g74 ( 
.A(n_35),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_42),
.Y(n_75)
);

OAI21x1_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_33),
.B(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_52),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

OAI21x1_ASAP7_75t_L g84 ( 
.A1(n_22),
.A2(n_23),
.B(n_7),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_16),
.A2(n_15),
.B1(n_25),
.B2(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_26),
.A2(n_10),
.B(n_49),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_92),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_2),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AND2x4_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_6),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_11),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_13),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_32),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_37),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_87),
.B(n_85),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_76),
.B(n_84),
.Y(n_108)
);

AOI21x1_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_78),
.B(n_75),
.Y(n_109)
);

AO31x2_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_68),
.A3(n_90),
.B(n_69),
.Y(n_110)
);

AOI211x1_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_90),
.B(n_67),
.C(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_104),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_77),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_95),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

AO21x1_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_100),
.B(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

AOI222xp33_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_86),
.B1(n_112),
.B2(n_108),
.C1(n_110),
.C2(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_41),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_123),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_126),
.B(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_134),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_131),
.B(n_126),
.Y(n_139)
);

NAND4xp25_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_138),
.C(n_133),
.D(n_135),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_133),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_129),
.C(n_50),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_47),
.B(n_53),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_54),
.Y(n_144)
);

OR2x6_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_56),
.Y(n_145)
);


endmodule