module fake_jpeg_28458_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_15),
.B(n_34),
.C(n_29),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_2),
.Y(n_66)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_45),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_41),
.C(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_37),
.C(n_4),
.Y(n_75)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_71),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_46),
.B1(n_44),
.B2(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_44),
.B1(n_43),
.B2(n_39),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_76),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_81),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_4),
.B(n_5),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_5),
.B(n_7),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_91),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_59),
.C(n_58),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_17),
.C(n_18),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_9),
.C(n_10),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_95),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_28),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_100),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_20),
.C(n_22),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_96),
.C(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_108),
.C(n_96),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_86),
.C(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_111),
.B1(n_104),
.B2(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_105),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_104),
.B(n_93),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_23),
.B(n_25),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

XNOR2x2_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_109),
.Y(n_116)
);


endmodule