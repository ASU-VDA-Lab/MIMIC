module fake_jpeg_2727_n_515 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_455;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_378;
wire n_419;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_57),
.Y(n_146)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_64),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_68),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_78),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_15),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_87),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_22),
.B(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_83),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_34),
.B(n_13),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_35),
.B(n_13),
.Y(n_87)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_16),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_101),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_18),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_23),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_49),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_122),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_52),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_130),
.Y(n_174)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_75),
.Y(n_130)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

NAND4xp25_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_48),
.C(n_26),
.D(n_47),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_136),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_55),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_29),
.B(n_16),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_147),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_97),
.A2(n_29),
.B(n_24),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_53),
.A2(n_48),
.B1(n_23),
.B2(n_27),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_166),
.B1(n_99),
.B2(n_88),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_56),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_160),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_46),
.Y(n_160)
);

OR2x4_ASAP7_75t_L g161 ( 
.A(n_58),
.B(n_26),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_60),
.B(n_41),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_144),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_69),
.A2(n_43),
.B1(n_31),
.B2(n_40),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_84),
.B1(n_73),
.B2(n_96),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_201),
.B1(n_151),
.B2(n_135),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_92),
.B1(n_90),
.B2(n_61),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_170),
.A2(n_180),
.B1(n_181),
.B2(n_212),
.Y(n_229)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_44),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_172),
.B(n_176),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_113),
.A2(n_54),
.B1(n_57),
.B2(n_24),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_153),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_179),
.B(n_109),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_110),
.A2(n_71),
.B1(n_102),
.B2(n_98),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_68),
.B1(n_67),
.B2(n_80),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_184),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_70),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_191),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_119),
.B(n_41),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_198),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_157),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_112),
.A2(n_37),
.B1(n_44),
.B2(n_47),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_197),
.A2(n_207),
.B1(n_214),
.B2(n_126),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_114),
.B(n_37),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_148),
.A2(n_28),
.B1(n_31),
.B2(n_40),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_106),
.B(n_81),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_49),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_209),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_112),
.A2(n_39),
.B1(n_46),
.B2(n_43),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_39),
.Y(n_209)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_108),
.A2(n_40),
.B1(n_31),
.B2(n_28),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_155),
.A2(n_28),
.B1(n_43),
.B2(n_103),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_126),
.A2(n_100),
.B1(n_26),
.B2(n_3),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_187),
.B1(n_191),
.B2(n_178),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_222),
.A2(n_125),
.B1(n_210),
.B2(n_208),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_228),
.B(n_232),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_185),
.Y(n_232)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_169),
.A2(n_162),
.B(n_107),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_213),
.B(n_203),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_174),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_183),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_249),
.B(n_179),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_178),
.A2(n_108),
.B1(n_140),
.B2(n_135),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_170),
.B1(n_168),
.B2(n_180),
.Y(n_254)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_253),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_254),
.A2(n_256),
.B1(n_273),
.B2(n_193),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_169),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_257),
.C(n_264),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_178),
.C(n_204),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_248),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_260),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_177),
.B(n_175),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_240),
.B(n_239),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_248),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_265),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_280),
.Y(n_306)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_167),
.C(n_172),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_203),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_267),
.A2(n_269),
.B(n_222),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_229),
.A2(n_212),
.B1(n_181),
.B2(n_140),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_268),
.A2(n_274),
.B1(n_256),
.B2(n_219),
.Y(n_309)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_244),
.B(n_200),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_277),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_220),
.A2(n_143),
.B1(n_145),
.B2(n_205),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_229),
.A2(n_193),
.B1(n_151),
.B2(n_190),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_199),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_216),
.B(n_171),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_239),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_221),
.Y(n_286)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_279),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_223),
.B(n_210),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_252),
.B(n_109),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_235),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_286),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_288),
.A2(n_291),
.B(n_295),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_221),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_305),
.C(n_301),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_230),
.B(n_240),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_259),
.A2(n_239),
.B(n_250),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_263),
.B(n_224),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_300),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_267),
.B(n_277),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_311),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_225),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_261),
.B(n_236),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_312),
.Y(n_335)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_284),
.A2(n_235),
.B(n_226),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_276),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_219),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_300),
.Y(n_339)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_274),
.B1(n_268),
.B2(n_254),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_309),
.B1(n_297),
.B2(n_291),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_289),
.B(n_272),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_318),
.B(n_334),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g320 ( 
.A(n_302),
.Y(n_320)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_294),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_329),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_233),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_324),
.B(n_340),
.Y(n_361)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_327),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_306),
.Y(n_333)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_262),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_337),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_289),
.A2(n_273),
.B1(n_260),
.B2(n_258),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_338),
.A2(n_311),
.B1(n_288),
.B2(n_287),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_233),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_226),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_341),
.B(n_342),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_282),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_281),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_343),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_301),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_285),
.B(n_271),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_345),
.B(n_346),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_270),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_347),
.A2(n_355),
.B1(n_360),
.B2(n_375),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_319),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_293),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_356),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_305),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_317),
.A2(n_299),
.B1(n_295),
.B2(n_290),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_358),
.A2(n_373),
.B1(n_349),
.B2(n_357),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_331),
.A2(n_317),
.B(n_321),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_369),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_343),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_362),
.A2(n_365),
.B1(n_328),
.B2(n_335),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_321),
.A2(n_286),
.B1(n_287),
.B2(n_296),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_363),
.A2(n_372),
.B1(n_377),
.B2(n_338),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_334),
.B(n_296),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_364),
.B(n_371),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_318),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_346),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_366),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_330),
.A2(n_286),
.B(n_302),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_218),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_322),
.A2(n_308),
.B1(n_219),
.B2(n_243),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_308),
.B(n_227),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_337),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_345),
.A2(n_308),
.B1(n_243),
.B2(n_238),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_344),
.C(n_319),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_381),
.C(n_383),
.Y(n_411)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_368),
.Y(n_379)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_331),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_402),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_368),
.B(n_335),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_382),
.B(n_353),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_331),
.C(n_342),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_376),
.Y(n_384)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_347),
.A2(n_365),
.B1(n_362),
.B2(n_349),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_385),
.A2(n_392),
.B1(n_372),
.B2(n_377),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_396),
.B1(n_398),
.B2(n_405),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_393),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_328),
.C(n_326),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_401),
.C(n_359),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_374),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_361),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_397),
.Y(n_418)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_360),
.A2(n_316),
.B1(n_327),
.B2(n_332),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_400),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_336),
.C(n_325),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_325),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_238),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_404),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_351),
.A2(n_320),
.B1(n_234),
.B2(n_231),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_406),
.A2(n_422),
.B1(n_426),
.B2(n_427),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_410),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_351),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_380),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_413),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_359),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_420),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_383),
.C(n_391),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_387),
.A2(n_353),
.B1(n_367),
.B2(n_320),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_218),
.Y(n_423)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_423),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_403),
.Y(n_424)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_385),
.A2(n_367),
.B1(n_231),
.B2(n_227),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_400),
.Y(n_427)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_415),
.A2(n_390),
.B(n_398),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_435),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_415),
.A2(n_390),
.B1(n_396),
.B2(n_401),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_432),
.A2(n_433),
.B1(n_448),
.B2(n_426),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_419),
.A2(n_382),
.B1(n_405),
.B2(n_279),
.Y(n_433)
);

INVx13_ASAP7_75t_L g434 ( 
.A(n_421),
.Y(n_434)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_434),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_279),
.C(n_253),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_182),
.Y(n_437)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_437),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_444),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_253),
.C(n_211),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_194),
.C(n_116),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_413),
.A2(n_107),
.B(n_184),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_447),
.B(n_410),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_406),
.A2(n_188),
.B(n_124),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_417),
.A2(n_154),
.B1(n_116),
.B2(n_124),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_414),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_454),
.Y(n_480)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_439),
.A2(n_425),
.B1(n_420),
.B2(n_408),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_408),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_458),
.Y(n_470)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_456),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_407),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_196),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_460),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_154),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_131),
.B(n_117),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_463),
.A2(n_457),
.B(n_452),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_441),
.A2(n_145),
.B1(n_12),
.B2(n_26),
.Y(n_465)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_117),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_466),
.B(n_429),
.C(n_443),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_438),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_475),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_472),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_L g469 ( 
.A1(n_450),
.A2(n_431),
.B(n_433),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_469),
.A2(n_481),
.B(n_125),
.Y(n_493)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_430),
.C(n_434),
.Y(n_472)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_452),
.B(n_461),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_449),
.A2(n_437),
.B(n_447),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_156),
.B(n_137),
.Y(n_491)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_479),
.Y(n_489)
);

HAxp5_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_440),
.CON(n_481),
.SN(n_481)
);

NOR2xp67_ASAP7_75t_SL g484 ( 
.A(n_480),
.B(n_455),
.Y(n_484)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_484),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_466),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_488),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_476),
.B(n_448),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_491),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_156),
.B1(n_137),
.B2(n_133),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_137),
.Y(n_490)
);

AOI322xp5_ASAP7_75t_L g499 ( 
.A1(n_490),
.A2(n_469),
.A3(n_164),
.B1(n_133),
.B2(n_165),
.C1(n_473),
.C2(n_6),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_133),
.C(n_26),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_493),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_470),
.C(n_481),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_498),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_499),
.A2(n_500),
.B(n_501),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_164),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_164),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_496),
.A2(n_489),
.B(n_485),
.Y(n_502)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_502),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_498),
.A2(n_501),
.B(n_495),
.Y(n_503)
);

AOI322xp5_ASAP7_75t_L g507 ( 
.A1(n_503),
.A2(n_506),
.A3(n_490),
.B1(n_1),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_497),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_508),
.Y(n_511)
);

AOI322xp5_ASAP7_75t_L g508 ( 
.A1(n_505),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_8),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_509),
.Y(n_510)
);

AOI322xp5_ASAP7_75t_L g512 ( 
.A1(n_510),
.A2(n_0),
.A3(n_3),
.B1(n_5),
.B2(n_8),
.C1(n_504),
.C2(n_511),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_512),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_0),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_514),
.Y(n_515)
);


endmodule