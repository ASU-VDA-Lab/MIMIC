module real_jpeg_24385_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_0),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_0),
.B(n_50),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_0),
.B(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_0),
.B(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_59),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_2),
.B(n_43),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_2),
.B(n_50),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_2),
.B(n_131),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_2),
.B(n_211),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_67),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_3),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_3),
.B(n_43),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_3),
.B(n_36),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_3),
.B(n_40),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_3),
.B(n_50),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_3),
.B(n_131),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_3),
.B(n_211),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_4),
.B(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_4),
.B(n_36),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_40),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_4),
.B(n_50),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_4),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_4),
.B(n_304),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx8_ASAP7_75t_SL g133 ( 
.A(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_8),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_8),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_8),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_8),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_8),
.B(n_50),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_8),
.B(n_131),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_230),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_9),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_59),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_9),
.B(n_43),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_9),
.B(n_36),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_9),
.B(n_40),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_9),
.B(n_50),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_9),
.B(n_131),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_9),
.B(n_211),
.Y(n_379)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_10),
.B(n_43),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_10),
.B(n_40),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_10),
.B(n_50),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_10),
.B(n_211),
.Y(n_389)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_12),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_12),
.B(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_12),
.B(n_40),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_12),
.B(n_50),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_12),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_12),
.B(n_230),
.Y(n_276)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_14),
.B(n_67),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_59),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_14),
.B(n_43),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_14),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_14),
.B(n_40),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_14),
.B(n_50),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_14),
.B(n_230),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_36),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_16),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_17),
.Y(n_209)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_385),
.B(n_386),
.C(n_390),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_375),
.C(n_384),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_360),
.C(n_361),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_338),
.C(n_339),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_308),
.C(n_309),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_282),
.C(n_283),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_250),
.C(n_251),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_213),
.C(n_214),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_173),
.C(n_174),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_140),
.C(n_141),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_112),
.C(n_113),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_70),
.C(n_83),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_53),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_33),
.B(n_45),
.C(n_53),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.C(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_34),
.A2(n_35),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_48),
.C(n_49),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_62),
.C(n_63),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_65),
.B(n_69),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.C(n_82),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_75),
.B1(n_82),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_81),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_108),
.C(n_109),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.C(n_98),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_90),
.C(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.C(n_103),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_126),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_127),
.C(n_139),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_121),
.C(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_120),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_122),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.CI(n_125),
.CON(n_122),
.SN(n_122)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_124),
.C(n_125),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_139),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_137),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_132),
.B(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_132),
.B(n_220),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_132),
.B(n_235),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_136),
.C(n_138),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_156),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_145),
.C(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_152),
.C(n_155),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_147),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.CI(n_150),
.CON(n_147),
.SN(n_147)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_163),
.C(n_171),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_163),
.B1(n_171),
.B2(n_172),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_162),
.B(n_199),
.C(n_200),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_169),
.C(n_170),
.Y(n_194)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_167),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_195),
.B2(n_212),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_196),
.C(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_179),
.C(n_188),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_184),
.C(n_187),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_182),
.B(n_235),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_192),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_210),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_205),
.C(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_204),
.B(n_235),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_248),
.B2(n_249),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_239),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_239),
.C(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_227),
.C(n_228),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_219),
.B(n_222),
.C(n_224),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_238),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_234),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_237),
.C(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_233),
.B(n_257),
.C(n_260),
.Y(n_306)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_246),
.C(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_254),
.C(n_281),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_268),
.B2(n_281),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_263),
.C(n_264),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_260),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_261),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_SL g323 ( 
.A(n_260),
.B(n_287),
.C(n_290),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_264),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.CI(n_267),
.CON(n_264),
.SN(n_264)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_280),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_276),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_278),
.B1(n_303),
.B2(n_305),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_305),
.C(n_306),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_307),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_297),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_297),
.C(n_307),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_292),
.C(n_293),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_290),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_SL g349 ( 
.A(n_290),
.B(n_316),
.C(n_318),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_293),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.CI(n_296),
.CON(n_293),
.SN(n_293)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_303),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_312),
.C(n_325),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_324),
.B2(n_325),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_320),
.B2(n_321),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_322),
.C(n_323),
.Y(n_341)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_318),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_318),
.A2(n_319),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_354),
.C(n_355),
.Y(n_367)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_328),
.C(n_331),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_334),
.C(n_337),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_336),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_339)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_342),
.C(n_359),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_348),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_349),
.C(n_350),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_344),
.B(n_362),
.C(n_364),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.CI(n_347),
.CON(n_344),
.SN(n_344)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_355),
.B2(n_356),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_351),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_352),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_353),
.A2(n_354),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_371),
.C(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_367),
.C(n_368),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_373),
.B2(n_374),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_371),
.A2(n_372),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_372),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_SL g391 ( 
.A(n_372),
.B(n_379),
.C(n_382),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_373),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_383),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_378),
.C(n_383),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_381),
.A2(n_382),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_382),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_389),
.Y(n_390)
);


endmodule