module fake_jpeg_4567_n_99 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_99);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_22),
.B1(n_13),
.B2(n_21),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_27),
.A2(n_30),
.B1(n_5),
.B2(n_8),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_44),
.Y(n_67)
);

HB1xp67_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_43),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_50),
.B1(n_9),
.B2(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_24),
.A2(n_16),
.B1(n_17),
.B2(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_24),
.A2(n_29),
.B1(n_17),
.B2(n_16),
.Y(n_51)
);

OAI22x1_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_32),
.B1(n_25),
.B2(n_3),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_3),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_25),
.B(n_32),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_34),
.C(n_52),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_38),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_66),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_11),
.B1(n_50),
.B2(n_38),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_51),
.B(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_64),
.B1(n_55),
.B2(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_40),
.B1(n_35),
.B2(n_47),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_77),
.C(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_76),
.Y(n_86)
);

XOR2x2_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_39),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_61),
.C(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_39),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_59),
.B(n_66),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_80),
.B(n_77),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_56),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_84),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_69),
.C(n_68),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_88),
.B(n_90),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_78),
.B(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

AOI21x1_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_68),
.B(n_81),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_52),
.A3(n_61),
.B1(n_65),
.B2(n_80),
.C1(n_82),
.C2(n_95),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.C(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_96),
.Y(n_99)
);


endmodule