module real_aes_18167_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_845, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_845;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g813 ( .A(n_0), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_1), .A2(n_33), .B1(n_125), .B2(n_148), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_2), .A2(n_9), .B1(n_167), .B2(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g814 ( .A(n_3), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_4), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_5), .A2(n_10), .B1(n_184), .B2(n_187), .Y(n_183) );
OR2x2_ASAP7_75t_L g797 ( .A(n_6), .B(n_30), .Y(n_797) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_7), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_8), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_11), .B(n_128), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_12), .A2(n_97), .B1(n_167), .B2(n_168), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_13), .A2(n_29), .B1(n_133), .B2(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_14), .A2(n_17), .B1(n_791), .B2(n_792), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_14), .Y(n_791) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_15), .B(n_128), .Y(n_127) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_16), .A2(n_45), .B(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g792 ( .A(n_17), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_18), .B(n_491), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_19), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_20), .A2(n_37), .B1(n_153), .B2(n_154), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_21), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_22), .A2(n_43), .B1(n_154), .B2(n_167), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_23), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_24), .B(n_133), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_25), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_26), .B(n_185), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_27), .B(n_142), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_28), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_31), .A2(n_81), .B1(n_125), .B2(n_223), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_32), .A2(n_36), .B1(n_124), .B2(n_125), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_34), .A2(n_48), .B1(n_167), .B2(n_171), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_35), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_38), .B(n_128), .Y(n_474) );
INVx2_ASAP7_75t_L g812 ( .A(n_39), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_40), .A2(n_51), .B1(n_826), .B2(n_827), .Y(n_825) );
INVx1_ASAP7_75t_L g827 ( .A(n_40), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_40), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_41), .B(n_129), .Y(n_486) );
BUFx3_ASAP7_75t_L g796 ( .A(n_42), .Y(n_796) );
INVx1_ASAP7_75t_L g807 ( .A(n_42), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_44), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g534 ( .A(n_46), .B(n_494), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_47), .B(n_201), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_49), .B(n_185), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_50), .B(n_153), .Y(n_610) );
INVx1_ASAP7_75t_L g826 ( .A(n_51), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_52), .A2(n_68), .B1(n_153), .B2(n_171), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_53), .A2(n_71), .B1(n_124), .B2(n_125), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_54), .B(n_519), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_55), .A2(n_226), .B(n_475), .C(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_56), .A2(n_93), .B1(n_167), .B2(n_187), .Y(n_213) );
INVx1_ASAP7_75t_L g120 ( .A(n_57), .Y(n_120) );
AND2x4_ASAP7_75t_L g139 ( .A(n_58), .B(n_140), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_59), .A2(n_60), .B1(n_154), .B2(n_204), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_61), .B(n_142), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_62), .B(n_494), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_63), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_64), .B(n_154), .Y(n_479) );
INVx1_ASAP7_75t_L g140 ( .A(n_65), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_66), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_67), .B(n_142), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_69), .B(n_125), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_70), .B(n_129), .C(n_148), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_72), .B(n_125), .Y(n_541) );
INVx2_ASAP7_75t_L g130 ( .A(n_73), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g461 ( .A(n_74), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_74), .A2(n_461), .B1(n_825), .B2(n_828), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_75), .B(n_190), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_76), .B(n_128), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_77), .B(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_78), .A2(n_94), .B1(n_154), .B2(n_226), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_79), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_80), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_82), .A2(n_88), .B1(n_185), .B2(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g817 ( .A(n_83), .B(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_84), .B(n_128), .Y(n_607) );
NAND2xp33_ASAP7_75t_SL g559 ( .A(n_85), .B(n_134), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_86), .B(n_169), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_87), .B(n_142), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_89), .Y(n_194) );
INVx1_ASAP7_75t_L g458 ( .A(n_90), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_90), .B(n_806), .Y(n_805) );
NAND2xp33_ASAP7_75t_L g135 ( .A(n_91), .B(n_128), .Y(n_135) );
NAND2xp33_ASAP7_75t_L g542 ( .A(n_92), .B(n_134), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_95), .B(n_494), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_96), .B(n_134), .C(n_190), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_98), .B(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_99), .B(n_125), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_100), .B(n_185), .Y(n_517) );
A2O1A1O1Ixp25_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_793), .B(n_798), .C(n_801), .D(n_815), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_789), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp33_ASAP7_75t_L g793 ( .A1(n_104), .A2(n_790), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_459), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_454), .Y(n_107) );
NAND2x1p5_ASAP7_75t_L g108 ( .A(n_109), .B(n_398), .Y(n_108) );
NOR3x1_ASAP7_75t_L g109 ( .A(n_110), .B(n_316), .C(n_353), .Y(n_109) );
NAND4xp75_ASAP7_75t_L g110 ( .A(n_111), .B(n_236), .C(n_270), .D(n_300), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI32xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_158), .A3(n_208), .B1(n_217), .B2(n_231), .Y(n_112) );
OR2x2_ASAP7_75t_L g217 ( .A(n_113), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_114), .A2(n_428), .B(n_430), .Y(n_427) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_143), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_115), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g299 ( .A(n_115), .B(n_245), .Y(n_299) );
AND2x2_ASAP7_75t_L g394 ( .A(n_115), .B(n_210), .Y(n_394) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g243 ( .A(n_116), .Y(n_243) );
OAI21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_141), .Y(n_116) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_117), .A2(n_121), .B(n_141), .Y(n_276) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx4_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_118), .B(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g205 ( .A(n_118), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_118), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_118), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g470 ( .A(n_118), .Y(n_470) );
AND2x4_ASAP7_75t_SL g549 ( .A(n_118), .B(n_480), .Y(n_549) );
INVx1_ASAP7_75t_SL g552 ( .A(n_118), .Y(n_552) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g175 ( .A(n_119), .Y(n_175) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_131), .B(n_137), .Y(n_121) );
O2A1O1Ixp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B(n_127), .C(n_129), .Y(n_122) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
INVx1_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_125), .A2(n_154), .B1(n_532), .B2(n_533), .Y(n_531) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_126), .Y(n_128) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_126), .Y(n_148) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx1_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
INVx1_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
INVx1_ASAP7_75t_L g201 ( .A(n_126), .Y(n_201) );
INVx1_ASAP7_75t_L g204 ( .A(n_126), .Y(n_204) );
INVx2_ASAP7_75t_L g224 ( .A(n_126), .Y(n_224) );
INVx1_ASAP7_75t_L g226 ( .A(n_126), .Y(n_226) );
INVx3_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx1_ASAP7_75t_L g491 ( .A(n_128), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_128), .A2(n_555), .B(n_556), .Y(n_554) );
INVx6_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_129), .A2(n_478), .B(n_479), .Y(n_477) );
O2A1O1Ixp5_ASAP7_75t_L g605 ( .A1(n_129), .A2(n_168), .B(n_606), .C(n_607), .Y(n_605) );
BUFx8_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g151 ( .A(n_130), .Y(n_151) );
INVx1_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
INVx1_ASAP7_75t_L g476 ( .A(n_130), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_135), .B(n_136), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g153 ( .A(n_134), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_136), .A2(n_147), .B1(n_149), .B2(n_152), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_136), .A2(n_149), .B1(n_166), .B2(n_170), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_136), .A2(n_183), .B1(n_188), .B2(n_189), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_136), .A2(n_149), .B1(n_199), .B2(n_202), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_136), .A2(n_189), .B1(n_213), .B2(n_214), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_136), .A2(n_222), .B1(n_225), .B2(n_227), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_136), .A2(n_149), .B1(n_261), .B2(n_262), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_136), .A2(n_149), .B1(n_497), .B2(n_499), .Y(n_496) );
INVx2_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_SL g228 ( .A(n_138), .Y(n_228) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx10_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx10_ASAP7_75t_L g480 ( .A(n_139), .Y(n_480) );
INVx2_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
INVx2_ASAP7_75t_L g267 ( .A(n_143), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_143), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_144), .Y(n_254) );
INVx1_ASAP7_75t_L g298 ( .A(n_144), .Y(n_298) );
AND2x2_ASAP7_75t_L g342 ( .A(n_144), .B(n_276), .Y(n_342) );
OR2x2_ASAP7_75t_L g396 ( .A(n_144), .B(n_220), .Y(n_396) );
AO31x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .A3(n_155), .B(n_156), .Y(n_144) );
INVx2_ASAP7_75t_L g164 ( .A(n_145), .Y(n_164) );
AO31x2_ASAP7_75t_L g181 ( .A1(n_145), .A2(n_182), .A3(n_191), .B(n_193), .Y(n_181) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_145), .A2(n_198), .A3(n_205), .B(n_206), .Y(n_197) );
AO31x2_ASAP7_75t_L g495 ( .A1(n_145), .A2(n_174), .A3(n_496), .B(n_500), .Y(n_495) );
INVx2_ASAP7_75t_L g519 ( .A(n_148), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_149), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g520 ( .A(n_150), .Y(n_520) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g546 ( .A(n_151), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_154), .A2(n_486), .B(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g498 ( .A(n_154), .Y(n_498) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_159), .A2(n_322), .B1(n_414), .B2(n_416), .Y(n_413) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_179), .Y(n_159) );
INVx4_ASAP7_75t_L g239 ( .A(n_160), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_160), .A2(n_219), .B1(n_251), .B2(n_253), .Y(n_250) );
OR2x2_ASAP7_75t_L g256 ( .A(n_160), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g375 ( .A(n_160), .B(n_274), .Y(n_375) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g295 ( .A(n_161), .B(n_180), .Y(n_295) );
AND2x2_ASAP7_75t_L g386 ( .A(n_161), .B(n_258), .Y(n_386) );
AND2x2_ASAP7_75t_L g441 ( .A(n_161), .B(n_197), .Y(n_441) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g235 ( .A(n_162), .Y(n_235) );
AND2x4_ASAP7_75t_L g362 ( .A(n_162), .B(n_258), .Y(n_362) );
AO31x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .A3(n_172), .B(n_176), .Y(n_162) );
AO31x2_ASAP7_75t_L g211 ( .A1(n_163), .A2(n_191), .A3(n_212), .B(n_215), .Y(n_211) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp67_ASAP7_75t_SL g525 ( .A(n_164), .B(n_173), .Y(n_525) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO31x2_ASAP7_75t_L g259 ( .A1(n_172), .A2(n_228), .A3(n_260), .B(n_263), .Y(n_259) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g193 ( .A(n_174), .B(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_174), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g178 ( .A(n_175), .Y(n_178) );
INVx2_ASAP7_75t_L g192 ( .A(n_175), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_178), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g494 ( .A(n_178), .Y(n_494) );
INVx2_ASAP7_75t_L g521 ( .A(n_178), .Y(n_521) );
NAND2x1_ASAP7_75t_L g238 ( .A(n_179), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_179), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_195), .Y(n_179) );
INVx2_ASAP7_75t_L g233 ( .A(n_180), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_180), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g281 ( .A(n_180), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_180), .B(n_283), .Y(n_308) );
AND2x2_ASAP7_75t_L g311 ( .A(n_180), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g371 ( .A(n_180), .Y(n_371) );
INVx4_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_181), .B(n_196), .Y(n_249) );
BUFx2_ASAP7_75t_L g287 ( .A(n_181), .Y(n_287) );
AND2x2_ASAP7_75t_L g336 ( .A(n_181), .B(n_197), .Y(n_336) );
AND2x2_ASAP7_75t_L g378 ( .A(n_181), .B(n_259), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_181), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx1_ASAP7_75t_L g492 ( .A(n_190), .Y(n_492) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_192), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_197), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g289 ( .A(n_197), .B(n_259), .Y(n_289) );
INVx1_ASAP7_75t_L g312 ( .A(n_197), .Y(n_312) );
INVx2_ASAP7_75t_L g332 ( .A(n_197), .Y(n_332) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_197), .Y(n_377) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AO31x2_ASAP7_75t_L g220 ( .A1(n_205), .A2(n_221), .A3(n_228), .B(n_229), .Y(n_220) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g296 ( .A(n_209), .B(n_297), .Y(n_296) );
NOR2x1p5_ASAP7_75t_L g402 ( .A(n_209), .B(n_396), .Y(n_402) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x4_ASAP7_75t_L g219 ( .A(n_210), .B(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_210), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_210), .B(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g244 ( .A(n_211), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g302 ( .A(n_211), .B(n_220), .Y(n_302) );
BUFx2_ASAP7_75t_L g415 ( .A(n_211), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_217), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g453 ( .A(n_217), .Y(n_453) );
INVx2_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g389 ( .A(n_219), .Y(n_389) );
AND2x4_ASAP7_75t_L g412 ( .A(n_219), .B(n_342), .Y(n_412) );
AND2x2_ASAP7_75t_L g436 ( .A(n_219), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g245 ( .A(n_220), .Y(n_245) );
BUFx2_ASAP7_75t_L g269 ( .A(n_220), .Y(n_269) );
INVx1_ASAP7_75t_L g325 ( .A(n_220), .Y(n_325) );
OR2x2_ASAP7_75t_L g447 ( .A(n_220), .B(n_304), .Y(n_447) );
INVx2_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_224), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g547 ( .A(n_226), .Y(n_547) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g293 ( .A(n_233), .Y(n_293) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_234), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_234), .Y(n_314) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g255 ( .A(n_235), .Y(n_255) );
OR2x2_ASAP7_75t_L g292 ( .A(n_235), .B(n_284), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_240), .B(n_246), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_241), .A2(n_335), .B1(n_337), .B2(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
OR2x2_ASAP7_75t_L g380 ( .A(n_243), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g388 ( .A(n_243), .Y(n_388) );
AND2x2_ASAP7_75t_L g401 ( .A(n_243), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g363 ( .A(n_244), .B(n_342), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_250), .B1(n_256), .B2(n_265), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g315 ( .A(n_249), .Y(n_315) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g273 ( .A(n_252), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g341 ( .A(n_252), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g350 ( .A(n_252), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_252), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_253), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g338 ( .A(n_255), .B(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g352 ( .A(n_255), .Y(n_352) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
AND2x4_ASAP7_75t_L g331 ( .A(n_259), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_259), .Y(n_347) );
INVx1_ASAP7_75t_L g411 ( .A(n_259), .Y(n_411) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
AND2x4_ASAP7_75t_L g303 ( .A(n_267), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g320 ( .A(n_267), .Y(n_320) );
INVx1_ASAP7_75t_L g278 ( .A(n_269), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_279), .B1(n_290), .B2(n_296), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2x1p5_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVxp67_ASAP7_75t_SL g328 ( .A(n_275), .Y(n_328) );
INVx1_ASAP7_75t_L g304 ( .A(n_276), .Y(n_304) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_285), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_281), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g433 ( .A(n_282), .Y(n_433) );
INVx1_ASAP7_75t_L g452 ( .A(n_282), .Y(n_452) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2x1_ASAP7_75t_L g429 ( .A(n_286), .B(n_352), .Y(n_429) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g445 ( .A(n_287), .Y(n_445) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx2_ASAP7_75t_L g383 ( .A(n_291), .Y(n_383) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx2_ASAP7_75t_L g372 ( .A(n_292), .Y(n_372) );
AND2x4_ASAP7_75t_L g374 ( .A(n_293), .B(n_331), .Y(n_374) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_297), .A2(n_443), .B1(n_446), .B2(n_448), .Y(n_442) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g367 ( .A(n_298), .Y(n_367) );
INVx1_ASAP7_75t_L g321 ( .A(n_299), .Y(n_321) );
AND2x4_ASAP7_75t_L g414 ( .A(n_299), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g422 ( .A(n_299), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
AND2x4_ASAP7_75t_SL g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_SL g365 ( .A(n_302), .Y(n_365) );
INVx2_ASAP7_75t_L g381 ( .A(n_302), .Y(n_381) );
INVx1_ASAP7_75t_L g408 ( .A(n_303), .Y(n_408) );
AND2x2_ASAP7_75t_L g439 ( .A(n_303), .B(n_350), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .C(n_313), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_310), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g351 ( .A(n_311), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_311), .B(n_386), .Y(n_419) );
INVx1_ASAP7_75t_L g339 ( .A(n_312), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_314), .B(n_378), .Y(n_404) );
INVx1_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
NAND3xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_333), .C(n_343), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .B(n_329), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g437 ( .A(n_320), .Y(n_437) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI32xp33_ASAP7_75t_L g373 ( .A1(n_324), .A2(n_374), .A3(n_375), .B1(n_376), .B2(n_379), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_324), .B(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g357 ( .A(n_331), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_331), .B(n_352), .Y(n_392) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_336), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g397 ( .A(n_336), .B(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g425 ( .A(n_339), .Y(n_425) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g343 ( .A1(n_341), .A2(n_344), .B1(n_348), .B2(n_351), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_342), .B(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_344), .A2(n_402), .B1(n_439), .B2(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g440 ( .A(n_346), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_348), .A2(n_391), .B1(n_393), .B2(n_397), .Y(n_390) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g432 ( .A(n_352), .Y(n_432) );
NAND4xp25_ASAP7_75t_L g353 ( .A(n_354), .B(n_373), .C(n_382), .D(n_390), .Y(n_353) );
O2A1O1Ixp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_360), .B(n_363), .C(n_364), .Y(n_354) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g418 ( .A(n_362), .B(n_377), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_362), .B(n_445), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B(n_368), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_369), .A2(n_407), .B1(n_409), .B2(n_412), .Y(n_406) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_374), .A2(n_379), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI21xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_387), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_R g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_397), .A2(n_414), .B1(n_451), .B2(n_453), .Y(n_450) );
NOR3x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_420), .C(n_434), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_413), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_405), .Y(n_400) );
INVx1_ASAP7_75t_L g426 ( .A(n_401), .Y(n_426) );
INVx2_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
INVx1_ASAP7_75t_L g423 ( .A(n_415), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_417), .A2(n_421), .B1(n_424), .B2(n_426), .C(n_427), .Y(n_420) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
NAND4xp25_ASAP7_75t_SL g434 ( .A(n_435), .B(n_438), .C(n_442), .D(n_450), .Y(n_434) );
AND2x2_ASAP7_75t_L g448 ( .A(n_441), .B(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx12f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g800 ( .A(n_457), .B(n_795), .Y(n_800) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g788 ( .A(n_458), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_785), .Y(n_459) );
XNOR2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
BUFx2_ASAP7_75t_L g822 ( .A(n_462), .Y(n_822) );
NAND2x1p5_ASAP7_75t_SL g462 ( .A(n_463), .B(n_719), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_655), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_577), .C(n_616), .D(n_645), .Y(n_464) );
O2A1O1Ixp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_502), .B(n_509), .C(n_561), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_482), .Y(n_466) );
INVx2_ASAP7_75t_L g505 ( .A(n_467), .Y(n_505) );
AND2x2_ASAP7_75t_L g643 ( .A(n_467), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_467), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_467), .B(n_563), .Y(n_738) );
OR2x2_ASAP7_75t_L g774 ( .A(n_467), .B(n_690), .Y(n_774) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g671 ( .A(n_468), .B(n_483), .Y(n_671) );
NOR2xp67_ASAP7_75t_L g697 ( .A(n_468), .B(n_507), .Y(n_697) );
BUFx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g632 ( .A(n_469), .Y(n_632) );
OAI21x1_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_481), .Y(n_469) );
OAI21x1_ASAP7_75t_L g483 ( .A1(n_470), .A2(n_484), .B(n_493), .Y(n_483) );
OAI21x1_ASAP7_75t_L g565 ( .A1(n_470), .A2(n_471), .B(n_481), .Y(n_565) );
OA21x2_ASAP7_75t_L g600 ( .A1(n_470), .A2(n_484), .B(n_493), .Y(n_600) );
OAI21x1_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_477), .B(n_480), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_475), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_475), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_475), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_475), .A2(n_558), .B(n_559), .Y(n_557) );
BUFx4f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI21x1_ASAP7_75t_L g484 ( .A1(n_480), .A2(n_485), .B(n_488), .Y(n_484) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_480), .A2(n_513), .B(n_516), .Y(n_512) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_480), .A2(n_554), .B(n_557), .Y(n_553) );
OAI21x1_ASAP7_75t_L g604 ( .A1(n_480), .A2(n_605), .B(n_608), .Y(n_604) );
AND2x2_ASAP7_75t_L g571 ( .A(n_482), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_482), .B(n_601), .Y(n_615) );
AND2x2_ASAP7_75t_L g623 ( .A(n_482), .B(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_482), .Y(n_646) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .Y(n_482) );
INVx1_ASAP7_75t_L g507 ( .A(n_483), .Y(n_507) );
INVx1_ASAP7_75t_L g563 ( .A(n_483), .Y(n_563) );
AND2x2_ASAP7_75t_L g633 ( .A(n_483), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g694 ( .A(n_483), .B(n_602), .Y(n_694) );
AOI21x1_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_492), .Y(n_488) );
INVx1_ASAP7_75t_L g508 ( .A(n_495), .Y(n_508) );
AND2x2_ASAP7_75t_L g564 ( .A(n_495), .B(n_565), .Y(n_564) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_495), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_495), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g677 ( .A(n_495), .B(n_632), .Y(n_677) );
OR2x2_ASAP7_75t_L g690 ( .A(n_495), .B(n_600), .Y(n_690) );
OR2x2_ASAP7_75t_L g700 ( .A(n_495), .B(n_565), .Y(n_700) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_505), .B(n_716), .Y(n_762) );
INVx1_ASAP7_75t_L g618 ( .A(n_506), .Y(n_618) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_L g702 ( .A(n_508), .B(n_565), .Y(n_702) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_535), .Y(n_509) );
AND2x2_ASAP7_75t_L g575 ( .A(n_510), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g637 ( .A(n_510), .Y(n_637) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_523), .Y(n_510) );
BUFx2_ASAP7_75t_L g744 ( .A(n_511), .Y(n_744) );
OAI21xp33_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_521), .B(n_522), .Y(n_511) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_512), .A2(n_521), .B(n_522), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_520), .Y(n_516) );
OAI21x1_ASAP7_75t_L g603 ( .A1(n_521), .A2(n_604), .B(n_611), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_521), .A2(n_604), .B(n_611), .Y(n_634) );
AND2x2_ASAP7_75t_L g583 ( .A(n_523), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g569 ( .A(n_524), .B(n_551), .Y(n_569) );
INVx2_ASAP7_75t_L g595 ( .A(n_524), .Y(n_595) );
AOI21x1_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_534), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_530), .Y(n_526) );
AND2x2_ASAP7_75t_L g741 ( .A(n_535), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_550), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx4_ASAP7_75t_L g568 ( .A(n_537), .Y(n_568) );
BUFx2_ASAP7_75t_L g576 ( .A(n_537), .Y(n_576) );
OR2x2_ASAP7_75t_L g580 ( .A(n_537), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g640 ( .A(n_537), .B(n_584), .Y(n_640) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .B(n_549), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_546), .B1(n_547), .B2(n_548), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_545), .A2(n_609), .B(n_610), .Y(n_608) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g627 ( .A(n_550), .Y(n_627) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_550), .Y(n_641) );
INVx2_ASAP7_75t_L g666 ( .A(n_550), .Y(n_666) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g581 ( .A(n_551), .Y(n_581) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B(n_560), .Y(n_551) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_566), .B1(n_570), .B2(n_574), .Y(n_561) );
INVx1_ASAP7_75t_L g651 ( .A(n_562), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g662 ( .A(n_563), .Y(n_662) );
AND2x2_ASAP7_75t_L g679 ( .A(n_564), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_564), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g573 ( .A(n_565), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_566), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_567), .B(n_583), .Y(n_674) );
AND2x2_ASAP7_75t_L g682 ( .A(n_567), .B(n_648), .Y(n_682) );
AND2x2_ASAP7_75t_L g758 ( .A(n_567), .B(n_705), .Y(n_758) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g593 ( .A(n_568), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g614 ( .A(n_568), .B(n_584), .Y(n_614) );
OR2x2_ASAP7_75t_L g626 ( .A(n_568), .B(n_627), .Y(n_626) );
NAND2x1_ASAP7_75t_L g660 ( .A(n_568), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g665 ( .A(n_568), .Y(n_665) );
INVx2_ASAP7_75t_L g659 ( .A(n_569), .Y(n_659) );
AND2x2_ASAP7_75t_L g685 ( .A(n_569), .B(n_649), .Y(n_685) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_572), .Y(n_621) );
INVx1_ASAP7_75t_L g688 ( .A(n_572), .Y(n_688) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g672 ( .A(n_573), .B(n_602), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_574), .A2(n_684), .B(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g745 ( .A(n_576), .B(n_685), .Y(n_745) );
INVx1_ASAP7_75t_L g781 ( .A(n_576), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_586), .B(n_590), .Y(n_577) );
AOI322xp5_ASAP7_75t_L g729 ( .A1(n_578), .A2(n_625), .A3(n_730), .B1(n_731), .B2(n_732), .C1(n_733), .C2(n_736), .Y(n_729) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g717 ( .A(n_580), .B(n_582), .C(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g596 ( .A(n_581), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g725 ( .A(n_581), .B(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_581), .Y(n_777) );
OR2x2_ASAP7_75t_L g673 ( .A(n_582), .B(n_626), .Y(n_673) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g661 ( .A(n_584), .Y(n_661) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g597 ( .A(n_585), .Y(n_597) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_587), .Y(n_722) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g693 ( .A(n_588), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_589), .B(n_716), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_598), .B(n_612), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_592), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
AND2x2_ASAP7_75t_L g648 ( .A(n_594), .B(n_649), .Y(n_648) );
AND3x2_ASAP7_75t_L g692 ( .A(n_594), .B(n_596), .C(n_665), .Y(n_692) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g654 ( .A(n_595), .Y(n_654) );
AND2x2_ASAP7_75t_L g705 ( .A(n_595), .B(n_666), .Y(n_705) );
INVx2_ASAP7_75t_L g728 ( .A(n_595), .Y(n_728) );
AND2x2_ASAP7_75t_L g732 ( .A(n_596), .B(n_728), .Y(n_732) );
INVx2_ASAP7_75t_L g649 ( .A(n_597), .Y(n_649) );
OR2x2_ASAP7_75t_L g783 ( .A(n_597), .B(n_666), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_598), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g735 ( .A(n_599), .Y(n_735) );
AND2x2_ASAP7_75t_L g644 ( .A(n_600), .B(n_634), .Y(n_644) );
AND2x2_ASAP7_75t_L g680 ( .A(n_600), .B(n_602), .Y(n_680) );
AND2x2_ASAP7_75t_L g676 ( .A(n_601), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_601), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g748 ( .A(n_601), .Y(n_748) );
BUFx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g619 ( .A(n_602), .Y(n_619) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_602), .Y(n_624) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_602), .Y(n_670) );
INVx1_ASAP7_75t_L g716 ( .A(n_602), .Y(n_716) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_625), .B(n_628), .Y(n_616) );
OAI31xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .A3(n_620), .B(n_622), .Y(n_617) );
INVx1_ASAP7_75t_L g699 ( .A(n_619), .Y(n_699) );
OAI32xp33_ASAP7_75t_L g657 ( .A1(n_620), .A2(n_629), .A3(n_658), .B1(n_662), .B2(n_663), .Y(n_657) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g650 ( .A(n_626), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_635), .B1(n_638), .B2(n_642), .Y(n_628) );
OAI22xp33_ASAP7_75t_SL g713 ( .A1(n_629), .A2(n_674), .B1(n_714), .B2(n_715), .Y(n_713) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx2_ASAP7_75t_L g771 ( .A(n_631), .Y(n_771) );
BUFx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g726 ( .A(n_634), .Y(n_726) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g652 ( .A(n_640), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g727 ( .A(n_640), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g778 ( .A(n_640), .Y(n_778) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g718 ( .A(n_644), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_651), .B2(n_652), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_647), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
AND2x2_ASAP7_75t_L g704 ( .A(n_649), .B(n_665), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_652), .A2(n_710), .B(n_713), .C(n_717), .Y(n_709) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_654), .Y(n_767) );
INVx1_ASAP7_75t_L g784 ( .A(n_654), .Y(n_784) );
NAND4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_678), .C(n_691), .D(n_709), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_667), .Y(n_656) );
OR2x6_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_661), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g766 ( .A(n_664), .B(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_667) );
NOR2xp33_ASAP7_75t_SL g668 ( .A(n_669), .B(n_672), .Y(n_668) );
BUFx2_ASAP7_75t_L g681 ( .A(n_669), .Y(n_681) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_675), .B(n_761), .Y(n_760) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g730 ( .A(n_677), .B(n_716), .Y(n_730) );
O2A1O1Ixp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B(n_682), .C(n_683), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_680), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g740 ( .A(n_687), .B(n_741), .Y(n_740) );
AND2x4_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_703), .C(n_706), .Y(n_691) );
AND2x2_ASAP7_75t_L g770 ( .A(n_694), .B(n_771), .Y(n_770) );
NAND3xp33_ASAP7_75t_SL g695 ( .A(n_696), .B(n_698), .C(n_701), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_699), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_699), .B(n_735), .Y(n_765) );
INVx1_ASAP7_75t_L g708 ( .A(n_700), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_700), .Y(n_712) );
AND2x2_ASAP7_75t_L g753 ( .A(n_702), .B(n_742), .Y(n_753) );
NAND2xp33_ASAP7_75t_SL g754 ( .A(n_702), .B(n_724), .Y(n_754) );
AND2x4_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g714 ( .A(n_705), .Y(n_714) );
NOR3x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_749), .C(n_768), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_729), .C(n_739), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g742 ( .A(n_726), .Y(n_742) );
INVx2_ASAP7_75t_L g731 ( .A(n_728), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_730), .A2(n_773), .B1(n_780), .B2(n_845), .Y(n_779) );
O2A1O1Ixp5_ASAP7_75t_L g751 ( .A1(n_731), .A2(n_743), .B(n_752), .C(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AO21x1_ASAP7_75t_L g755 ( .A1(n_734), .A2(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g747 ( .A(n_738), .B(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B1(n_745), .B2(n_746), .Y(n_739) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND4xp75_ASAP7_75t_L g749 ( .A(n_750), .B(n_755), .C(n_759), .D(n_763), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .C(n_779), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_775), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVxp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OR2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
AND2x4_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
NOR2x1p5_ASAP7_75t_SL g782 ( .A(n_783), .B(n_784), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g808 ( .A(n_797), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_809), .Y(n_801) );
INVx3_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
CKINVDCx8_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_L g818 ( .A(n_804), .Y(n_818) );
INVx3_ASAP7_75t_L g831 ( .A(n_804), .Y(n_831) );
AND2x6_ASAP7_75t_SL g804 ( .A(n_805), .B(n_808), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g809 ( .A(n_810), .B(n_813), .Y(n_809) );
BUFx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_811), .B(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_812), .B(n_831), .Y(n_843) );
INVx2_ASAP7_75t_SL g840 ( .A(n_813), .Y(n_840) );
A2O1A1Ixp33_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_819), .B(n_834), .C(n_841), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVxp67_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI22xp5_ASAP7_75t_SL g820 ( .A1(n_821), .A2(n_822), .B1(n_823), .B2(n_832), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_829), .Y(n_823) );
INVx1_ASAP7_75t_L g833 ( .A(n_824), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_825), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_829), .B(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
INVx4_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
BUFx3_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
OR2x4_ASAP7_75t_L g842 ( .A(n_839), .B(n_843), .Y(n_842) );
BUFx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
endmodule