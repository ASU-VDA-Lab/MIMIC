module fake_netlist_6_4584_n_1264 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1264);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1264;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_1094;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_177;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_172;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_87),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_7),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_25),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_86),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_104),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_33),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_74),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_45),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_58),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_48),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_50),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_55),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_67),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_129),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_27),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_31),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_21),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_16),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_55),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_58),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_18),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_48),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_128),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_166),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_60),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_28),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_79),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_28),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_95),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_0),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_159),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_98),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_49),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_17),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_101),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_30),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_168),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_19),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_139),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_54),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_6),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_41),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_12),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_82),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_85),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_81),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_24),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_3),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_150),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_66),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_72),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_68),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_4),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_54),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_124),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_130),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_116),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_153),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_8),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_61),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_143),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_120),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_19),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_13),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_117),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_93),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_91),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_165),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_69),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_7),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_64),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_126),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_158),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_33),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_144),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_9),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_152),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_140),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_147),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_30),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_108),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_146),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_51),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_88),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_134),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_154),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_11),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_59),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_197),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_0),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_178),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_194),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_203),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_207),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_222),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_1),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_210),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_171),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_1),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_241),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_213),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_221),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_246),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_171),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_252),
.B(n_2),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_172),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_224),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_190),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_190),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_190),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_190),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_190),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_195),
.B(n_3),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_192),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_191),
.B(n_196),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_226),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_192),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_268),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_229),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_277),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_172),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_240),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_214),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_215),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_180),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_242),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_214),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_244),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_263),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_255),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_219),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_244),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_256),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_257),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_211),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_261),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_217),
.B(n_4),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_262),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_266),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_267),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_206),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_216),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_218),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_195),
.B(n_5),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_211),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_232),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_223),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_201),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_232),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_217),
.B(n_6),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_202),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_173),
.B(n_9),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_227),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_184),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_204),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_170),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_228),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_208),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_225),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_184),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_R g374 ( 
.A(n_170),
.B(n_62),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_174),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_231),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_235),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_236),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_237),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_238),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_245),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_291),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_351),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_250),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_291),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_318),
.B(n_250),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_174),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_258),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_298),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_175),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_304),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_291),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_291),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_291),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_302),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_313),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_302),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_305),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_305),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_307),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_316),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_307),
.B(n_258),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_308),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_308),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_315),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_315),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_306),
.B(n_173),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_347),
.B(n_233),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_360),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

BUFx8_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_324),
.Y(n_423)
);

CKINVDCx8_ASAP7_75t_R g424 ( 
.A(n_353),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_314),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_233),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_364),
.B(n_175),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_357),
.B(n_177),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_362),
.B(n_177),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_327),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_334),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_327),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_333),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_363),
.B(n_181),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_325),
.A2(n_269),
.B(n_179),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_333),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_337),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_363),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_370),
.B(n_181),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_335),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_337),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_338),
.B(n_269),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_342),
.B(n_176),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_342),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_345),
.Y(n_451)
);

BUFx8_ASAP7_75t_SL g452 ( 
.A(n_384),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_292),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_426),
.B(n_251),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_397),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_424),
.B(n_296),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_397),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_385),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_297),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_418),
.A2(n_309),
.B1(n_300),
.B2(n_323),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_303),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_310),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_393),
.A2(n_341),
.B1(n_375),
.B2(n_368),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_397),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_414),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_445),
.A2(n_234),
.B1(n_205),
.B2(n_293),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_433),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_359),
.C(n_355),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

OAI22xp33_ASAP7_75t_L g475 ( 
.A1(n_393),
.A2(n_199),
.B1(n_356),
.B2(n_254),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_408),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_418),
.A2(n_282),
.B1(n_276),
.B2(n_253),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_417),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_383),
.Y(n_479)
);

NOR2x1p5_ASAP7_75t_L g480 ( 
.A(n_429),
.B(n_264),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_384),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_388),
.B(n_311),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_445),
.A2(n_180),
.B1(n_183),
.B2(n_188),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_412),
.B(n_243),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_388),
.B(n_317),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_426),
.B(n_430),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_417),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_418),
.A2(n_251),
.B1(n_325),
.B2(n_370),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_426),
.B(n_326),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_426),
.B(n_329),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_424),
.B(n_332),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_402),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_426),
.B(n_336),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_430),
.B(n_340),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_424),
.B(n_344),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_392),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_435),
.B(n_346),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_418),
.B(n_348),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_392),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_418),
.A2(n_251),
.B1(n_371),
.B2(n_372),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_429),
.B(n_444),
.C(n_437),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_418),
.A2(n_251),
.B1(n_371),
.B2(n_372),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_412),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_385),
.B(n_350),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

BUFx6f_ASAP7_75t_SL g518 ( 
.A(n_412),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_385),
.B(n_352),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_412),
.B(n_182),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_435),
.B(n_365),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_435),
.B(n_438),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_483),
.B(n_412),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_487),
.B(n_405),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_501),
.B(n_405),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_471),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_459),
.B(n_490),
.Y(n_529)
);

NAND3xp33_ASAP7_75t_SL g530 ( 
.A(n_469),
.B(n_339),
.C(n_485),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_405),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_369),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_510),
.B(n_422),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_405),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_461),
.B(n_453),
.C(n_472),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_464),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_376),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_493),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_493),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_493),
.B(n_422),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_468),
.B(n_405),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_513),
.B(n_520),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_468),
.B(n_478),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_478),
.B(n_415),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_513),
.B(n_422),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_513),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_466),
.B(n_433),
.C(n_404),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_491),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_498),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_471),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_498),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_469),
.B(n_380),
.C(n_379),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_460),
.B(n_198),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_463),
.B(n_422),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_454),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_470),
.B(n_294),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_471),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_477),
.B(n_381),
.C(n_437),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_505),
.B(n_444),
.C(n_404),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_521),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_456),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_473),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_465),
.B(n_415),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_495),
.A2(n_438),
.B(n_415),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_499),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_499),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_514),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_500),
.B(n_422),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_486),
.B(n_422),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_520),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_514),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_457),
.B(n_394),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_518),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_486),
.B(n_480),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_486),
.B(n_520),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_520),
.B(n_387),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_486),
.B(n_415),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_480),
.B(n_419),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_516),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_522),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_497),
.B(n_295),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_494),
.B(n_419),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_522),
.A2(n_438),
.B1(n_415),
.B2(n_387),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_522),
.A2(n_387),
.B1(n_407),
.B2(n_406),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_516),
.B(n_408),
.Y(n_589)
);

NOR2x1p5_ASAP7_75t_L g590 ( 
.A(n_470),
.B(n_183),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_496),
.A2(n_522),
.B1(n_518),
.B2(n_502),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_522),
.A2(n_328),
.B1(n_330),
.B2(n_312),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_509),
.B(n_419),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_473),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_517),
.B(n_387),
.Y(n_595)
);

NAND2x1_ASAP7_75t_L g596 ( 
.A(n_455),
.B(n_382),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_479),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_517),
.B(n_408),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_511),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_512),
.B(n_408),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_458),
.B(n_408),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_458),
.B(n_408),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_458),
.B(n_387),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_511),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_475),
.B(n_406),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_479),
.B(n_406),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_518),
.A2(n_387),
.B1(n_416),
.B2(n_406),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_458),
.B(n_407),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_492),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_492),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_504),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_504),
.B(n_407),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_467),
.B(n_407),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_452),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_507),
.B(n_508),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_507),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_455),
.B(n_200),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_485),
.B(n_411),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_535),
.A2(n_301),
.B1(n_299),
.B2(n_518),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_525),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_529),
.A2(n_489),
.B(n_476),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_579),
.A2(n_489),
.B(n_476),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_602),
.A2(n_474),
.B(n_467),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_576),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_603),
.A2(n_474),
.B(n_467),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_579),
.A2(n_581),
.B(n_523),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_578),
.A2(n_455),
.B1(n_489),
.B2(n_476),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_606),
.A2(n_544),
.B(n_531),
.C(n_548),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_567),
.A2(n_489),
.B(n_476),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_568),
.A2(n_508),
.B(n_507),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_574),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_532),
.B(n_508),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_601),
.A2(n_474),
.B(n_467),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_525),
.Y(n_637)
);

AOI21x1_ASAP7_75t_L g638 ( 
.A1(n_618),
.A2(n_416),
.B(n_395),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_537),
.A2(n_411),
.B(n_425),
.C(n_247),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_587),
.A2(n_484),
.B(n_474),
.Y(n_641)
);

NOR2x1p5_ASAP7_75t_SL g642 ( 
.A(n_552),
.B(n_560),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_604),
.A2(n_481),
.B(n_456),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_564),
.B(n_543),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_536),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_540),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_551),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_574),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_SL g649 ( 
.A1(n_606),
.A2(n_283),
.B(n_286),
.C(n_281),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_552),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_527),
.A2(n_488),
.B(n_484),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_524),
.A2(n_488),
.B(n_484),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_543),
.B(n_427),
.Y(n_653)
);

AND2x4_ASAP7_75t_SL g654 ( 
.A(n_540),
.B(n_425),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_560),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_534),
.A2(n_488),
.B(n_484),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_553),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_617),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_582),
.B(n_358),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_543),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_586),
.B(n_488),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_562),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_L g663 ( 
.A(n_584),
.B(n_455),
.Y(n_663)
);

BUFx8_ASAP7_75t_L g664 ( 
.A(n_582),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_526),
.B(n_361),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_550),
.A2(n_586),
.B(n_584),
.C(n_538),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_539),
.A2(n_455),
.B1(n_209),
.B2(n_212),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_547),
.A2(n_427),
.B(n_441),
.C(n_442),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_588),
.A2(n_503),
.B(n_416),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_556),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_593),
.B(n_569),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_542),
.A2(n_455),
.B(n_503),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_528),
.A2(n_503),
.B(n_416),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_593),
.A2(n_427),
.B(n_443),
.C(n_442),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_570),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_580),
.A2(n_455),
.B1(n_230),
.B2(n_248),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_562),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_559),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_595),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_571),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_575),
.B(n_503),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_583),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_558),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_545),
.B(n_456),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_540),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_595),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_566),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_561),
.B(n_185),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_595),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_566),
.B(n_456),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_580),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_621),
.B(n_185),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_580),
.A2(n_272),
.B1(n_249),
.B2(n_449),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_592),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_591),
.A2(n_186),
.B1(n_189),
.B2(n_193),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_573),
.A2(n_481),
.B(n_456),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_SL g697 ( 
.A(n_617),
.B(n_187),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_573),
.A2(n_481),
.B(n_462),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_556),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_594),
.B(n_597),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_594),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_597),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_563),
.B(n_391),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_599),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_609),
.A2(n_481),
.B(n_462),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_616),
.A2(n_481),
.B(n_462),
.Y(n_706)
);

AOI21xp33_ASAP7_75t_L g707 ( 
.A1(n_554),
.A2(n_265),
.B(n_188),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_599),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_598),
.A2(n_481),
.B(n_462),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_530),
.B(n_186),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_557),
.A2(n_462),
.B(n_401),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_557),
.A2(n_462),
.B(n_401),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_610),
.B(n_619),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_556),
.A2(n_401),
.B(n_400),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_549),
.B(n_585),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_608),
.A2(n_284),
.B1(n_189),
.B2(n_193),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_556),
.B(n_270),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_572),
.A2(n_401),
.B(n_400),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_590),
.B(n_391),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_565),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_610),
.B(n_391),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_555),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_577),
.B(n_446),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_618),
.A2(n_449),
.B(n_395),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_619),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_533),
.A2(n_443),
.B(n_441),
.C(n_449),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_572),
.A2(n_401),
.B(n_400),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_629),
.A2(n_589),
.B(n_600),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_658),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_653),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_653),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_627),
.B(n_577),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_629),
.A2(n_565),
.B(n_546),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_650),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_R g735 ( 
.A(n_646),
.B(n_577),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_635),
.A2(n_565),
.B(n_546),
.Y(n_736)
);

BUFx2_ASAP7_75t_SL g737 ( 
.A(n_670),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_692),
.A2(n_533),
.B(n_541),
.C(n_605),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_634),
.B(n_565),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_655),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_701),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_683),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_624),
.A2(n_541),
.B(n_620),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_662),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_677),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_659),
.B(n_555),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_660),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_644),
.Y(n_748)
);

OAI21xp33_ASAP7_75t_SL g749 ( 
.A1(n_647),
.A2(n_589),
.B(n_611),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_670),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_685),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_624),
.A2(n_620),
.B(n_614),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_665),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_704),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_632),
.A2(n_625),
.B(n_643),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_634),
.B(n_612),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_710),
.A2(n_555),
.B1(n_615),
.B2(n_613),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_694),
.A2(n_689),
.B1(n_686),
.B2(n_691),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_679),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_670),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_634),
.B(n_270),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_SL g762 ( 
.A1(n_661),
.A2(n_614),
.B(n_607),
.C(n_596),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_708),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_671),
.B(n_555),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_678),
.B(n_607),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_664),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_648),
.B(n_273),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_648),
.B(n_273),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_632),
.A2(n_401),
.B(n_400),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_703),
.B(n_555),
.Y(n_770)
);

AOI21x1_ASAP7_75t_L g771 ( 
.A1(n_633),
.A2(n_395),
.B(n_390),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_707),
.B(n_275),
.C(n_271),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_625),
.A2(n_401),
.B(n_400),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_648),
.B(n_660),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_719),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_623),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_622),
.B(n_271),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_679),
.B(n_274),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_691),
.B(n_555),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_657),
.B(n_434),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_640),
.A2(n_377),
.B(n_378),
.C(n_447),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_687),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_675),
.B(n_274),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_664),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_684),
.A2(n_663),
.B(n_641),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_699),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_641),
.A2(n_401),
.B(n_400),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_725),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_631),
.A2(n_669),
.B(n_633),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_669),
.A2(n_400),
.B(n_386),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_696),
.A2(n_400),
.B(n_386),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_699),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_680),
.B(n_279),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_R g794 ( 
.A(n_715),
.B(n_279),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_682),
.B(n_447),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_639),
.B(n_447),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_755),
.A2(n_696),
.B(n_656),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_777),
.A2(n_666),
.B(n_674),
.C(n_668),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_769),
.A2(n_628),
.B(n_626),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_741),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_743),
.A2(n_785),
.B(n_733),
.Y(n_801)
);

OAI21x1_ASAP7_75t_SL g802 ( 
.A1(n_746),
.A2(n_726),
.B(n_698),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_753),
.B(n_654),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_775),
.A2(n_697),
.B1(n_695),
.B2(n_693),
.Y(n_804)
);

AO31x2_ASAP7_75t_L g805 ( 
.A1(n_738),
.A2(n_727),
.A3(n_718),
.B(n_722),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_729),
.B(n_717),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_789),
.A2(n_736),
.B(n_752),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_761),
.A2(n_688),
.B1(n_716),
.B2(n_637),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_750),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_796),
.B(n_645),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_741),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_754),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_728),
.A2(n_656),
.B(n_652),
.Y(n_813)
);

OR2x6_ASAP7_75t_L g814 ( 
.A(n_737),
.B(n_723),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_760),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_794),
.B(n_630),
.Y(n_816)
);

AO21x1_ASAP7_75t_L g817 ( 
.A1(n_770),
.A2(n_718),
.B(n_727),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_796),
.B(n_721),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_781),
.A2(n_642),
.B(n_698),
.C(n_652),
.Y(n_819)
);

BUFx4_ASAP7_75t_SL g820 ( 
.A(n_766),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_SL g821 ( 
.A1(n_779),
.A2(n_723),
.B(n_672),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_767),
.A2(n_676),
.B1(n_667),
.B2(n_288),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_758),
.A2(n_700),
.B1(n_713),
.B2(n_702),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_730),
.B(n_731),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_787),
.A2(n_638),
.B(n_636),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_734),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_773),
.A2(n_636),
.B(n_651),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_742),
.B(n_649),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_754),
.Y(n_829)
);

AO32x2_ASAP7_75t_L g830 ( 
.A1(n_760),
.A2(n_651),
.A3(n_724),
.B1(n_712),
.B2(n_711),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_763),
.B(n_720),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_730),
.B(n_232),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_791),
.A2(n_712),
.B(n_711),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_750),
.Y(n_834)
);

AO31x2_ASAP7_75t_L g835 ( 
.A1(n_764),
.A2(n_673),
.A3(n_709),
.B(n_706),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_790),
.A2(n_706),
.B(n_705),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_757),
.A2(n_673),
.B(n_681),
.C(n_709),
.Y(n_837)
);

AO32x2_ASAP7_75t_L g838 ( 
.A1(n_760),
.A2(n_705),
.A3(n_259),
.B1(n_690),
.B2(n_720),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_734),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_731),
.B(n_259),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_763),
.B(n_714),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_788),
.Y(n_842)
);

OAI21x1_ASAP7_75t_SL g843 ( 
.A1(n_788),
.A2(n_396),
.B(n_389),
.Y(n_843)
);

OA21x2_ASAP7_75t_L g844 ( 
.A1(n_771),
.A2(n_398),
.B(n_390),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_776),
.B(n_446),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_771),
.A2(n_396),
.B(n_389),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_740),
.Y(n_847)
);

AO31x2_ASAP7_75t_L g848 ( 
.A1(n_740),
.A2(n_398),
.A3(n_399),
.B(n_403),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_765),
.B(n_446),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_765),
.B(n_446),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_759),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_744),
.Y(n_852)
);

AO31x2_ASAP7_75t_L g853 ( 
.A1(n_744),
.A2(n_745),
.A3(n_782),
.B(n_792),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_SL g854 ( 
.A1(n_732),
.A2(n_409),
.B(n_390),
.C(n_398),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_745),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_782),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_729),
.B(n_63),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_853),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_816),
.A2(n_772),
.B1(n_748),
.B2(n_793),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_853),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_809),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_804),
.A2(n_783),
.B1(n_778),
.B2(n_768),
.Y(n_862)
);

CKINVDCx6p67_ASAP7_75t_R g863 ( 
.A(n_803),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_809),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_844),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_844),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_824),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_835),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_832),
.A2(n_779),
.B1(n_780),
.B2(n_784),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_824),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_SL g871 ( 
.A1(n_806),
.A2(n_766),
.B1(n_735),
.B2(n_779),
.Y(n_871)
);

INVx6_ASAP7_75t_L g872 ( 
.A(n_809),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_835),
.Y(n_873)
);

BUFx12f_ASAP7_75t_L g874 ( 
.A(n_840),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_853),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_806),
.A2(n_780),
.B1(n_759),
.B2(n_187),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_800),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_808),
.A2(n_747),
.B1(n_751),
.B2(n_780),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_830),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_828),
.A2(n_759),
.B1(n_187),
.B2(n_795),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_810),
.B(n_751),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_818),
.A2(n_747),
.B1(n_756),
.B2(n_774),
.Y(n_883)
);

BUFx4f_ASAP7_75t_SL g884 ( 
.A(n_834),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_818),
.A2(n_792),
.B1(n_786),
.B2(n_259),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_812),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_822),
.A2(n_786),
.B1(n_374),
.B2(n_739),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_810),
.A2(n_275),
.B1(n_289),
.B2(n_285),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_830),
.Y(n_889)
);

BUFx8_ASAP7_75t_SL g890 ( 
.A(n_820),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_829),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_834),
.Y(n_892)
);

CKINVDCx6p67_ASAP7_75t_R g893 ( 
.A(n_834),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_849),
.B(n_850),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_815),
.Y(n_895)
);

BUFx2_ASAP7_75t_SL g896 ( 
.A(n_815),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_814),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_842),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_831),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_SL g900 ( 
.A1(n_823),
.A2(n_289),
.B1(n_285),
.B2(n_802),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_830),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_849),
.A2(n_749),
.B1(n_287),
.B2(n_280),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_850),
.A2(n_280),
.B1(n_288),
.B2(n_287),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_826),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_851),
.A2(n_284),
.B1(n_378),
.B2(n_377),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_827),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_851),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_798),
.A2(n_421),
.B1(n_420),
.B2(n_439),
.Y(n_908)
);

OAI22xp33_ASAP7_75t_L g909 ( 
.A1(n_857),
.A2(n_841),
.B1(n_814),
.B2(n_831),
.Y(n_909)
);

INVx6_ASAP7_75t_L g910 ( 
.A(n_814),
.Y(n_910)
);

CKINVDCx11_ASAP7_75t_R g911 ( 
.A(n_839),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_847),
.A2(n_750),
.B1(n_737),
.B2(n_345),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_852),
.B(n_750),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_855),
.A2(n_856),
.B1(n_841),
.B2(n_823),
.Y(n_914)
);

OAI22xp33_ASAP7_75t_L g915 ( 
.A1(n_845),
.A2(n_750),
.B1(n_420),
.B2(n_421),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_848),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_843),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_817),
.A2(n_434),
.B1(n_451),
.B2(n_436),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_819),
.A2(n_436),
.B1(n_451),
.B2(n_434),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_858),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_865),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_858),
.Y(n_922)
);

OA21x2_ASAP7_75t_L g923 ( 
.A1(n_916),
.A2(n_807),
.B(n_797),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_897),
.B(n_807),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_860),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_868),
.Y(n_926)
);

NOR2x1_ASAP7_75t_SL g927 ( 
.A(n_896),
.B(n_846),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_910),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_865),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_860),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_875),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_862),
.A2(n_845),
.B1(n_837),
.B2(n_821),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_875),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_916),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_859),
.A2(n_451),
.B1(n_436),
.B2(n_439),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_910),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_866),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_910),
.Y(n_939)
);

OAI22xp33_ASAP7_75t_L g940 ( 
.A1(n_874),
.A2(n_813),
.B1(n_801),
.B2(n_797),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_866),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_900),
.A2(n_439),
.B1(n_813),
.B2(n_413),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_866),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_877),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_868),
.A2(n_836),
.B(n_833),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_899),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_897),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_868),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_877),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_879),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_879),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_919),
.A2(n_799),
.B(n_825),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_868),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_886),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_880),
.B(n_805),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_880),
.B(n_838),
.Y(n_956)
);

AO31x2_ASAP7_75t_L g957 ( 
.A1(n_880),
.A2(n_838),
.A3(n_805),
.B(n_835),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_886),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_944),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_937),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_947),
.B(n_867),
.Y(n_961)
);

AOI211xp5_ASAP7_75t_L g962 ( 
.A1(n_940),
.A2(n_909),
.B(n_878),
.C(n_882),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_946),
.B(n_894),
.Y(n_963)
);

O2A1O1Ixp5_ASAP7_75t_L g964 ( 
.A1(n_932),
.A2(n_914),
.B(n_873),
.C(n_906),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_932),
.A2(n_876),
.B(n_881),
.C(n_902),
.Y(n_965)
);

NOR2x1_ASAP7_75t_SL g966 ( 
.A(n_928),
.B(n_896),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_942),
.A2(n_908),
.B(n_871),
.C(n_887),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_956),
.B(n_889),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_956),
.B(n_889),
.Y(n_969)
);

AO32x1_ASAP7_75t_L g970 ( 
.A1(n_922),
.A2(n_901),
.A3(n_889),
.B1(n_906),
.B2(n_898),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_946),
.B(n_873),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_924),
.B(n_937),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_944),
.B(n_891),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_947),
.B(n_867),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_SL g975 ( 
.A1(n_937),
.A2(n_895),
.B(n_898),
.C(n_891),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_942),
.A2(n_908),
.B(n_903),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_L g977 ( 
.A1(n_935),
.A2(n_888),
.B1(n_885),
.B2(n_869),
.C(n_905),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_935),
.A2(n_863),
.B1(n_874),
.B2(n_883),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_949),
.Y(n_979)
);

INVx5_ASAP7_75t_SL g980 ( 
.A(n_924),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_956),
.B(n_901),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_923),
.A2(n_915),
.B(n_906),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_949),
.B(n_901),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_924),
.A2(n_863),
.B1(n_911),
.B2(n_910),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_958),
.B(n_904),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_928),
.B(n_939),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_928),
.B(n_870),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_950),
.B(n_873),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_950),
.B(n_873),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_L g990 ( 
.A1(n_924),
.A2(n_917),
.B(n_918),
.Y(n_990)
);

AOI221xp5_ASAP7_75t_L g991 ( 
.A1(n_951),
.A2(n_854),
.B1(n_917),
.B2(n_870),
.C(n_913),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_939),
.B(n_870),
.Y(n_992)
);

AND2x4_ASAP7_75t_SL g993 ( 
.A(n_951),
.B(n_897),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_954),
.B(n_838),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_939),
.A2(n_917),
.B1(n_897),
.B2(n_912),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_954),
.B(n_907),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_958),
.B(n_907),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_936),
.B(n_897),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_934),
.B(n_864),
.Y(n_999)
);

NOR2x1_ASAP7_75t_R g1000 ( 
.A(n_960),
.B(n_890),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_959),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_970),
.Y(n_1002)
);

INVx3_ASAP7_75t_SL g1003 ( 
.A(n_972),
.Y(n_1003)
);

AND2x2_ASAP7_75t_SL g1004 ( 
.A(n_993),
.B(n_923),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_979),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_983),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_983),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_973),
.Y(n_1008)
);

NOR2xp67_ASAP7_75t_L g1009 ( 
.A(n_984),
.B(n_921),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_989),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_968),
.B(n_969),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_970),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_968),
.B(n_957),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_970),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_960),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_969),
.B(n_957),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_963),
.B(n_934),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_981),
.B(n_957),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_981),
.B(n_955),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_972),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_978),
.B(n_955),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_970),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_994),
.B(n_957),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_971),
.B(n_957),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_988),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_1021),
.A2(n_967),
.B(n_976),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_1025),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1011),
.B(n_972),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1001),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_1021),
.A2(n_967),
.B1(n_977),
.B2(n_965),
.C(n_962),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1011),
.B(n_972),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1011),
.B(n_980),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1008),
.A2(n_965),
.B1(n_964),
.B2(n_990),
.C(n_1017),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1001),
.Y(n_1034)
);

OAI33xp33_ASAP7_75t_L g1035 ( 
.A1(n_1017),
.A2(n_1008),
.A3(n_1002),
.B1(n_1022),
.B2(n_1014),
.B3(n_1025),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1009),
.A2(n_995),
.B1(n_991),
.B2(n_985),
.Y(n_1036)
);

AO21x2_ASAP7_75t_L g1037 ( 
.A1(n_1002),
.A2(n_982),
.B(n_975),
.Y(n_1037)
);

AOI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_1002),
.A2(n_1014),
.B1(n_1022),
.B2(n_1012),
.C(n_1023),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_1019),
.B(n_994),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_1020),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_1000),
.B(n_986),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1019),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_1020),
.B(n_999),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_L g1044 ( 
.A(n_1009),
.B(n_986),
.C(n_997),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1001),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1015),
.A2(n_992),
.B1(n_987),
.B2(n_980),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_1020),
.B(n_999),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_1020),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1043),
.B(n_1020),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1045),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1033),
.B(n_1006),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1042),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1029),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1033),
.B(n_1006),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1029),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1031),
.B(n_1003),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1034),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1052),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1051),
.B(n_1039),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1053),
.B(n_1057),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_1055),
.B(n_1039),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1052),
.B(n_1038),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1053),
.B(n_1043),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1054),
.B(n_1038),
.Y(n_1066)
);

AOI21xp33_ASAP7_75t_SL g1067 ( 
.A1(n_1057),
.A2(n_1026),
.B(n_1041),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1067),
.B(n_1026),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1061),
.B(n_1063),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_1064),
.B(n_1058),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1062),
.B(n_1058),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1064),
.B(n_1027),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1071),
.B(n_1065),
.Y(n_1073)
);

AOI211xp5_ASAP7_75t_L g1074 ( 
.A1(n_1068),
.A2(n_1030),
.B(n_1036),
.C(n_1066),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_1072),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1070),
.A2(n_1030),
.B1(n_1069),
.B2(n_1066),
.Y(n_1076)
);

OAI21xp33_ASAP7_75t_SL g1077 ( 
.A1(n_1068),
.A2(n_1060),
.B(n_1032),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1072),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1071),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1072),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1068),
.A2(n_1046),
.B1(n_1048),
.B2(n_1049),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1068),
.B(n_1044),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_1068),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1068),
.A2(n_1015),
.B(n_1012),
.C(n_1040),
.Y(n_1084)
);

NAND2x1_ASAP7_75t_L g1085 ( 
.A(n_1079),
.B(n_1048),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1074),
.B(n_1054),
.Y(n_1086)
);

AOI221xp5_ASAP7_75t_L g1087 ( 
.A1(n_1083),
.A2(n_1035),
.B1(n_1056),
.B2(n_1059),
.C(n_1037),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1079),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1075),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1073),
.B(n_1048),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1078),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1076),
.A2(n_1012),
.B1(n_1010),
.B2(n_1015),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1082),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1080),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1076),
.B(n_1048),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1081),
.Y(n_1096)
);

XOR2x2_ASAP7_75t_L g1097 ( 
.A(n_1077),
.B(n_1000),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1084),
.B(n_1031),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1084),
.B(n_1056),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_1079),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_1075),
.B(n_1015),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1095),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1101),
.A2(n_1096),
.B1(n_1097),
.B2(n_1089),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1100),
.B(n_1049),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1088),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1093),
.B(n_1094),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1091),
.Y(n_1107)
);

AOI222xp33_ASAP7_75t_L g1108 ( 
.A1(n_1086),
.A2(n_1012),
.B1(n_1059),
.B2(n_1023),
.C1(n_1050),
.C2(n_1049),
.Y(n_1108)
);

OAI221xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1087),
.A2(n_1040),
.B1(n_1032),
.B2(n_1010),
.C(n_1050),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1086),
.A2(n_1040),
.B(n_1050),
.C(n_1049),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1085),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1099),
.Y(n_1112)
);

OA21x2_ASAP7_75t_L g1113 ( 
.A1(n_1099),
.A2(n_1045),
.B(n_1034),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_1092),
.Y(n_1114)
);

XNOR2xp5_ASAP7_75t_L g1115 ( 
.A(n_1092),
.B(n_10),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1090),
.A2(n_1037),
.B1(n_1040),
.B2(n_1003),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_SL g1117 ( 
.A1(n_1098),
.A2(n_1045),
.B(n_1024),
.C(n_12),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1100),
.B(n_1043),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1100),
.B(n_1037),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1101),
.B(n_1047),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1086),
.A2(n_1037),
.B(n_975),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1103),
.B(n_1047),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1106),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1115),
.B(n_1047),
.Y(n_1124)
);

AO22x1_ASAP7_75t_L g1125 ( 
.A1(n_1102),
.A2(n_1047),
.B1(n_892),
.B2(n_864),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1111),
.B(n_1007),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_SL g1127 ( 
.A(n_1107),
.B(n_413),
.C(n_10),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1114),
.B(n_1007),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1112),
.A2(n_966),
.B(n_927),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1117),
.A2(n_927),
.B(n_998),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1105),
.B(n_1007),
.Y(n_1131)
);

AND3x2_ASAP7_75t_L g1132 ( 
.A(n_1104),
.B(n_11),
.C(n_14),
.Y(n_1132)
);

OAI221xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1121),
.A2(n_1024),
.B1(n_1023),
.B2(n_16),
.C(n_17),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1118),
.B(n_1007),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1110),
.B(n_1001),
.Y(n_1135)
);

NOR3x1_ASAP7_75t_L g1136 ( 
.A(n_1120),
.B(n_861),
.C(n_1024),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1119),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1113),
.Y(n_1138)
);

OAI221xp5_ASAP7_75t_L g1139 ( 
.A1(n_1133),
.A2(n_1109),
.B1(n_1108),
.B2(n_1116),
.C(n_1113),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1122),
.A2(n_1108),
.B1(n_980),
.B2(n_1004),
.Y(n_1140)
);

AOI211xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1133),
.A2(n_884),
.B(n_15),
.C(n_18),
.Y(n_1141)
);

OAI222xp33_ASAP7_75t_L g1142 ( 
.A1(n_1138),
.A2(n_1019),
.B1(n_961),
.B2(n_974),
.C1(n_1005),
.C2(n_999),
.Y(n_1142)
);

AOI211xp5_ASAP7_75t_L g1143 ( 
.A1(n_1123),
.A2(n_1124),
.B(n_1137),
.C(n_1128),
.Y(n_1143)
);

AOI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1131),
.A2(n_14),
.B(n_15),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1127),
.A2(n_1004),
.B1(n_1005),
.B2(n_993),
.Y(n_1145)
);

OAI211xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1135),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_L g1147 ( 
.A(n_1136),
.B(n_864),
.C(n_23),
.D(n_24),
.Y(n_1147)
);

NAND2xp33_ASAP7_75t_L g1148 ( 
.A(n_1126),
.B(n_892),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1132),
.B(n_1005),
.Y(n_1149)
);

AOI21xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1125),
.A2(n_20),
.B(n_23),
.Y(n_1150)
);

AOI211xp5_ASAP7_75t_L g1151 ( 
.A1(n_1129),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1134),
.A2(n_1004),
.B1(n_1005),
.B2(n_1013),
.Y(n_1152)
);

AOI32xp33_ASAP7_75t_L g1153 ( 
.A1(n_1130),
.A2(n_1018),
.A3(n_1016),
.B1(n_1013),
.B2(n_996),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1132),
.B(n_26),
.Y(n_1154)
);

OAI211xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1123),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1132),
.Y(n_1156)
);

OAI21xp33_ASAP7_75t_SL g1157 ( 
.A1(n_1138),
.A2(n_1004),
.B(n_1016),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_L g1158 ( 
.A1(n_1133),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.C(n_35),
.Y(n_1158)
);

OAI211xp5_ASAP7_75t_SL g1159 ( 
.A1(n_1123),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1122),
.A2(n_872),
.B1(n_1016),
.B2(n_1013),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_R g1161 ( 
.A(n_1132),
.B(n_36),
.Y(n_1161)
);

AOI221xp5_ASAP7_75t_L g1162 ( 
.A1(n_1133),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.C(n_40),
.Y(n_1162)
);

AOI322xp5_ASAP7_75t_L g1163 ( 
.A1(n_1156),
.A2(n_1018),
.A3(n_930),
.B1(n_920),
.B2(n_933),
.C1(n_925),
.C2(n_922),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1140),
.A2(n_872),
.B1(n_925),
.B2(n_931),
.Y(n_1164)
);

OAI211xp5_ASAP7_75t_L g1165 ( 
.A1(n_1161),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1165)
);

AOI222xp33_ASAP7_75t_L g1166 ( 
.A1(n_1139),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.C1(n_44),
.C2(n_45),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1158),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.C(n_46),
.Y(n_1167)
);

OAI22xp33_ASAP7_75t_R g1168 ( 
.A1(n_1143),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_1168)
);

OAI321xp33_ASAP7_75t_L g1169 ( 
.A1(n_1147),
.A2(n_861),
.A3(n_892),
.B1(n_895),
.B2(n_53),
.C(n_56),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1162),
.A2(n_893),
.B1(n_872),
.B2(n_864),
.Y(n_1170)
);

NAND5xp2_ASAP7_75t_L g1171 ( 
.A(n_1141),
.B(n_47),
.C(n_51),
.D(n_52),
.E(n_53),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1154),
.B(n_52),
.Y(n_1172)
);

NOR4xp75_ASAP7_75t_L g1173 ( 
.A(n_1149),
.B(n_56),
.C(n_57),
.D(n_59),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1146),
.A2(n_1159),
.B(n_1155),
.C(n_1144),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_1151),
.B(n_892),
.C(n_60),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1160),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_L g1177 ( 
.A(n_1150),
.B(n_423),
.C(n_440),
.Y(n_1177)
);

AOI222xp33_ASAP7_75t_L g1178 ( 
.A1(n_1148),
.A2(n_57),
.B1(n_1018),
.B2(n_933),
.C1(n_931),
.C2(n_872),
.Y(n_1178)
);

NOR4xp25_ASAP7_75t_L g1179 ( 
.A(n_1157),
.B(n_423),
.C(n_431),
.D(n_440),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1145),
.A2(n_1152),
.B1(n_1153),
.B2(n_1142),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1161),
.B(n_440),
.C(n_431),
.Y(n_1181)
);

AOI211xp5_ASAP7_75t_L g1182 ( 
.A1(n_1158),
.A2(n_892),
.B(n_431),
.C(n_423),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1141),
.A2(n_762),
.B(n_431),
.C(n_440),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1161),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_L g1185 ( 
.A(n_1156),
.B(n_423),
.C(n_446),
.Y(n_1185)
);

AOI211xp5_ASAP7_75t_L g1186 ( 
.A1(n_1158),
.A2(n_410),
.B(n_403),
.C(n_409),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1184),
.A2(n_1176),
.B1(n_1164),
.B2(n_1175),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_L g1188 ( 
.A(n_1165),
.B(n_410),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1173),
.B(n_920),
.Y(n_1189)
);

XNOR2xp5_ASAP7_75t_L g1190 ( 
.A(n_1170),
.B(n_65),
.Y(n_1190)
);

NOR3xp33_ASAP7_75t_L g1191 ( 
.A(n_1181),
.B(n_409),
.C(n_403),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1172),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1167),
.B(n_893),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_SL g1194 ( 
.A(n_1171),
.B(n_399),
.C(n_71),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_1168),
.B(n_432),
.Y(n_1195)
);

NOR2x1_ASAP7_75t_L g1196 ( 
.A(n_1183),
.B(n_1174),
.Y(n_1196)
);

NAND4xp75_ASAP7_75t_L g1197 ( 
.A(n_1180),
.B(n_399),
.C(n_923),
.D(n_75),
.Y(n_1197)
);

NAND4xp75_ASAP7_75t_L g1198 ( 
.A(n_1166),
.B(n_923),
.C(n_73),
.D(n_77),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1170),
.A2(n_1169),
.B1(n_1178),
.B2(n_1163),
.Y(n_1199)
);

XOR2x1_ASAP7_75t_L g1200 ( 
.A(n_1177),
.B(n_70),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1185),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1182),
.B(n_78),
.Y(n_1202)
);

NOR2xp67_ASAP7_75t_L g1203 ( 
.A(n_1179),
.B(n_80),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1186),
.B(n_957),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1184),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1172),
.B(n_432),
.Y(n_1206)
);

AND2x2_ASAP7_75t_SL g1207 ( 
.A(n_1184),
.B(n_432),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1184),
.B(n_930),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1205),
.A2(n_432),
.B(n_448),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1189),
.B(n_83),
.Y(n_1210)
);

NAND4xp75_ASAP7_75t_L g1211 ( 
.A(n_1196),
.B(n_84),
.C(n_89),
.D(n_90),
.Y(n_1211)
);

OAI221xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1187),
.A2(n_938),
.B1(n_936),
.B2(n_943),
.C(n_941),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1189),
.B(n_432),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1188),
.B(n_432),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1195),
.B(n_1192),
.Y(n_1215)
);

OAI221xp5_ASAP7_75t_L g1216 ( 
.A1(n_1199),
.A2(n_923),
.B1(n_941),
.B2(n_943),
.C(n_938),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1194),
.A2(n_948),
.B(n_953),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1193),
.B(n_450),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1200),
.B(n_92),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1203),
.A2(n_945),
.B(n_953),
.C(n_926),
.Y(n_1220)
);

NAND2x1_ASAP7_75t_L g1221 ( 
.A(n_1201),
.B(n_1208),
.Y(n_1221)
);

OAI211xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1202),
.A2(n_94),
.B(n_96),
.C(n_97),
.Y(n_1222)
);

OR3x2_ASAP7_75t_L g1223 ( 
.A(n_1204),
.B(n_99),
.C(n_102),
.Y(n_1223)
);

AOI22x1_ASAP7_75t_L g1224 ( 
.A1(n_1210),
.A2(n_1190),
.B1(n_1206),
.B2(n_1207),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1217),
.A2(n_1191),
.B(n_1197),
.C(n_1198),
.Y(n_1225)
);

AOI221xp5_ASAP7_75t_L g1226 ( 
.A1(n_1212),
.A2(n_432),
.B1(n_448),
.B2(n_450),
.C(n_948),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1213),
.B(n_1218),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_SL g1228 ( 
.A(n_1215),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1214),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1211),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1219),
.B(n_450),
.Y(n_1231)
);

OAI21xp33_ASAP7_75t_L g1232 ( 
.A1(n_1221),
.A2(n_953),
.B(n_926),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1223),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1222),
.A2(n_926),
.B1(n_929),
.B2(n_921),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1209),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1220),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1216),
.B(n_105),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1210),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1228),
.A2(n_926),
.B1(n_450),
.B2(n_432),
.Y(n_1239)
);

AO22x2_ASAP7_75t_L g1240 ( 
.A1(n_1229),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_1240)
);

AOI211xp5_ASAP7_75t_L g1241 ( 
.A1(n_1237),
.A2(n_450),
.B(n_448),
.C(n_115),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1238),
.Y(n_1242)
);

OAI22x1_ASAP7_75t_L g1243 ( 
.A1(n_1224),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1227),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1233),
.A2(n_450),
.B1(n_448),
.B2(n_921),
.Y(n_1245)
);

OAI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1230),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1236),
.A2(n_450),
.B1(n_448),
.B2(n_929),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1225),
.A2(n_929),
.B1(n_952),
.B2(n_450),
.Y(n_1248)
);

OAI22x1_ASAP7_75t_L g1249 ( 
.A1(n_1242),
.A2(n_1235),
.B1(n_1231),
.B2(n_1234),
.Y(n_1249)
);

OAI22x1_ASAP7_75t_L g1250 ( 
.A1(n_1244),
.A2(n_1235),
.B1(n_1232),
.B2(n_1226),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1240),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1243),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1246),
.A2(n_448),
.B1(n_133),
.B2(n_137),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1240),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1252),
.B(n_1248),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1251),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1254),
.A2(n_1239),
.B1(n_1245),
.B2(n_1241),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1253),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1256),
.A2(n_1247),
.B1(n_1249),
.B2(n_1250),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1259),
.A2(n_1255),
.B(n_1257),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1260),
.A2(n_1258),
.B(n_138),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1261),
.Y(n_1262)
);

AOI221xp5_ASAP7_75t_L g1263 ( 
.A1(n_1262),
.A2(n_448),
.B1(n_386),
.B2(n_382),
.C(n_145),
.Y(n_1263)
);

AOI211xp5_ASAP7_75t_L g1264 ( 
.A1(n_1263),
.A2(n_448),
.B(n_141),
.C(n_142),
.Y(n_1264)
);


endmodule