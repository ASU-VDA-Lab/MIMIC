module fake_jpeg_2407_n_216 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_55),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_67),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_91),
.Y(n_99)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_81),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_71),
.B1(n_58),
.B2(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_82),
.B1(n_79),
.B2(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_104),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_111),
.B1(n_88),
.B2(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_65),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_82),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_79),
.B1(n_71),
.B2(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_116),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_62),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_123),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_96),
.B(n_68),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_137),
.B(n_5),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_0),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_62),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_132),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_59),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_136),
.B1(n_21),
.B2(n_52),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_60),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_61),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_58),
.B1(n_72),
.B2(n_77),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_77),
.B(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_142),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_147),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_64),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_24),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_146),
.C(n_9),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_25),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_0),
.C(n_1),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_26),
.B1(n_51),
.B2(n_50),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_2),
.B(n_3),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_11),
.B(n_12),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_7),
.B(n_8),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_5),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_6),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_136),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_20),
.Y(n_191)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_167),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_36),
.B(n_49),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_176),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_178),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_161),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_150),
.B1(n_146),
.B2(n_145),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_168),
.B1(n_175),
.B2(n_169),
.Y(n_197)
);

OA21x2_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_37),
.B(n_48),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_187),
.Y(n_198)
);

OAI322xp33_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_33),
.A3(n_46),
.B1(n_45),
.B2(n_42),
.C1(n_41),
.C2(n_18),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_173),
.C(n_179),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_200),
.C(n_183),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_178),
.B(n_172),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_185),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_186),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_204),
.C(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

AOI321xp33_ASAP7_75t_L g211 ( 
.A1(n_208),
.A2(n_209),
.A3(n_205),
.B1(n_202),
.B2(n_206),
.C(n_38),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_193),
.B1(n_191),
.B2(n_198),
.Y(n_209)
);

AOI21x1_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_53),
.B(n_40),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_210),
.C(n_30),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_64),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_13),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_14),
.Y(n_216)
);


endmodule