module fake_jpeg_9918_n_38 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_3),
.B(n_9),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_6),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx9p33_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.C(n_28),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_16),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_13),
.B1(n_23),
.B2(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_17),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_30),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_29),
.Y(n_36)
);

AOI31xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_15),
.A3(n_21),
.B(n_13),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_21),
.B(n_17),
.Y(n_38)
);


endmodule