module real_aes_4171_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_393;
wire n_84;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g295 ( .A(n_0), .B(n_233), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_1), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g366 ( .A1(n_2), .A2(n_238), .B(n_367), .C(n_368), .Y(n_366) );
OAI22xp33_ASAP7_75t_L g300 ( .A1(n_3), .A2(n_66), .B1(n_244), .B2(n_301), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_4), .A2(n_31), .B1(n_119), .B2(n_126), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_5), .A2(n_48), .B1(n_139), .B2(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g159 ( .A(n_6), .Y(n_159) );
AOI211x1_ASAP7_75t_L g143 ( .A1(n_7), .A2(n_144), .B(n_149), .C(n_180), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_8), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_9), .A2(n_37), .B1(n_161), .B2(n_170), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_10), .A2(n_56), .B1(n_264), .B2(n_301), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_11), .Y(n_330) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVxp67_ASAP7_75t_L g169 ( .A(n_12), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_12), .B(n_58), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_13), .A2(n_51), .B1(n_244), .B2(n_249), .Y(n_344) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_14), .A2(n_55), .B(n_236), .Y(n_235) );
OA21x2_ASAP7_75t_L g279 ( .A1(n_14), .A2(n_55), .B(n_236), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g100 ( .A(n_15), .B(n_90), .Y(n_100) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_16), .A2(n_18), .B1(n_131), .B2(n_135), .Y(n_130) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_17), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_19), .Y(n_283) );
BUFx3_ASAP7_75t_L g210 ( .A(n_20), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_21), .A2(n_246), .B(n_373), .C(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g189 ( .A(n_22), .Y(n_189) );
OAI22xp33_ASAP7_75t_SL g298 ( .A1(n_23), .A2(n_39), .B1(n_241), .B2(n_244), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_24), .A2(n_30), .B1(n_241), .B2(n_260), .Y(n_259) );
OAI22xp33_ASAP7_75t_SL g588 ( .A1(n_25), .A2(n_81), .B1(n_191), .B2(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_25), .Y(n_589) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_26), .Y(n_90) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_27), .Y(n_196) );
O2A1O1Ixp5_ASAP7_75t_L g309 ( .A1(n_28), .A2(n_238), .B(n_310), .C(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g91 ( .A(n_29), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_29), .B(n_57), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_32), .B(n_271), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_33), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_34), .A2(n_38), .B1(n_85), .B2(n_108), .Y(n_84) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_35), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_36), .Y(n_370) );
INVx1_ASAP7_75t_L g236 ( .A(n_40), .Y(n_236) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_41), .Y(n_221) );
AND2x4_ASAP7_75t_L g251 ( .A(n_41), .B(n_219), .Y(n_251) );
AND2x4_ASAP7_75t_L g277 ( .A(n_41), .B(n_219), .Y(n_277) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_42), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_43), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_44), .A2(n_238), .B(n_287), .C(n_289), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_45), .Y(n_318) );
INVx2_ASAP7_75t_L g335 ( .A(n_46), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_47), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_49), .B(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_50), .Y(n_80) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_50), .A2(n_64), .B1(n_263), .B2(n_265), .Y(n_262) );
OA22x2_ASAP7_75t_L g95 ( .A1(n_52), .A2(n_58), .B1(n_90), .B2(n_94), .Y(n_95) );
INVx1_ASAP7_75t_L g115 ( .A(n_52), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_53), .Y(n_250) );
NAND2xp33_ASAP7_75t_R g348 ( .A(n_54), .B(n_279), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_54), .A2(n_76), .B1(n_271), .B2(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g107 ( .A(n_57), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_57), .B(n_113), .Y(n_179) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_57), .Y(n_213) );
OAI21xp33_ASAP7_75t_L g116 ( .A1(n_58), .A2(n_65), .B(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_59), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_60), .Y(n_334) );
INVx1_ASAP7_75t_L g150 ( .A(n_61), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_62), .Y(n_331) );
INVx1_ASAP7_75t_L g185 ( .A(n_63), .Y(n_185) );
INVx1_ASAP7_75t_L g93 ( .A(n_65), .Y(n_93) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_65), .B(n_73), .Y(n_177) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_67), .Y(n_242) );
BUFx5_ASAP7_75t_L g244 ( .A(n_67), .Y(n_244) );
INVx1_ASAP7_75t_L g261 ( .A(n_67), .Y(n_261) );
INVx2_ASAP7_75t_L g378 ( .A(n_68), .Y(n_378) );
INVx2_ASAP7_75t_L g292 ( .A(n_69), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_70), .Y(n_375) );
INVx2_ASAP7_75t_SL g219 ( .A(n_71), .Y(n_219) );
INVx1_ASAP7_75t_L g316 ( .A(n_72), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g98 ( .A(n_73), .B(n_99), .Y(n_98) );
INVx2_ASAP7_75t_L g322 ( .A(n_74), .Y(n_322) );
OAI21xp33_ASAP7_75t_SL g281 ( .A1(n_75), .A2(n_244), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_76), .B(n_271), .Y(n_325) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_76), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_205), .B1(n_222), .B2(n_574), .C(n_581), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_192), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_190), .B2(n_191), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_80), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_81), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_81), .A2(n_191), .B1(n_583), .B2(n_584), .Y(n_582) );
INVxp33_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_143), .Y(n_82) );
AND4x1_ASAP7_75t_L g83 ( .A(n_84), .B(n_118), .C(n_130), .D(n_138), .Y(n_83) );
BUFx8_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_96), .Y(n_86) );
AND2x4_ASAP7_75t_L g132 ( .A(n_87), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g154 ( .A(n_87), .B(n_128), .Y(n_154) );
AND2x2_ASAP7_75t_L g188 ( .A(n_87), .B(n_124), .Y(n_188) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
INVx1_ASAP7_75t_L g122 ( .A(n_88), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
NAND2xp33_ASAP7_75t_L g89 ( .A(n_90), .B(n_91), .Y(n_89) );
INVx2_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx3_ASAP7_75t_L g99 ( .A(n_90), .Y(n_99) );
NAND2xp33_ASAP7_75t_L g106 ( .A(n_90), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g117 ( .A(n_90), .Y(n_117) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_91), .B(n_115), .Y(n_114) );
INVxp67_ASAP7_75t_L g214 ( .A(n_91), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g92 ( .A(n_93), .B(n_94), .Y(n_92) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_93), .A2(n_117), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g123 ( .A(n_95), .Y(n_123) );
AND2x2_ASAP7_75t_L g148 ( .A(n_95), .B(n_122), .Y(n_148) );
AND2x2_ASAP7_75t_L g167 ( .A(n_95), .B(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g110 ( .A(n_96), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g140 ( .A(n_96), .B(n_121), .Y(n_140) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_101), .Y(n_96) );
AND2x4_ASAP7_75t_L g124 ( .A(n_97), .B(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g129 ( .A(n_97), .Y(n_129) );
OR2x2_ASAP7_75t_L g134 ( .A(n_97), .B(n_102), .Y(n_134) );
AND2x2_ASAP7_75t_L g163 ( .A(n_97), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_99), .B(n_105), .Y(n_104) );
INVxp67_ASAP7_75t_L g113 ( .A(n_99), .Y(n_113) );
NAND3xp33_ASAP7_75t_L g178 ( .A(n_100), .B(n_112), .C(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g125 ( .A(n_103), .Y(n_125) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx8_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g136 ( .A(n_111), .B(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g184 ( .A(n_111), .B(n_128), .Y(n_184) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_116), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_115), .Y(n_215) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
AND2x2_ASAP7_75t_L g127 ( .A(n_121), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g142 ( .A(n_121), .B(n_137), .Y(n_142) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x4_ASAP7_75t_L g147 ( .A(n_124), .B(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g128 ( .A(n_125), .B(n_129), .Y(n_128) );
BUFx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g158 ( .A(n_128), .B(n_148), .Y(n_158) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g137 ( .A(n_134), .Y(n_137) );
BUFx12f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_155), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI21xp5_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_159), .B(n_160), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx4f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_167), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g174 ( .A(n_165), .Y(n_174) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_166), .Y(n_211) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_178), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_185), .B1(n_186), .B2(n_189), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B1(n_203), .B2(n_204), .Y(n_192) );
INVx1_ASAP7_75t_L g203 ( .A(n_193), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_194), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_198) );
INVx1_ASAP7_75t_L g202 ( .A(n_199), .Y(n_202) );
INVx1_ASAP7_75t_L g201 ( .A(n_200), .Y(n_201) );
BUFx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_216), .Y(n_207) );
INVxp67_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g586 ( .A(n_209), .B(n_216), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .C(n_215), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_220), .Y(n_216) );
OR2x2_ASAP7_75t_L g591 ( .A(n_217), .B(n_221), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_217), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_217), .B(n_220), .Y(n_595) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVxp33_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND3x4_ASAP7_75t_L g223 ( .A(n_224), .B(n_477), .C(n_528), .Y(n_223) );
NOR2x1_ASAP7_75t_L g224 ( .A(n_225), .B(n_422), .Y(n_224) );
NAND3xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_395), .C(n_407), .Y(n_225) );
AOI221xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_303), .B1(n_337), .B2(n_362), .C(n_379), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_272), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_228), .B(n_355), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_228), .B(n_436), .Y(n_472) );
AND2x2_ASAP7_75t_L g531 ( .A(n_228), .B(n_411), .Y(n_531) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g396 ( .A(n_229), .Y(n_396) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_255), .Y(n_229) );
AND2x2_ASAP7_75t_L g356 ( .A(n_230), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g426 ( .A(n_230), .B(n_412), .Y(n_426) );
AND2x2_ASAP7_75t_L g461 ( .A(n_230), .B(n_294), .Y(n_461) );
AND2x2_ASAP7_75t_L g489 ( .A(n_230), .B(n_490), .Y(n_489) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_237), .B(n_252), .Y(n_230) );
OA21x2_ASAP7_75t_L g353 ( .A1(n_231), .A2(n_237), .B(n_252), .Y(n_353) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g447 ( .A(n_232), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_SL g376 ( .A(n_233), .B(n_319), .Y(n_376) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g271 ( .A(n_234), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_234), .B(n_251), .Y(n_302) );
NOR2xp33_ASAP7_75t_SL g377 ( .A(n_234), .B(n_378), .Y(n_377) );
INVx4_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g254 ( .A(n_235), .Y(n_254) );
BUFx3_ASAP7_75t_L g268 ( .A(n_235), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .B1(n_246), .B2(n_247), .C(n_251), .Y(n_237) );
INVx1_ASAP7_75t_L g336 ( .A(n_238), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_238), .A2(n_285), .B1(n_344), .B2(n_345), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_238), .A2(n_285), .B1(n_329), .B2(n_333), .Y(n_446) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g246 ( .A(n_239), .Y(n_246) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_239), .Y(n_258) );
INVx1_ASAP7_75t_L g266 ( .A(n_239), .Y(n_266) );
INVx4_ASAP7_75t_L g285 ( .A(n_239), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_239), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_239), .B(n_316), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_241), .A2(n_243), .B1(n_244), .B2(n_245), .Y(n_240) );
INVx2_ASAP7_75t_SL g265 ( .A(n_241), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_241), .A2(n_244), .B1(n_330), .B2(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g369 ( .A(n_241), .Y(n_369) );
INVx6_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g249 ( .A(n_242), .Y(n_249) );
INVx3_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
INVx2_ASAP7_75t_L g301 ( .A(n_242), .Y(n_301) );
INVx1_ASAP7_75t_L g597 ( .A(n_243), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_244), .A2(n_248), .B1(n_249), .B2(n_250), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_244), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_244), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_244), .B(n_318), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_246), .A2(n_300), .B(n_302), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_249), .A2(n_260), .B1(n_334), .B2(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g373 ( .A(n_249), .Y(n_373) );
INVx1_ASAP7_75t_L g583 ( .A(n_250), .Y(n_583) );
INVx1_ASAP7_75t_L g347 ( .A(n_251), .Y(n_347) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_251), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g346 ( .A(n_253), .B(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_254), .B(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g320 ( .A(n_254), .Y(n_320) );
AND2x4_ASAP7_75t_L g456 ( .A(n_255), .B(n_352), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_267), .B(n_269), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_257), .A2(n_270), .B(n_359), .Y(n_358) );
OA22x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B1(n_262), .B2(n_266), .Y(n_257) );
INVx4_ASAP7_75t_L g580 ( .A(n_258), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_260), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_260), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g264 ( .A(n_261), .Y(n_264) );
INVx1_ASAP7_75t_L g367 ( .A(n_263), .Y(n_367) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_293), .Y(n_273) );
BUFx2_ASAP7_75t_L g350 ( .A(n_274), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_274), .B(n_294), .Y(n_355) );
INVx2_ASAP7_75t_L g383 ( .A(n_274), .Y(n_383) );
AND2x2_ASAP7_75t_L g400 ( .A(n_274), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g416 ( .A(n_274), .B(n_412), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_274), .B(n_353), .Y(n_476) );
INVx1_ASAP7_75t_L g482 ( .A(n_274), .Y(n_482) );
INVx2_ASAP7_75t_L g501 ( .A(n_274), .Y(n_501) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI21x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B(n_291), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx4_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_277), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g323 ( .A(n_279), .Y(n_323) );
BUFx3_ASAP7_75t_L g361 ( .A(n_279), .Y(n_361) );
INVx2_ASAP7_75t_L g394 ( .A(n_279), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B(n_286), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_284), .A2(n_319), .B1(n_328), .B2(n_332), .C(n_336), .Y(n_327) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_285), .A2(n_314), .B1(n_315), .B2(n_317), .Y(n_313) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g310 ( .A(n_288), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
AND2x4_ASAP7_75t_L g351 ( .A(n_293), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g552 ( .A(n_293), .B(n_357), .Y(n_552) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g399 ( .A(n_294), .Y(n_399) );
INVx3_ASAP7_75t_L g412 ( .A(n_294), .Y(n_412) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_324), .Y(n_305) );
AND2x4_ASAP7_75t_L g339 ( .A(n_306), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g568 ( .A(n_306), .B(n_501), .Y(n_568) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g389 ( .A(n_307), .Y(n_389) );
AND2x2_ASAP7_75t_L g403 ( .A(n_307), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_307), .B(n_364), .Y(n_441) );
BUFx2_ASAP7_75t_R g451 ( .A(n_307), .Y(n_451) );
AND2x2_ASAP7_75t_L g527 ( .A(n_307), .B(n_507), .Y(n_527) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_307), .Y(n_535) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_320), .B(n_321), .Y(n_307) );
NOR3xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_313), .C(n_319), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_320), .B(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g363 ( .A(n_324), .B(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g406 ( .A(n_324), .B(n_364), .Y(n_406) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_324), .Y(n_414) );
AND2x2_ASAP7_75t_L g537 ( .A(n_324), .B(n_433), .Y(n_537) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g390 ( .A(n_326), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_349), .B(n_354), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g480 ( .A(n_339), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g516 ( .A(n_339), .B(n_386), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_339), .B(n_483), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g538 ( .A(n_339), .B(n_425), .C(n_481), .D(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g547 ( .A(n_339), .B(n_470), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_339), .B(n_452), .Y(n_560) );
INVx1_ASAP7_75t_L g421 ( .A(n_340), .Y(n_421) );
AND2x2_ASAP7_75t_L g545 ( .A(n_340), .B(n_507), .Y(n_545) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g404 ( .A(n_341), .Y(n_404) );
AND2x2_ASAP7_75t_L g442 ( .A(n_341), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g495 ( .A(n_341), .B(n_389), .Y(n_495) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_341), .Y(n_513) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_348), .Y(n_341) );
AND2x2_ASAP7_75t_L g391 ( .A(n_342), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_349), .A2(n_530), .B1(n_532), .B2(n_536), .C(n_538), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_351), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_351), .B(n_382), .Y(n_459) );
AND2x4_ASAP7_75t_L g485 ( .A(n_351), .B(n_474), .Y(n_485) );
AND2x2_ASAP7_75t_L g496 ( .A(n_351), .B(n_425), .Y(n_496) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g401 ( .A(n_353), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g380 ( .A(n_356), .Y(n_380) );
AOI322xp5_ASAP7_75t_L g479 ( .A1(n_356), .A2(n_388), .A3(n_469), .B1(n_480), .B2(n_483), .C1(n_485), .C2(n_486), .Y(n_479) );
INVx3_ASAP7_75t_L g410 ( .A(n_357), .Y(n_410) );
INVx1_ASAP7_75t_L g490 ( .A(n_357), .Y(n_490) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g384 ( .A(n_358), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_360), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI32xp33_ASAP7_75t_L g550 ( .A1(n_362), .A2(n_551), .A3(n_553), .B1(n_554), .B2(n_555), .Y(n_550) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_363), .B(n_451), .Y(n_493) );
AND2x2_ASAP7_75t_L g497 ( .A(n_363), .B(n_403), .Y(n_497) );
INVx1_ASAP7_75t_L g387 ( .A(n_364), .Y(n_387) );
INVx1_ASAP7_75t_L g433 ( .A(n_364), .Y(n_433) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_364), .Y(n_453) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_364), .Y(n_463) );
AND2x4_ASAP7_75t_L g470 ( .A(n_364), .B(n_443), .Y(n_470) );
INVx2_ASAP7_75t_L g507 ( .A(n_364), .Y(n_507) );
AO31x2_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_371), .A3(n_376), .B(n_377), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_373), .Y(n_577) );
AOI21xp33_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_381), .B(n_385), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g509 ( .A(n_381), .B(n_426), .Y(n_509) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g508 ( .A(n_382), .B(n_426), .Y(n_508) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g437 ( .A(n_383), .Y(n_437) );
INVx1_ASAP7_75t_L g455 ( .A(n_383), .Y(n_455) );
AND2x2_ASAP7_75t_L g551 ( .A(n_383), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_384), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g474 ( .A(n_384), .Y(n_474) );
OR2x2_ASAP7_75t_L g499 ( .A(n_384), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g564 ( .A(n_385), .Y(n_564) );
NAND2x1p5_ASAP7_75t_SL g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g540 ( .A(n_387), .Y(n_540) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g420 ( .A(n_389), .Y(n_420) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_389), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_402), .Y(n_395) );
AOI321xp33_ASAP7_75t_L g565 ( .A1(n_396), .A2(n_467), .A3(n_566), .B1(n_567), .B2(n_569), .C(n_570), .Y(n_565) );
AND2x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NOR2xp67_ASAP7_75t_L g475 ( .A(n_399), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_401), .B(n_482), .Y(n_556) );
INVx2_ASAP7_75t_L g572 ( .A(n_401), .Y(n_572) );
AOI22x1_ASAP7_75t_L g407 ( .A1(n_402), .A2(n_408), .B1(n_413), .B2(n_417), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_402), .A2(n_424), .B(n_427), .Y(n_423) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
AND2x4_ASAP7_75t_L g469 ( .A(n_403), .B(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_403), .A2(n_406), .B1(n_483), .B2(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_403), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g553 ( .A(n_403), .Y(n_553) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g522 ( .A(n_406), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g570 ( .A(n_409), .B(n_568), .C(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx3_ASAP7_75t_L g425 ( .A(n_410), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_410), .B(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g467 ( .A(n_410), .B(n_426), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_410), .B(n_416), .Y(n_468) );
BUFx3_ASAP7_75t_L g549 ( .A(n_411), .Y(n_549) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_412), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_SL g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NAND2xp33_ASAP7_75t_L g498 ( .A(n_415), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g458 ( .A(n_419), .B(n_453), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_438), .C(n_464), .Y(n_422) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AND2x2_ASAP7_75t_L g515 ( .A(n_425), .B(n_461), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_425), .B(n_426), .Y(n_524) );
OAI22xp33_ASAP7_75t_SL g427 ( .A1(n_428), .A2(n_431), .B1(n_432), .B2(n_435), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx2_ASAP7_75t_L g566 ( .A(n_432), .Y(n_566) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AND2x2_ASAP7_75t_L g554 ( .A(n_433), .B(n_442), .Y(n_554) );
OR2x2_ASAP7_75t_L g462 ( .A(n_434), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
O2A1O1Ixp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_449), .B(n_454), .C(n_457), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_439), .A2(n_485), .B1(n_489), .B2(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g439 ( .A(n_440), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_442), .A2(n_465), .B1(n_469), .B2(n_471), .Y(n_464) );
AND2x2_ASAP7_75t_L g526 ( .A(n_442), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g484 ( .A(n_443), .Y(n_484) );
OAI21x1_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B(n_447), .Y(n_443) );
AND2x2_ASAP7_75t_SL g575 ( .A(n_445), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g543 ( .A(n_455), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B1(n_460), .B2(n_462), .Y(n_457) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_462), .B(n_568), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_467), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_467), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_470), .B(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g533 ( .A(n_470), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
BUFx2_ASAP7_75t_SL g562 ( .A(n_475), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_502), .C(n_521), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
INVx1_ASAP7_75t_L g487 ( .A(n_481), .Y(n_487) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g519 ( .A(n_489), .B(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_491) );
NAND2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AND2x2_ASAP7_75t_L g504 ( .A(n_495), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g523 ( .A(n_495), .Y(n_523) );
INVx1_ASAP7_75t_L g563 ( .A(n_500), .Y(n_563) );
BUFx2_ASAP7_75t_L g520 ( .A(n_501), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_507), .Y(n_573) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_517), .B2(n_519), .Y(n_514) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_524), .B(n_525), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_541), .C(n_557), .Y(n_528) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_544), .B1(n_546), .B2(n_548), .C(n_550), .Y(n_541) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .C(n_565), .Y(n_557) );
INVxp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_564), .Y(n_561) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_576), .A2(n_594), .B(n_595), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI222xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B1(n_587), .B2(n_590), .C1(n_592), .C2(n_596), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_583), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
endmodule