module fake_jpeg_19111_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_8),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_16),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_27),
.C(n_19),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_21),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_30),
.B1(n_6),
.B2(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_8),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_2),
.B(n_3),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_7),
.Y(n_38)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_18),
.CI(n_37),
.CON(n_39),
.SN(n_39)
);


endmodule