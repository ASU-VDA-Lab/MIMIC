module real_jpeg_16058_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_213;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_0),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g16 ( 
.A1(n_1),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_17),
.B1(n_95),
.B2(n_97),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_17),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_2),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_6),
.Y(n_134)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_55),
.A3(n_56),
.B1(n_62),
.B2(n_65),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_7),
.A2(n_45),
.B1(n_73),
.B2(n_76),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_7),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_7),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_7),
.B(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_157),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_155),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_150),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_13),
.B(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_91),
.B1(n_92),
.B2(n_149),
.Y(n_13)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_14),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_53),
.B1(n_89),
.B2(n_90),
.Y(n_14)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_15),
.B(n_168),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_26),
.B1(n_36),
.B2(n_44),
.Y(n_15)
);

AO22x2_ASAP7_75t_L g154 ( 
.A1(n_16),
.A2(n_26),
.B1(n_36),
.B2(n_44),
.Y(n_154)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_36),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_36),
.Y(n_207)
);

AO22x2_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_36)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_39),
.Y(n_145)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_42),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B(n_50),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_50),
.A2(n_83),
.A3(n_174),
.B1(n_178),
.B2(n_182),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_70),
.Y(n_53)
);

XOR2x2_ASAP7_75t_SL g153 ( 
.A(n_54),
.B(n_70),
.Y(n_153)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_79),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_71),
.A2(n_139),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_72),
.B(n_80),
.Y(n_146)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_75),
.Y(n_200)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_85),
.Y(n_202)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_163),
.C(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_124),
.B1(n_125),
.B2(n_148),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_93),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_99),
.B1(n_106),
.B2(n_115),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_94),
.A2(n_99),
.B1(n_106),
.B2(n_115),
.Y(n_152)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2x1p5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

OA22x2_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_129)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_135),
.B2(n_147),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_195),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_139),
.B(n_146),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_147),
.B(n_210),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_147),
.B(n_210),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_154),
.A2(n_161),
.B1(n_173),
.B2(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_170),
.B(n_214),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_162),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_192),
.B(n_213),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_188),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_188),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_209),
.B(n_212),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_203),
.B(n_208),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);


endmodule