module fake_netlist_1_8210_n_718 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_718, n_391);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_718;
output n_391;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_703;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_195;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_77), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_18), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_76), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_52), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_31), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g86 ( .A(n_73), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_20), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_44), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_51), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_36), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_53), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_37), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_70), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_58), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_60), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_16), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_9), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_34), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_17), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_26), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_28), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_46), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_30), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_41), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_32), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_17), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_5), .Y(n_111) );
BUFx5_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_39), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_23), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_42), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_3), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_72), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_67), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_54), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_55), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_19), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_5), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_10), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_22), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_119), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_112), .B(n_0), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_96), .B(n_0), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_121), .B(n_1), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_87), .B(n_1), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_82), .B(n_2), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_81), .B(n_2), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_108), .B(n_4), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_87), .B(n_88), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_83), .B(n_4), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_86), .B(n_6), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_101), .B(n_109), .Y(n_148) );
INVxp67_ASAP7_75t_L g149 ( .A(n_111), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_102), .B(n_6), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_126), .B(n_7), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_112), .B(n_7), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_119), .B(n_40), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_97), .B(n_8), .Y(n_155) );
BUFx2_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_112), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_89), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_97), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_122), .B(n_8), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_89), .Y(n_162) );
BUFx8_ASAP7_75t_L g163 ( .A(n_112), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_126), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_93), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_104), .B(n_9), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_93), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_127), .B(n_10), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_112), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_127), .B(n_11), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_94), .Y(n_171) );
NAND2xp33_ASAP7_75t_R g172 ( .A(n_95), .B(n_45), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_110), .B(n_11), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_88), .B(n_12), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_132), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_136), .A2(n_113), .B1(n_128), .B2(n_98), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
NOR3xp33_ASAP7_75t_L g179 ( .A(n_134), .B(n_113), .C(n_128), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_159), .Y(n_180) );
NAND3xp33_ASAP7_75t_L g181 ( .A(n_163), .B(n_98), .C(n_107), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_143), .B(n_105), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_156), .B(n_90), .Y(n_183) );
INVx1_ASAP7_75t_SL g184 ( .A(n_147), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_143), .B(n_105), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_143), .B(n_94), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_149), .B(n_106), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_143), .B(n_125), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_135), .B(n_92), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_151), .B(n_125), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_135), .B(n_92), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_151), .B(n_124), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_168), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_130), .B(n_107), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_168), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_130), .B(n_124), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_139), .B(n_116), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_144), .B(n_12), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
OR2x2_ASAP7_75t_SL g215 ( .A(n_144), .B(n_120), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_161), .Y(n_216) );
BUFx10_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_157), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_153), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_158), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_148), .B(n_13), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_161), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_154), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_158), .B(n_95), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_163), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_162), .Y(n_229) );
AO22x2_ASAP7_75t_L g230 ( .A1(n_162), .A2(n_117), .B1(n_114), .B2(n_115), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_165), .B(n_123), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_165), .A2(n_106), .B1(n_118), .B2(n_129), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_167), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_167), .B(n_112), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_171), .B(n_146), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_171), .B(n_91), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_146), .B(n_100), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_131), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_157), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_157), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_217), .Y(n_241) );
NOR2x1_ASAP7_75t_L g242 ( .A(n_181), .B(n_173), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_179), .A2(n_172), .B1(n_163), .B2(n_145), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_217), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_217), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_196), .B(n_174), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_187), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_228), .B(n_163), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_187), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_227), .B(n_166), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_187), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_240), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_231), .B(n_150), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_228), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_193), .A2(n_142), .B1(n_138), .B2(n_174), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_176), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_231), .B(n_236), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_213), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_193), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_240), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_193), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_184), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_234), .Y(n_264) );
INVxp67_ASAP7_75t_SL g265 ( .A(n_213), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_178), .Y(n_266) );
AND2x6_ASAP7_75t_SL g267 ( .A(n_237), .B(n_138), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_231), .B(n_140), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_240), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_193), .Y(n_271) );
NOR2x2_ASAP7_75t_L g272 ( .A(n_232), .B(n_169), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_214), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_193), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_193), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_183), .B(n_160), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_237), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_188), .B(n_155), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_198), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_236), .B(n_146), .Y(n_280) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_237), .B(n_164), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_218), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_236), .B(n_196), .Y(n_283) );
INVx5_ASAP7_75t_L g284 ( .A(n_226), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_200), .B(n_133), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_202), .B(n_164), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_198), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_198), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_198), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_204), .B(n_164), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_238), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_177), .B(n_164), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_203), .A2(n_152), .B1(n_154), .B2(n_146), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_221), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_198), .A2(n_154), .B1(n_169), .B2(n_131), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_222), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_200), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_206), .B(n_154), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_223), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_224), .B(n_169), .Y(n_301) );
BUFx4f_ASAP7_75t_SL g302 ( .A(n_224), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_198), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
AOI22xp33_ASAP7_75t_SL g306 ( .A1(n_230), .A2(n_154), .B1(n_112), .B2(n_131), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_180), .Y(n_307) );
AND2x4_ASAP7_75t_SL g308 ( .A(n_211), .B(n_131), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_180), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_182), .B(n_131), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_265), .B(n_207), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_260), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_259), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_259), .Y(n_314) );
BUFx12f_ASAP7_75t_L g315 ( .A(n_256), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_260), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_246), .B(n_211), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_246), .A2(n_230), .B1(n_209), .B2(n_201), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_283), .A2(n_230), .B1(n_201), .B2(n_186), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_256), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_260), .B(n_211), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_273), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_301), .B(n_208), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_247), .A2(n_186), .B1(n_201), .B2(n_182), .Y(n_324) );
NOR2x1_ASAP7_75t_L g325 ( .A(n_266), .B(n_182), .Y(n_325) );
BUFx4f_ASAP7_75t_L g326 ( .A(n_247), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_274), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_252), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_254), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_186), .B1(n_199), .B2(n_197), .C1(n_208), .C2(n_235), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_263), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_274), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_266), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_301), .B(n_208), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_302), .B(n_215), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_270), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_249), .B(n_226), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_282), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_270), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_254), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_277), .A2(n_230), .B1(n_215), .B2(n_154), .Y(n_342) );
AOI21x1_ASAP7_75t_L g343 ( .A1(n_298), .A2(n_239), .B(n_175), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_249), .B(n_226), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_277), .Y(n_345) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_267), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_252), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_254), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_281), .Y(n_349) );
O2A1O1Ixp5_ASAP7_75t_L g350 ( .A1(n_248), .A2(n_239), .B(n_175), .C(n_189), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_261), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_251), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_250), .B(n_219), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_275), .Y(n_354) );
INVx5_ASAP7_75t_L g355 ( .A(n_254), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_282), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_281), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_251), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_304), .A2(n_154), .B1(n_226), .B2(n_191), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_257), .B(n_219), .Y(n_360) );
BUFx2_ASAP7_75t_SL g361 ( .A(n_275), .Y(n_361) );
OAI33xp33_ASAP7_75t_L g362 ( .A1(n_253), .A2(n_191), .A3(n_189), .B1(n_185), .B2(n_190), .B3(n_205), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_276), .A2(n_226), .B1(n_154), .B2(n_131), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_241), .Y(n_364) );
BUFx6f_ASAP7_75t_SL g365 ( .A(n_279), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_315), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_337), .A2(n_241), .B1(n_244), .B2(n_245), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_316), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_320), .B(n_268), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_315), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_326), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_320), .A2(n_272), .B1(n_304), .B2(n_279), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_316), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_328), .Y(n_375) );
BUFx10_ASAP7_75t_L g376 ( .A(n_321), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_326), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_334), .A2(n_292), .B1(n_278), .B2(n_258), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_352), .B(n_258), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_318), .A2(n_255), .B1(n_243), .B2(n_296), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_337), .B(n_286), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_316), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_352), .B(n_264), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_334), .B(n_264), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_328), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_357), .A2(n_340), .B1(n_345), .B2(n_346), .Y(n_386) );
O2A1O1Ixp5_ASAP7_75t_SL g387 ( .A1(n_322), .A2(n_285), .B(n_296), .C(n_294), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_353), .A2(n_294), .B(n_300), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_326), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_357), .A2(n_288), .B1(n_300), .B2(n_299), .Y(n_390) );
UNKNOWN g391 ( );
AND2x2_ASAP7_75t_L g392 ( .A(n_358), .B(n_299), .Y(n_392) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_338), .B(n_244), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_345), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_336), .A2(n_280), .B1(n_290), .B2(n_306), .C(n_303), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_324), .A2(n_288), .B1(n_303), .B2(n_245), .Y(n_396) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_311), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_332), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_373), .A2(n_342), .B1(n_340), .B2(n_313), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_391), .A2(n_314), .B1(n_325), .B2(n_319), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_388), .A2(n_362), .B(n_339), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_392), .B(n_358), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_383), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g405 ( .A1(n_394), .A2(n_349), .B1(n_364), .B2(n_317), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_376), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_375), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_385), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_392), .B(n_330), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_380), .A2(n_356), .B1(n_286), .B2(n_242), .Y(n_411) );
BUFx12f_ASAP7_75t_L g412 ( .A(n_366), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_381), .A2(n_286), .B1(n_242), .B2(n_335), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_394), .A2(n_364), .B1(n_323), .B2(n_321), .Y(n_415) );
BUFx5_ASAP7_75t_L g416 ( .A(n_389), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_379), .B(n_321), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_383), .A2(n_298), .B1(n_360), .B2(n_365), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_369), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_390), .A2(n_359), .B1(n_355), .B2(n_361), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_368), .Y(n_421) );
NOR2xp33_ASAP7_75t_SL g422 ( .A(n_389), .B(n_355), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_384), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
INVx4_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_379), .B(n_347), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_378), .A2(n_293), .B1(n_310), .B2(n_350), .C(n_363), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_383), .B(n_347), .Y(n_428) );
OA21x2_ASAP7_75t_L g429 ( .A1(n_402), .A2(n_395), .B(n_387), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_415), .B(n_387), .C(n_367), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_415), .A2(n_386), .B1(n_396), .B2(n_384), .Y(n_431) );
OAI211xp5_ASAP7_75t_SL g432 ( .A1(n_405), .A2(n_399), .B(n_370), .C(n_372), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_400), .A2(n_370), .B1(n_371), .B2(n_376), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g434 ( .A1(n_405), .A2(n_377), .B(n_382), .Y(n_434) );
OA21x2_ASAP7_75t_L g435 ( .A1(n_402), .A2(n_295), .B(n_343), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_406), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_412), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_426), .B(n_351), .Y(n_440) );
INVx5_ASAP7_75t_L g441 ( .A(n_425), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_421), .A2(n_366), .B1(n_397), .B2(n_371), .C(n_308), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_421), .A2(n_308), .B1(n_298), .B2(n_374), .C(n_369), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_408), .Y(n_444) );
OAI31xp33_ASAP7_75t_L g445 ( .A1(n_420), .A2(n_310), .A3(n_374), .B(n_369), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_413), .A2(n_393), .B(n_382), .C(n_374), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_408), .Y(n_447) );
AOI31xp33_ASAP7_75t_L g448 ( .A1(n_420), .A2(n_310), .A3(n_351), .B(n_344), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_404), .A2(n_382), .B1(n_365), .B2(n_333), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_426), .B(n_338), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_409), .A2(n_414), .B(n_411), .Y(n_452) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_427), .A2(n_194), .B(n_190), .Y(n_453) );
AOI31xp33_ASAP7_75t_L g454 ( .A1(n_423), .A2(n_344), .A3(n_338), .B(n_365), .Y(n_454) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_427), .A2(n_192), .B(n_194), .Y(n_455) );
OAI211xp5_ASAP7_75t_L g456 ( .A1(n_423), .A2(n_355), .B(n_269), .C(n_261), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g457 ( .A1(n_424), .A2(n_341), .B(n_329), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_409), .Y(n_458) );
BUFx3_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_424), .A2(n_269), .B1(n_344), .B2(n_287), .C(n_262), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_426), .B(n_355), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_403), .A2(n_333), .B1(n_341), .B2(n_354), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_428), .B(n_355), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_414), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_447), .B(n_414), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_431), .A2(n_403), .B1(n_410), .B2(n_401), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_436), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_439), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_447), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_436), .Y(n_470) );
OAI31xp33_ASAP7_75t_L g471 ( .A1(n_432), .A2(n_403), .A3(n_410), .B(n_407), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_432), .A2(n_417), .B1(n_428), .B2(n_425), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_441), .B(n_419), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_464), .B(n_428), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_440), .B(n_417), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_439), .Y(n_477) );
AOI211x1_ASAP7_75t_SL g478 ( .A1(n_430), .A2(n_419), .B(n_15), .C(n_18), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_439), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_440), .B(n_417), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_464), .B(n_419), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_449), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_444), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_449), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_438), .Y(n_487) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_442), .A2(n_418), .B(n_425), .C(n_407), .Y(n_488) );
OAI211xp5_ASAP7_75t_SL g489 ( .A1(n_442), .A2(n_192), .B(n_195), .C(n_205), .Y(n_489) );
OAI31xp33_ASAP7_75t_L g490 ( .A1(n_434), .A2(n_422), .A3(n_262), .B(n_271), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_449), .B(n_416), .Y(n_491) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_448), .B(n_425), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_430), .A2(n_422), .B(n_185), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_458), .B(n_416), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_441), .B(n_329), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_458), .B(n_416), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_441), .B(n_329), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_458), .B(n_416), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
AO221x2_ASAP7_75t_L g500 ( .A1(n_434), .A2(n_14), .B1(n_15), .B2(n_19), .C(n_20), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_429), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_461), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_433), .A2(n_412), .B1(n_416), .B2(n_354), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_441), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_441), .Y(n_505) );
OAI31xp33_ASAP7_75t_SL g506 ( .A1(n_446), .A2(n_416), .A3(n_412), .B(n_14), .Y(n_506) );
BUFx2_ASAP7_75t_SL g507 ( .A(n_441), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_429), .Y(n_508) );
OAI33xp33_ASAP7_75t_L g509 ( .A1(n_445), .A2(n_212), .A3(n_210), .B1(n_195), .B2(n_225), .B3(n_448), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_463), .B(n_416), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_463), .B(n_416), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_441), .B(n_416), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_445), .B(n_220), .C(n_216), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_459), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_468), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_491), .B(n_453), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_504), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_474), .B(n_459), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g519 ( .A(n_506), .B(n_443), .C(n_459), .D(n_462), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_474), .B(n_454), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
BUFx3_ASAP7_75t_L g522 ( .A(n_473), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_499), .B(n_452), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_510), .B(n_455), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_470), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_476), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_487), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_481), .Y(n_528) );
NOR2xp33_ASAP7_75t_SL g529 ( .A(n_507), .B(n_416), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_500), .A2(n_446), .B1(n_456), .B2(n_443), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_502), .B(n_452), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_465), .B(n_469), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_465), .B(n_454), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_496), .B(n_455), .Y(n_534) );
AND2x6_ASAP7_75t_L g535 ( .A(n_512), .B(n_456), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_466), .B(n_429), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_488), .B(n_457), .C(n_460), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_468), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_507), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_491), .B(n_453), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_494), .B(n_453), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_485), .B(n_429), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_509), .B(n_457), .C(n_460), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_483), .B(n_429), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_483), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_475), .B(n_450), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_477), .Y(n_547) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_505), .B(n_435), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_494), .B(n_435), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_492), .B(n_329), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_496), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_498), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_514), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_477), .Y(n_554) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_513), .B(n_435), .Y(n_555) );
NOR2x1_ASAP7_75t_L g556 ( .A(n_473), .B(n_435), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_511), .B(n_435), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_480), .B(n_348), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_500), .B(n_348), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_492), .B(n_348), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_479), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_500), .B(n_348), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_498), .B(n_225), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_479), .Y(n_564) );
AND4x1_ASAP7_75t_L g565 ( .A(n_471), .B(n_21), .C(n_24), .D(n_25), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_472), .B(n_348), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_501), .B(n_212), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_484), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_473), .B(n_27), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_472), .B(n_329), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_484), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_571), .Y(n_572) );
OAI33xp33_ASAP7_75t_L g573 ( .A1(n_536), .A2(n_521), .A3(n_526), .B1(n_525), .B2(n_528), .B3(n_546), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_532), .B(n_482), .Y(n_574) );
AOI322xp5_ASAP7_75t_L g575 ( .A1(n_527), .A2(n_508), .A3(n_501), .B1(n_503), .B2(n_478), .C1(n_486), .C2(n_497), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_545), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_571), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_552), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_553), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_551), .B(n_508), .Y(n_580) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_550), .A2(n_490), .B(n_493), .C(n_489), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_517), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_515), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_537), .B(n_482), .C(n_486), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_533), .B(n_497), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_554), .Y(n_586) );
NAND3xp33_ASAP7_75t_SL g587 ( .A(n_565), .B(n_497), .C(n_495), .Y(n_587) );
NAND2xp33_ASAP7_75t_SL g588 ( .A(n_550), .B(n_495), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_531), .B(n_495), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_522), .B(n_29), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_561), .Y(n_591) );
NOR2xp33_ASAP7_75t_R g592 ( .A(n_529), .B(n_35), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_523), .B(n_210), .Y(n_593) );
NAND2x2_ASAP7_75t_L g594 ( .A(n_520), .B(n_38), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_522), .B(n_43), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_518), .B(n_47), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_564), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_539), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_534), .B(n_220), .Y(n_599) );
AOI322xp5_ASAP7_75t_L g600 ( .A1(n_560), .A2(n_220), .A3(n_216), .B1(n_312), .B2(n_287), .C1(n_271), .C2(n_262), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_557), .B(n_216), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_530), .A2(n_216), .B(n_220), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_544), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_542), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_519), .B(n_48), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_568), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_515), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_538), .Y(n_608) );
INVxp33_ASAP7_75t_L g609 ( .A(n_560), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_569), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_559), .B(n_49), .Y(n_611) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_548), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_538), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_569), .B(n_254), .Y(n_614) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_569), .B(n_333), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_524), .B(n_50), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_563), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_549), .B(n_56), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_541), .B(n_57), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_537), .A2(n_312), .B(n_289), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_547), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_516), .B(n_59), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_605), .A2(n_540), .B1(n_535), .B2(n_543), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_603), .B(n_516), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_603), .B(n_540), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_604), .B(n_540), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g627 ( .A1(n_575), .A2(n_556), .B(n_562), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_579), .Y(n_628) );
NAND2xp33_ASAP7_75t_L g629 ( .A(n_592), .B(n_535), .Y(n_629) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_615), .B(n_535), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_604), .B(n_547), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_583), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_576), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_580), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_607), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_617), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_582), .B(n_535), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_574), .B(n_586), .Y(n_638) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_572), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_578), .B(n_555), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g641 ( .A(n_598), .B(n_563), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_572), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_577), .B(n_558), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_591), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_589), .B(n_567), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_597), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_606), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_608), .B(n_535), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_613), .B(n_543), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_621), .B(n_567), .Y(n_650) );
OAI21xp33_ASAP7_75t_L g651 ( .A1(n_605), .A2(n_570), .B(n_566), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_601), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_592), .Y(n_653) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_590), .B(n_312), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_612), .B(n_63), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_584), .B(n_64), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_609), .A2(n_65), .B(n_68), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_593), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_573), .A2(n_305), .B1(n_291), .B2(n_354), .C(n_327), .Y(n_659) );
XNOR2xp5_ASAP7_75t_L g660 ( .A(n_585), .B(n_74), .Y(n_660) );
NAND4xp25_ASAP7_75t_SL g661 ( .A(n_581), .B(n_75), .C(n_78), .D(n_79), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_612), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_588), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_599), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_610), .B(n_307), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_573), .A2(n_271), .B1(n_287), .B2(n_289), .C(n_307), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_594), .A2(n_289), .B1(n_284), .B2(n_309), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_SL g668 ( .A1(n_611), .A2(n_284), .B(n_618), .C(n_622), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_616), .B(n_284), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_619), .B(n_284), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_595), .Y(n_671) );
OAI21xp33_ASAP7_75t_SL g672 ( .A1(n_614), .A2(n_284), .B(n_611), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_614), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_596), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_602), .B(n_284), .Y(n_675) );
XOR2xp5_ASAP7_75t_L g676 ( .A(n_587), .B(n_594), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_587), .Y(n_677) );
NOR3xp33_ASAP7_75t_L g678 ( .A(n_620), .B(n_605), .C(n_432), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g679 ( .A(n_600), .B(n_487), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_617), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_603), .B(n_604), .Y(n_681) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_676), .A2(n_660), .A3(n_653), .B(n_677), .Y(n_682) );
NAND4xp25_ASAP7_75t_L g683 ( .A(n_623), .B(n_678), .C(n_627), .D(n_668), .Y(n_683) );
INVxp67_ASAP7_75t_L g684 ( .A(n_649), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_681), .A2(n_663), .B1(n_628), .B2(n_634), .C(n_662), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g686 ( .A(n_641), .B(n_636), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g687 ( .A1(n_679), .A2(n_668), .B(n_660), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_681), .Y(n_688) );
NOR2xp33_ASAP7_75t_R g689 ( .A(n_629), .B(n_636), .Y(n_689) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_629), .B(n_630), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_637), .A2(n_625), .B1(n_626), .B2(n_641), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_662), .B(n_642), .C(n_673), .Y(n_692) );
NAND4xp75_ASAP7_75t_L g693 ( .A(n_672), .B(n_654), .C(n_655), .D(n_640), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g694 ( .A1(n_661), .A2(n_651), .B(n_680), .C(n_640), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_630), .A2(n_667), .B(n_654), .C(n_639), .Y(n_695) );
AOI322xp5_ASAP7_75t_L g696 ( .A1(n_688), .A2(n_624), .A3(n_625), .B1(n_626), .B2(n_638), .C1(n_642), .C2(n_674), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_684), .A2(n_633), .B1(n_647), .B2(n_646), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_682), .A2(n_631), .B(n_648), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_690), .A2(n_671), .B1(n_634), .B2(n_643), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_683), .A2(n_658), .B(n_655), .C(n_656), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_684), .A2(n_644), .B1(n_645), .B2(n_664), .C(n_671), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_692), .Y(n_702) );
AOI22x1_ASAP7_75t_L g703 ( .A1(n_686), .A2(n_671), .B1(n_669), .B2(n_675), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_691), .B1(n_685), .B2(n_687), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_697), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_700), .B(n_695), .C(n_694), .Y(n_706) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_702), .B(n_689), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_699), .A2(n_645), .B1(n_632), .B2(n_635), .C(n_650), .Y(n_708) );
AOI22xp5_ASAP7_75t_SL g709 ( .A1(n_705), .A2(n_698), .B1(n_693), .B2(n_696), .Y(n_709) );
BUFx3_ASAP7_75t_L g710 ( .A(n_707), .Y(n_710) );
AO22x2_ASAP7_75t_L g711 ( .A1(n_706), .A2(n_701), .B1(n_635), .B2(n_632), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_710), .A2(n_704), .B1(n_708), .B2(n_666), .C(n_657), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_711), .A2(n_652), .B1(n_650), .B2(n_670), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_713), .A2(n_709), .B1(n_711), .B2(n_665), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_714), .Y(n_716) );
BUFx2_ASAP7_75t_SL g717 ( .A(n_716), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_715), .B(n_659), .Y(n_718) );
endmodule