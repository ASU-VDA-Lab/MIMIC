module real_jpeg_4732_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_366;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_1),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_1),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_1),
.A2(n_91),
.B1(n_104),
.B2(n_264),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_1),
.A2(n_91),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_2),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_50),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_50),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_3),
.A2(n_50),
.B1(n_272),
.B2(n_276),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_4),
.A2(n_37),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_4),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_4),
.A2(n_28),
.B1(n_85),
.B2(n_227),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_4),
.A2(n_85),
.B1(n_116),
.B2(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_4),
.A2(n_85),
.B1(n_295),
.B2(n_298),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_5),
.A2(n_157),
.B1(n_162),
.B2(n_166),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_5),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_5),
.A2(n_166),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_6),
.A2(n_46),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_6),
.B(n_257),
.C(n_260),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_6),
.B(n_72),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_6),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_6),
.B(n_251),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_6),
.B(n_333),
.Y(n_332)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_108),
.B1(n_110),
.B2(n_113),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_8),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_8),
.A2(n_113),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_9),
.Y(n_169)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_9),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_9),
.Y(n_270)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_9),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_9),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_10),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_10),
.Y(n_214)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_13),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_13),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_14),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_14),
.Y(n_174)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_15),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_15),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_15),
.Y(n_259)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_234),
.B1(n_235),
.B2(n_366),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_18),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_233),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_199),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_20),
.B(n_199),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_135),
.C(n_176),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_21),
.B(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_55),
.B2(n_134),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_22),
.B(n_56),
.C(n_95),
.Y(n_218)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_42),
.B(n_47),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_24),
.B(n_49),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_36),
.Y(n_334)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_41),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_42),
.A2(n_139),
.A3(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_138)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_46),
.CON(n_42),
.SN(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_46),
.B(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_46),
.A2(n_151),
.B(n_268),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_SL g327 ( 
.A1(n_46),
.A2(n_328),
.B(n_331),
.Y(n_327)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.Y(n_48)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_54),
.Y(n_198)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_95),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_56)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_57),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_72),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_67),
.B2(n_70),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_63),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_66),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_66),
.Y(n_185)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_72),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_75),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_76),
.Y(n_324)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_80),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_82),
.A2(n_86),
.B(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_86),
.B(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_87),
.Y(n_231)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_89),
.A2(n_332),
.A3(n_341),
.B1(n_344),
.B2(n_346),
.Y(n_340)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_90),
.Y(n_330)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_107),
.B(n_114),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_96),
.A2(n_107),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_96),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_96),
.A2(n_114),
.B(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_96),
.A2(n_203),
.B1(n_280),
.B2(n_319),
.Y(n_318)
);

AOI22x1_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_103),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_104),
.B(n_288),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_112),
.Y(n_245)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_112),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_115),
.B(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_123),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_132),
.Y(n_255)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_135),
.A2(n_136),
.B1(n_176),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_149),
.B2(n_150),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_138),
.B(n_149),
.Y(n_222)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_155),
.B1(n_167),
.B2(n_170),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_151),
.A2(n_263),
.B(n_268),
.Y(n_262)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_156),
.B1(n_188),
.B2(n_194),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_152),
.A2(n_171),
.B1(n_210),
.B2(n_216),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_152),
.B(n_271),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_152),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_154),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_158),
.Y(n_276)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_172),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_173),
.Y(n_267)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_176),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_187),
.C(n_197),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_177),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_186),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_186),
.A2(n_232),
.B(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_187),
.B(n_197),
.Y(n_357)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_188),
.Y(n_337)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_190),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_226),
.B(n_228),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_221),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_203),
.A2(n_242),
.B(n_250),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_203),
.A2(n_250),
.B(n_319),
.Y(n_354)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_208),
.Y(n_321)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_230),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_360),
.B(n_365),
.Y(n_235)
);

AO21x2_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_349),
.B(n_359),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_313),
.B(n_348),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_284),
.B(n_312),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_261),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_240),
.B(n_261),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_252),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_241),
.A2(n_252),
.B1(n_253),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_241),
.Y(n_310)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_249),
.Y(n_343)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_277),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_278),
.C(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_282),
.B2(n_283),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_303),
.B(n_311),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_292),
.B(n_302),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.Y(n_286)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_301),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_299),
.B(n_300),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_300),
.A2(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_309),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_309),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_308),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_315),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_335),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_325),
.B2(n_326),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_325),
.C(n_335),
.Y(n_350)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g346 ( 
.A(n_321),
.B(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_340),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_350),
.B(n_351),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_356),
.B2(n_358),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_355),
.C(n_358),
.Y(n_361)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_361),
.B(n_362),
.Y(n_365)
);


endmodule