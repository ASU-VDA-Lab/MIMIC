module fake_jpeg_11938_n_378 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_76),
.Y(n_90)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_27),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_64),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_74),
.Y(n_123)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_73),
.Y(n_104)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_18),
.B(n_12),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_42),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_0),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_9),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_21),
.B1(n_24),
.B2(n_33),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_85),
.A2(n_97),
.B1(n_117),
.B2(n_120),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_87),
.A2(n_89),
.B1(n_98),
.B2(n_112),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_34),
.B1(n_26),
.B2(n_32),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_88),
.A2(n_107),
.B1(n_122),
.B2(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_24),
.B1(n_26),
.B2(n_40),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_19),
.B1(n_20),
.B2(n_40),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_20),
.B1(n_17),
.B2(n_16),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_62),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_16),
.B(n_3),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_106),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_56),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_22),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_113),
.A2(n_114),
.B1(n_125),
.B2(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_44),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_72),
.A2(n_1),
.B(n_8),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_121),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_57),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_53),
.A2(n_10),
.B1(n_65),
.B2(n_66),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_81),
.B1(n_69),
.B2(n_73),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_60),
.A2(n_10),
.B1(n_58),
.B2(n_46),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_104),
.B1(n_100),
.B2(n_86),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_47),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_132),
.B(n_133),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_47),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_59),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_62),
.C(n_52),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_138),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_172),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_140),
.A2(n_164),
.B1(n_160),
.B2(n_155),
.Y(n_192)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_145),
.B1(n_147),
.B2(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_143),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_90),
.B(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_148),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_89),
.A2(n_86),
.B1(n_98),
.B2(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_105),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_119),
.B1(n_124),
.B2(n_94),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_121),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_150),
.B(n_157),
.Y(n_206)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_92),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_163),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_92),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_159),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_95),
.B(n_111),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_87),
.A2(n_95),
.B(n_119),
.C(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_110),
.B(n_91),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_175),
.B1(n_143),
.B2(n_165),
.Y(n_213)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_174),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_90),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_152),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_137),
.B(n_167),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_196),
.C(n_210),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_187),
.B(n_184),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_176),
.B(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_195),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_194),
.B1(n_197),
.B2(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_140),
.A2(n_145),
.B1(n_156),
.B2(n_147),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_147),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_145),
.A2(n_147),
.B1(n_168),
.B2(n_169),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_131),
.B1(n_170),
.B2(n_151),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_174),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_135),
.A2(n_149),
.B1(n_134),
.B2(n_141),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_217),
.B(n_219),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_154),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_228),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_149),
.B1(n_175),
.B2(n_172),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_230),
.B1(n_207),
.B2(n_202),
.Y(n_265)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_139),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_171),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_171),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_180),
.C(n_203),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_234),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_192),
.B1(n_195),
.B2(n_182),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_178),
.B(n_184),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_231),
.B(n_232),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_186),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_239),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_179),
.Y(n_237)
);

HB1xp67_ASAP7_75t_SL g269 ( 
.A(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_184),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_182),
.B1(n_211),
.B2(n_200),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_240),
.A2(n_225),
.B1(n_243),
.B2(n_241),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_182),
.B(n_200),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_196),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_199),
.B(n_183),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_185),
.C(n_212),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_210),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_232),
.Y(n_276)
);

AOI22x1_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_183),
.B1(n_212),
.B2(n_199),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_250),
.A2(n_262),
.B(n_266),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_253),
.B(n_234),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_191),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_261),
.C(n_264),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_270),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_191),
.B(n_185),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_215),
.C(n_207),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_225),
.B1(n_244),
.B2(n_246),
.Y(n_292)
);

OAI31xp33_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_235),
.A3(n_221),
.B(n_230),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_215),
.C(n_202),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_277),
.C(n_275),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_217),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_248),
.B1(n_238),
.B2(n_218),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_226),
.A2(n_236),
.B(n_243),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_224),
.B(n_237),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_274),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_216),
.C(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_279),
.A2(n_295),
.B1(n_265),
.B2(n_250),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_282),
.B(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_286),
.C(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_229),
.C(n_239),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_228),
.B(n_219),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_220),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_296),
.B(n_262),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_260),
.B1(n_250),
.B2(n_272),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_264),
.C(n_276),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_267),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_294),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_222),
.B1(n_223),
.B2(n_233),
.Y(n_295)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_233),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_268),
.C(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_263),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_254),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_298),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_254),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_252),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_312),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_297),
.C(n_281),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_309),
.B(n_300),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_252),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_281),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_266),
.B1(n_259),
.B2(n_251),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_288),
.A2(n_253),
.B(n_259),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_296),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_272),
.B1(n_288),
.B2(n_299),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_279),
.B1(n_291),
.B2(n_290),
.Y(n_324)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_286),
.C(n_285),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_330),
.C(n_327),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_327),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_335),
.B1(n_313),
.B2(n_306),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_325),
.A2(n_329),
.B(n_333),
.C(n_315),
.Y(n_342)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_326),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_319),
.B(n_280),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_303),
.C(n_305),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_331),
.A2(n_332),
.B(n_334),
.Y(n_343)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_287),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_333),
.A2(n_316),
.B1(n_307),
.B2(n_318),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_344),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_338),
.B(n_341),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_310),
.C(n_311),
.Y(n_341)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_342),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_308),
.C(n_309),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_347),
.C(n_322),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_302),
.C(n_306),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_347),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_356),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_287),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_354),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_339),
.A2(n_324),
.B1(n_312),
.B2(n_320),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_351),
.A2(n_333),
.B1(n_342),
.B2(n_304),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_325),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_339),
.B(n_301),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_355),
.B(n_301),
.Y(n_361)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_343),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_357),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_345),
.C(n_336),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_365),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_361),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_336),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_364),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_353),
.A2(n_317),
.B1(n_304),
.B2(n_283),
.Y(n_365)
);

NAND2x1_ASAP7_75t_SL g370 ( 
.A(n_362),
.B(n_353),
.Y(n_370)
);

AOI21xp33_ASAP7_75t_L g372 ( 
.A1(n_370),
.A2(n_360),
.B(n_364),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_367),
.B(n_359),
.C(n_352),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_373),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_372),
.Y(n_375)
);

AOI322xp5_ASAP7_75t_L g373 ( 
.A1(n_369),
.A2(n_332),
.A3(n_365),
.B1(n_348),
.B2(n_278),
.C1(n_356),
.C2(n_358),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_375),
.A2(n_366),
.B(n_368),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_374),
.B(n_370),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_377),
.Y(n_378)
);


endmodule