module fake_jpeg_16051_n_52 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_52);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_52;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_1),
.B1(n_2),
.B2(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_25),
.C(n_26),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_38),
.B(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_35),
.B2(n_37),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_45),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_33),
.Y(n_49)
);

AOI322xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_10),
.A3(n_11),
.B1(n_14),
.B2(n_15),
.C1(n_17),
.C2(n_18),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_20),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_21),
.C(n_24),
.Y(n_52)
);


endmodule