module real_jpeg_6084_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_1),
.A2(n_26),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_45),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_1),
.A2(n_45),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_1),
.A2(n_45),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_2),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_159),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_4),
.A2(n_159),
.B1(n_277),
.B2(n_280),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_4),
.A2(n_28),
.B1(n_159),
.B2(n_414),
.Y(n_413)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_6),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_6),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_6),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_6),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_6),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_12),
.A2(n_25),
.B1(n_137),
.B2(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_12),
.B(n_33),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_12),
.A2(n_25),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_12),
.A2(n_25),
.B1(n_39),
.B2(n_219),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_12),
.A2(n_302),
.B(n_305),
.C(n_309),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_12),
.B(n_122),
.C(n_164),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_12),
.B(n_111),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_12),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_12),
.B(n_127),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_13),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_13),
.A2(n_71),
.B1(n_107),
.B2(n_110),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_13),
.A2(n_71),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_13),
.A2(n_71),
.B1(n_131),
.B2(n_335),
.Y(n_334)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_437),
.Y(n_19)
);

OAI221xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_55),
.B1(n_59),
.B2(n_432),
.C(n_435),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_21),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_21),
.B(n_55),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_22),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_23),
.B(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_48),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_29),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_25),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_29),
.Y(n_152)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_33),
.B(n_44),
.Y(n_212)
);

AO22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_41),
.Y(n_33)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_34),
.Y(n_149)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_36),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_37),
.Y(n_220)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_38),
.Y(n_148)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_39),
.Y(n_309)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_40),
.Y(n_156)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_43),
.B(n_68),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_43),
.A2(n_57),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_48),
.B(n_69),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_51),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_53),
.B(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_55),
.A2(n_257),
.B1(n_262),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_55),
.A2(n_262),
.B(n_268),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B(n_58),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_56),
.A2(n_212),
.B(n_413),
.Y(n_428)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_392),
.B(n_422),
.C(n_425),
.D(n_431),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_384),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_245),
.C(n_291),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_221),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_194),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_64),
.B(n_194),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_143),
.C(n_179),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_65),
.B(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_73),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_66),
.B(n_74),
.C(n_113),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_67),
.B(n_212),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_112),
.B1(n_113),
.B2(n_142),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_105),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_76),
.A2(n_111),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_76),
.B(n_216),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_100),
.Y(n_76)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_77),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_90),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_83),
.B2(n_87),
.Y(n_78)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_80),
.Y(n_304)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_90),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_99),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_95),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_95),
.Y(n_318)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_98),
.Y(n_205)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_98),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_98),
.Y(n_317)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_101),
.B(n_111),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_102),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_105),
.B(n_255),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_106),
.B(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_111),
.A2(n_183),
.B(n_218),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_112),
.A2(n_113),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_112),
.B(n_399),
.C(n_402),
.Y(n_420)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_113),
.B(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_113),
.B(n_418),
.C(n_419),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_134),
.B(n_135),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_114),
.A2(n_202),
.B(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_115),
.B(n_136),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_115),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_115),
.B(n_314),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_127),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_122),
.B2(n_125),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_118),
.Y(n_308)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_127),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_127),
.B(n_314),
.Y(n_329)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_133),
.Y(n_127)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_131),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_134),
.A2(n_231),
.B(n_236),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_134),
.B(n_135),
.Y(n_284)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_143),
.A2(n_144),
.B1(n_179),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_157),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_145),
.B(n_157),
.Y(n_209)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.A3(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_148),
.Y(n_279)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_165),
.B(n_169),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_191),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_170),
.A2(n_188),
.B(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_170),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_171),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_172),
.Y(n_338)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_179),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_186),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_180),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_181),
.B(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_181),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_183),
.B(n_218),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_183),
.A2(n_276),
.B(n_403),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_186),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_187),
.B(n_350),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_191),
.B(n_333),
.Y(n_362)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_208),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_197),
.C(n_208),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_200),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_201),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_202),
.B(n_313),
.Y(n_340)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_205),
.Y(n_326)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_211),
.C(n_214),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_221),
.A2(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_244),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_222),
.B(n_244),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_223),
.B(n_225),
.C(n_237),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_237),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_230),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_227),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_229),
.B(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_236),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_236),
.B(n_329),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_240),
.B(n_428),
.C(n_429),
.Y(n_434)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_242),
.B(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_288),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_246),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_264),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_247),
.B(n_264),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.C(n_263),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_248),
.B(n_256),
.CI(n_263),
.CON(n_289),
.SN(n_289)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_253),
.C(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_261),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_257),
.A2(n_262),
.B1(n_301),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_287),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_273),
.B2(n_274),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_267),
.B(n_273),
.C(n_287),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_283),
.B(n_286),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_283),
.Y(n_286)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_286),
.A2(n_396),
.B1(n_397),
.B2(n_404),
.Y(n_395)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_286),
.Y(n_404)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_288),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_289),
.B(n_290),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g439 ( 
.A(n_289),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_319),
.B(n_383),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_293),
.B(n_296),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.C(n_310),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_297),
.B(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_300),
.A2(n_310),
.B1(n_311),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx11_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_377),
.B(n_382),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_367),
.B(n_376),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_344),
.B(n_366),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_330),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_330),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_325),
.B1(n_328),
.B2(n_347),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_339),
.Y(n_330)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_351),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_342),
.C(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_353),
.B(n_365),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_348),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_361),
.B(n_364),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_360),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_363),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_370),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_374),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_373),
.C(n_374),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_381),
.Y(n_382)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_386),
.B(n_389),
.C(n_390),
.D(n_391),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_407),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_406),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_406),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_405),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_404),
.C(n_405),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_398),
.A2(n_399),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_410),
.C(n_420),
.Y(n_430)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_407),
.A2(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_421),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_421),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_420),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_415),
.B1(n_416),
.B2(n_419),
.Y(n_411)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_412),
.Y(n_419)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_430),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_430),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_434),
.Y(n_436)
);


endmodule