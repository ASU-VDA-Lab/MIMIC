module fake_jpeg_22342_n_281 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_28),
.B1(n_18),
.B2(n_27),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_53),
.B1(n_39),
.B2(n_23),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_27),
.B(n_18),
.Y(n_44)
);

NAND2x1p5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_28),
.B1(n_27),
.B2(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_28),
.B1(n_16),
.B2(n_15),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_16),
.B1(n_17),
.B2(n_15),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_17),
.B1(n_26),
.B2(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_50),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_17),
.B1(n_26),
.B2(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_70),
.Y(n_90)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_66),
.Y(n_88)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_59),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_22),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_73),
.B(n_19),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_78),
.B1(n_81),
.B2(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_39),
.B1(n_23),
.B2(n_24),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_39),
.B1(n_19),
.B2(n_31),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_52),
.B1(n_54),
.B2(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_101),
.B1(n_69),
.B2(n_77),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_34),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_103),
.C(n_104),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_55),
.B1(n_38),
.B2(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_38),
.B1(n_49),
.B2(n_34),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_100),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_68),
.B1(n_65),
.B2(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_49),
.B(n_21),
.C(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_9),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_21),
.B1(n_36),
.B2(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_21),
.B1(n_36),
.B2(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_105),
.B(n_7),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_7),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_103),
.B1(n_101),
.B2(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_113),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_85),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_124),
.B1(n_127),
.B2(n_61),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_126),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_80),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_101),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_131),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_94),
.C(n_93),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_137),
.C(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_106),
.B1(n_116),
.B2(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_100),
.C(n_82),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_145),
.B(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_101),
.B1(n_67),
.B2(n_86),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_127),
.B1(n_112),
.B2(n_108),
.Y(n_160)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_141),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_101),
.C(n_36),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_143),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_99),
.B(n_86),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_92),
.C(n_14),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_14),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_155),
.B1(n_167),
.B2(n_174),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_120),
.B1(n_119),
.B2(n_109),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_139),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_147),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_172),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

INVxp33_ASAP7_75t_SL g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_105),
.B1(n_115),
.B2(n_108),
.Y(n_167)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_110),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_158),
.C(n_137),
.Y(n_189)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_110),
.B1(n_124),
.B2(n_114),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_114),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_185),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_161),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_139),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_133),
.B(n_148),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_195),
.C(n_164),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_196),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_151),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_132),
.C(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_161),
.B(n_157),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_180),
.B(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_209),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_197),
.A2(n_155),
.B1(n_157),
.B2(n_152),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_181),
.B1(n_180),
.B2(n_215),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_212),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_0),
.Y(n_231)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_213),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_189),
.C(n_195),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_196),
.B1(n_193),
.B2(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_220),
.B(n_1),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_2),
.C(n_3),
.Y(n_237)
);

BUFx12f_ASAP7_75t_SL g220 ( 
.A(n_200),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_183),
.C(n_185),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_5),
.C(n_8),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_224),
.A2(n_226),
.B1(n_211),
.B2(n_202),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_187),
.B1(n_129),
.B2(n_165),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_206),
.B1(n_198),
.B2(n_214),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_231),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_6),
.CI(n_12),
.CON(n_229),
.SN(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_9),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_230),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_222),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_238),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_239),
.C(n_221),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_224),
.B(n_2),
.CI(n_3),
.CON(n_238),
.SN(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_4),
.C(n_5),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_245),
.C(n_8),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_13),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_246),
.B(n_252),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_247),
.B(n_254),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_223),
.B(n_229),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_256),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_251),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_222),
.C(n_227),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_228),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_238),
.B1(n_244),
.B2(n_11),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_8),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_10),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_241),
.B1(n_243),
.B2(n_236),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_253),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_238),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_265),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_11),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_266),
.A2(n_271),
.B(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_269),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_13),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_274),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_275),
.B(n_258),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_276),
.C(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_280),
.B(n_262),
.Y(n_281)
);


endmodule