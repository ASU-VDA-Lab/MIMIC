module fake_jpeg_153_n_589 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_589);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_589;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_18),
.C(n_17),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_57),
.B(n_32),
.C(n_55),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_58),
.Y(n_159)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_61),
.Y(n_202)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_62),
.Y(n_168)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_64),
.B(n_68),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_65),
.B(n_71),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_67),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_70),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_20),
.B(n_17),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_73),
.Y(n_194)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_75),
.Y(n_171)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_76),
.Y(n_215)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_77),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_25),
.B(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_78),
.B(n_89),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_79),
.Y(n_218)
);

CKINVDCx9p33_ASAP7_75t_R g80 ( 
.A(n_21),
.Y(n_80)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

HAxp5_ASAP7_75t_SL g82 ( 
.A(n_21),
.B(n_0),
.CON(n_82),
.SN(n_82)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_2),
.B(n_3),
.Y(n_133)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_29),
.Y(n_84)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_86),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_30),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_91),
.Y(n_198)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_92),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_93),
.Y(n_205)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_20),
.B(n_15),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_109),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_96),
.Y(n_222)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_39),
.B(n_15),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_101),
.Y(n_139)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_39),
.B(n_15),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_39),
.B(n_0),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_112),
.B(n_114),
.Y(n_206)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g212 ( 
.A(n_117),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g213 ( 
.A(n_118),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_54),
.B(n_0),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_122),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_121),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_125),
.Y(n_165)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_54),
.B(n_2),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_38),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_54),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_127),
.A2(n_28),
.B1(n_8),
.B2(n_10),
.Y(n_204)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_34),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_129),
.B(n_136),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_36),
.B(n_55),
.C(n_32),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_131),
.A2(n_139),
.B(n_135),
.C(n_140),
.Y(n_256)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_28),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_132),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_133),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_58),
.A2(n_56),
.B1(n_52),
.B2(n_38),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_134),
.A2(n_148),
.B1(n_195),
.B2(n_211),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_70),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_143),
.B(n_169),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_84),
.A2(n_56),
.B1(n_52),
.B2(n_34),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_56),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_150),
.B(n_155),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_60),
.A2(n_36),
.B1(n_50),
.B2(n_44),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_151),
.A2(n_76),
.B1(n_104),
.B2(n_62),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_87),
.B(n_52),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_37),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_172),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_162),
.B(n_174),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_66),
.A2(n_26),
.B1(n_44),
.B2(n_40),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_166),
.A2(n_187),
.B1(n_213),
.B2(n_175),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_96),
.B(n_37),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_72),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_100),
.B(n_38),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_180),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_37),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_73),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_181),
.B(n_182),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_107),
.A2(n_25),
.B1(n_40),
.B2(n_35),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_111),
.A2(n_50),
.B1(n_35),
.B2(n_26),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_201),
.B1(n_210),
.B2(n_141),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_108),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_75),
.B(n_3),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_196),
.B(n_197),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_61),
.B(n_117),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_61),
.B(n_6),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_199),
.B(n_203),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_121),
.A2(n_28),
.B1(n_29),
.B2(n_8),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_117),
.B(n_6),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_159),
.B(n_169),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_118),
.B(n_7),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_132),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_11),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_209),
.B(n_216),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_97),
.A2(n_28),
.B1(n_12),
.B2(n_13),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_82),
.A2(n_28),
.B1(n_12),
.B2(n_13),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_11),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_115),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_219),
.A2(n_122),
.B1(n_13),
.B2(n_14),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_103),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_223),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_103),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_227),
.A2(n_231),
.B1(n_266),
.B2(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_150),
.Y(n_228)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_229),
.B(n_243),
.Y(n_321)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_160),
.A2(n_127),
.B1(n_63),
.B2(n_81),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_232),
.A2(n_241),
.B1(n_252),
.B2(n_304),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_152),
.A2(n_14),
.B1(n_165),
.B2(n_176),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_233),
.A2(n_254),
.B1(n_269),
.B2(n_295),
.Y(n_327)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_234),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_172),
.A2(n_180),
.B1(n_200),
.B2(n_184),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_235),
.A2(n_240),
.B1(n_265),
.B2(n_297),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_236),
.A2(n_277),
.B1(n_286),
.B2(n_243),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_237),
.Y(n_339)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_239),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_184),
.A2(n_185),
.B1(n_200),
.B2(n_208),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_242),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

AO22x1_ASAP7_75t_SL g246 ( 
.A1(n_206),
.A2(n_185),
.B1(n_152),
.B2(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_246),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_164),
.B(n_140),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_247),
.B(n_258),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_212),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_249),
.B(n_256),
.Y(n_360)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_250),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_151),
.A2(n_141),
.B1(n_214),
.B2(n_149),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_143),
.A2(n_207),
.B1(n_204),
.B2(n_217),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_153),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_255),
.B(n_268),
.Y(n_311)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_257),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_259),
.B(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_260),
.B(n_264),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_133),
.A2(n_131),
.B(n_132),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_261),
.A2(n_303),
.B(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_149),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_167),
.A2(n_222),
.B1(n_205),
.B2(n_130),
.Y(n_266)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

BUFx24_ASAP7_75t_L g348 ( 
.A(n_267),
.Y(n_348)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_146),
.A2(n_178),
.B1(n_163),
.B2(n_189),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_163),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_270),
.B(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_178),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_168),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_273),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_168),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_186),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_275),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_171),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_198),
.A2(n_130),
.B1(n_189),
.B2(n_221),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_179),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_278),
.Y(n_352)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_183),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_282),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_146),
.A2(n_222),
.B1(n_205),
.B2(n_167),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_218),
.A2(n_194),
.B1(n_193),
.B2(n_142),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_302),
.B1(n_306),
.B2(n_258),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_190),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_283),
.B(n_287),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_214),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_292),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_190),
.A2(n_221),
.B1(n_218),
.B2(n_145),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_157),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_157),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_138),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_145),
.A2(n_191),
.B(n_183),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_SL g316 ( 
.A(n_290),
.B(n_250),
.C(n_233),
.Y(n_316)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_161),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_298),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_142),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_301),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_144),
.A2(n_194),
.B1(n_193),
.B2(n_158),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_144),
.A2(n_215),
.B1(n_186),
.B2(n_177),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_137),
.B(n_215),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_192),
.B(n_156),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_158),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_147),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_156),
.A2(n_173),
.B1(n_192),
.B2(n_147),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_191),
.A2(n_177),
.B1(n_147),
.B2(n_173),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_156),
.A2(n_173),
.B1(n_192),
.B2(n_191),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_313),
.A2(n_323),
.B(n_318),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_316),
.B(n_279),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_322),
.B(n_316),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_251),
.A2(n_229),
.B1(n_254),
.B2(n_230),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_228),
.A2(n_231),
.B1(n_238),
.B2(n_248),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_325),
.A2(n_349),
.B1(n_356),
.B2(n_345),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_225),
.A2(n_238),
.B1(n_248),
.B2(n_251),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_331),
.B1(n_358),
.B2(n_361),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_225),
.A2(n_251),
.B1(n_260),
.B2(n_261),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_246),
.B(n_305),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_341),
.Y(n_373)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_294),
.A2(n_255),
.A3(n_236),
.B1(n_298),
.B2(n_284),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_343),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_253),
.B(n_244),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_245),
.B(n_246),
.C(n_262),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_347),
.C(n_321),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_253),
.B(n_256),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_289),
.Y(n_343)
);

AOI32xp33_ASAP7_75t_L g344 ( 
.A1(n_276),
.A2(n_272),
.A3(n_273),
.B1(n_226),
.B2(n_299),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_353),
.Y(n_372)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_345),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_270),
.B(n_271),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_227),
.A2(n_280),
.B1(n_281),
.B2(n_269),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_264),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_259),
.B(n_263),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_357),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_295),
.A2(n_265),
.B1(n_239),
.B2(n_234),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_283),
.B(n_288),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_293),
.A2(n_287),
.B1(n_300),
.B2(n_274),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g361 ( 
.A1(n_301),
.A2(n_275),
.B1(n_257),
.B2(n_268),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_242),
.A2(n_241),
.B1(n_187),
.B2(n_166),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_267),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_396),
.C(n_406),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_366),
.B(n_365),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_351),
.A2(n_334),
.B1(n_308),
.B2(n_307),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_367),
.A2(n_392),
.B(n_369),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_351),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_369),
.B(n_395),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_371),
.B(n_383),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_344),
.A2(n_313),
.B(n_338),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_378),
.B(n_372),
.Y(n_427)
);

NOR2x1_ASAP7_75t_L g443 ( 
.A(n_378),
.B(n_391),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_325),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_388),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_320),
.A2(n_327),
.B1(n_308),
.B2(n_307),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_327),
.A2(n_314),
.B1(n_326),
.B2(n_349),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_381),
.A2(n_370),
.B1(n_367),
.B2(n_364),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_319),
.Y(n_382)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_360),
.B(n_363),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_311),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_385),
.B(n_389),
.Y(n_428)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_387),
.B(n_373),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_309),
.B(n_329),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_335),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_329),
.B(n_309),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_397),
.Y(n_421)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_391),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_346),
.Y(n_393)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

AOI32xp33_ASAP7_75t_L g395 ( 
.A1(n_323),
.A2(n_322),
.A3(n_318),
.B1(n_312),
.B2(n_357),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_340),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_339),
.B(n_352),
.Y(n_397)
);

OA21x2_ASAP7_75t_L g398 ( 
.A1(n_314),
.A2(n_356),
.B(n_315),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_324),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_346),
.Y(n_399)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_401),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_342),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_350),
.A2(n_342),
.B1(n_354),
.B2(n_336),
.Y(n_402)
);

AOI22x1_ASAP7_75t_SL g410 ( 
.A1(n_402),
.A2(n_361),
.B1(n_324),
.B2(n_348),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_339),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_403),
.B(n_359),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_358),
.A2(n_352),
.B1(n_333),
.B2(n_310),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_330),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_383),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_317),
.B(n_310),
.C(n_359),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_415),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g448 ( 
.A1(n_410),
.A2(n_414),
.B(n_435),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_401),
.B(n_348),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_403),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_416),
.B(n_417),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_371),
.B(n_348),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_374),
.A2(n_348),
.B(n_378),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_420),
.A2(n_427),
.B(n_433),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_396),
.C(n_392),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_439),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_424),
.B(n_431),
.Y(n_466)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_405),
.Y(n_426)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_430),
.A2(n_398),
.B1(n_370),
.B2(n_400),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_385),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_434),
.B(n_413),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_389),
.A2(n_373),
.B(n_379),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_395),
.A2(n_402),
.B(n_366),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_443),
.B(n_382),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_388),
.B(n_377),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_398),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_390),
.B(n_394),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_441),
.B(n_377),
.Y(n_447)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_445),
.A2(n_462),
.B(n_432),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_429),
.A2(n_381),
.B1(n_370),
.B2(n_364),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_446),
.A2(n_465),
.B1(n_467),
.B2(n_472),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_447),
.B(n_457),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_368),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_454),
.C(n_474),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_406),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_409),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_455),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_397),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_456),
.B(n_477),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_426),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_458),
.A2(n_407),
.B1(n_436),
.B2(n_432),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_426),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_459),
.B(n_460),
.Y(n_505)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_437),
.A2(n_433),
.B(n_427),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_429),
.A2(n_376),
.B1(n_398),
.B2(n_384),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_414),
.A2(n_384),
.B1(n_399),
.B2(n_393),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_471),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_415),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_473),
.Y(n_498)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_418),
.Y(n_470)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_435),
.B(n_413),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_414),
.A2(n_416),
.B1(n_419),
.B2(n_412),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_417),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_443),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_421),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_423),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_423),
.B(n_428),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_479),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_443),
.C(n_420),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_482),
.C(n_493),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_451),
.B(n_408),
.C(n_418),
.Y(n_482)
);

A2O1A1Ixp33_ASAP7_75t_SL g483 ( 
.A1(n_460),
.A2(n_430),
.B(n_410),
.C(n_441),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_483),
.A2(n_484),
.B(n_494),
.Y(n_508)
);

O2A1O1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_445),
.A2(n_408),
.B(n_421),
.C(n_436),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_449),
.Y(n_485)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_485),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_449),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_497),
.Y(n_506)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_490),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_440),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_495),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_441),
.C(n_412),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_476),
.A2(n_432),
.B(n_425),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_425),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_496),
.A2(n_502),
.B(n_448),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_453),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_438),
.C(n_407),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_474),
.C(n_462),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_476),
.A2(n_407),
.B(n_438),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_453),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_504),
.B(n_459),
.Y(n_507)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_507),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_455),
.Y(n_509)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_520),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_478),
.B(n_475),
.C(n_472),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_517),
.C(n_526),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_514),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_501),
.A2(n_458),
.B1(n_469),
.B2(n_473),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_515),
.A2(n_465),
.B1(n_444),
.B2(n_483),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_450),
.C(n_461),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_450),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_503),
.Y(n_521)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_521),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_481),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_487),
.Y(n_536)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_503),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_524),
.A2(n_489),
.B1(n_501),
.B2(n_505),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_457),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_525),
.B(n_499),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_482),
.B(n_463),
.C(n_464),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_444),
.C(n_447),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_500),
.C(n_494),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_486),
.B(n_466),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_528),
.B(n_493),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_515),
.Y(n_530)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_530),
.Y(n_550)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_531),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_533),
.A2(n_535),
.B1(n_540),
.B2(n_542),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_521),
.A2(n_505),
.B1(n_446),
.B2(n_483),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_543),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_544),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_488),
.C(n_496),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_545),
.C(n_510),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_523),
.A2(n_485),
.B1(n_504),
.B2(n_479),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_448),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_502),
.C(n_480),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_546),
.A2(n_514),
.B(n_508),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_547),
.B(n_559),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_530),
.A2(n_524),
.B1(n_519),
.B2(n_508),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_548),
.A2(n_549),
.B1(n_553),
.B2(n_541),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_519),
.B1(n_509),
.B2(n_506),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_551),
.B(n_552),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_534),
.B(n_526),
.C(n_512),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_538),
.A2(n_506),
.B1(n_525),
.B2(n_507),
.Y(n_553)
);

AO221x1_ASAP7_75t_L g557 ( 
.A1(n_540),
.A2(n_484),
.B1(n_527),
.B2(n_520),
.C(n_483),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_557),
.A2(n_538),
.B1(n_545),
.B2(n_535),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_529),
.C(n_539),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_529),
.C(n_537),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_546),
.A2(n_448),
.B(n_483),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_561),
.B(n_562),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_556),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_556),
.Y(n_563)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_563),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_564),
.A2(n_565),
.B1(n_570),
.B2(n_555),
.Y(n_572)
);

BUFx24_ASAP7_75t_SL g568 ( 
.A(n_560),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_568),
.B(n_549),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_511),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_569),
.A2(n_566),
.B(n_570),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_558),
.B(n_550),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_571),
.A2(n_572),
.B1(n_541),
.B2(n_518),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_563),
.B(n_548),
.C(n_554),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_575),
.B(n_554),
.C(n_543),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_547),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_567),
.B(n_553),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_577),
.B(n_516),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_578),
.B(n_579),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_580),
.A2(n_581),
.B(n_575),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_583),
.B(n_559),
.C(n_536),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_579),
.B(n_573),
.C(n_574),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_516),
.Y(n_585)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_585),
.A2(n_586),
.B(n_582),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_518),
.C(n_513),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_588),
.B(n_513),
.Y(n_589)
);


endmodule