module fake_jpeg_14847_n_303 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_14;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_0),
.C(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_33),
.Y(n_43)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_46),
.Y(n_51)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_27),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_31),
.B1(n_34),
.B2(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_55),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_36),
.B1(n_35),
.B2(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_21),
.B1(n_20),
.B2(n_17),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_34),
.B1(n_28),
.B2(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_60),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_34),
.B1(n_28),
.B2(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_33),
.B1(n_29),
.B2(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_67),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_33),
.B(n_29),
.C(n_15),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_29),
.B1(n_18),
.B2(n_15),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_46),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_18),
.B1(n_23),
.B2(n_13),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_20),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_74),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_89),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_48),
.C(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_61),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_42),
.B1(n_46),
.B2(n_66),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_59),
.Y(n_97)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_86),
.B(n_71),
.Y(n_125)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_52),
.B1(n_50),
.B2(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_110),
.B1(n_82),
.B2(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_64),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_53),
.B1(n_63),
.B2(n_54),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_112),
.B(n_79),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_135),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_81),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_121),
.C(n_111),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_81),
.C(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_83),
.B(n_85),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_79),
.B(n_104),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_71),
.B(n_86),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_53),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_92),
.Y(n_143)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_108),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_146),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_155),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_70),
.Y(n_148)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_78),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_78),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_53),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_157),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_57),
.C(n_110),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_134),
.B1(n_131),
.B2(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_78),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_110),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_161),
.B(n_55),
.Y(n_187)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_126),
.B(n_124),
.Y(n_168)
);

XOR2x1_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_125),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_168),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_127),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_174),
.B(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_122),
.B1(n_121),
.B2(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_113),
.B1(n_104),
.B2(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

NOR4xp25_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_148),
.C(n_147),
.D(n_150),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_128),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_179),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_138),
.B1(n_137),
.B2(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_155),
.A2(n_104),
.B(n_133),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_186),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_137),
.A2(n_94),
.B1(n_130),
.B2(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_94),
.B(n_87),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_95),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_210),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_144),
.C(n_154),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_194),
.C(n_196),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_152),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_144),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_58),
.C(n_45),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_202),
.C(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_58),
.C(n_145),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_185),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_68),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_208),
.C(n_209),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_66),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_65),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_166),
.B(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_187),
.B1(n_188),
.B2(n_172),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_217),
.B1(n_20),
.B2(n_22),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_206),
.B(n_176),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_9),
.B(n_12),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_173),
.B1(n_169),
.B2(n_180),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_174),
.C(n_186),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_219),
.C(n_223),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_177),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_170),
.B1(n_182),
.B2(n_101),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_170),
.B(n_12),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_48),
.C(n_45),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_197),
.B1(n_205),
.B2(n_200),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_13),
.B1(n_19),
.B2(n_16),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_225),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_48),
.C(n_37),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_37),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_46),
.B1(n_42),
.B2(n_41),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_233),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_41),
.B1(n_40),
.B2(n_2),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_237),
.B1(n_244),
.B2(n_40),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_41),
.B1(n_40),
.B2(n_2),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_37),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_0),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_23),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_240),
.B(n_247),
.Y(n_248)
);

OAI321xp33_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_69),
.A3(n_18),
.B1(n_11),
.B2(n_10),
.C(n_6),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_219),
.C(n_227),
.Y(n_257)
);

AOI21x1_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_37),
.B(n_40),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_218),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_253),
.C(n_256),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_26),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_211),
.C(n_212),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_217),
.B(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_211),
.C(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_214),
.B1(n_229),
.B2(n_22),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_259),
.B1(n_17),
.B2(n_13),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_214),
.B1(n_22),
.B2(n_17),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_236),
.C(n_234),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_265),
.C(n_267),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_273),
.B1(n_19),
.B2(n_16),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_244),
.C(n_231),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_25),
.Y(n_267)
);

XOR2x1_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_11),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_248),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_1),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_251),
.B(n_261),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.C(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_252),
.C(n_24),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_281),
.C(n_282),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_26),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_25),
.C(n_26),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_14),
.B(n_6),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_270),
.C(n_14),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_10),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_266),
.C(n_25),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.C(n_8),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_10),
.C(n_9),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_274),
.B1(n_6),
.B2(n_3),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_284),
.C(n_288),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_293),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_285),
.C(n_295),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_5),
.C(n_3),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_3),
.C(n_4),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_4),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_4),
.C(n_5),
.Y(n_303)
);


endmodule