module fake_jpeg_17981_n_154 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_154);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_29),
.B1(n_26),
.B2(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_54),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_32),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_24),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_22),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_66),
.C(n_68),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_15),
.C(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_46),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_76),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_23),
.B(n_21),
.C(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_50),
.B1(n_48),
.B2(n_46),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_52),
.B1(n_59),
.B2(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_49),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_64),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_88),
.B(n_95),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_44),
.C(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_93),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_55),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_96),
.B1(n_75),
.B2(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_1),
.B(n_3),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_16),
.B1(n_11),
.B2(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_73),
.C(n_78),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_79),
.Y(n_107)
);

XOR2x1_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_60),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_95),
.B(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_66),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_88),
.B(n_81),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_117),
.B(n_127),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_71),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_92),
.B1(n_97),
.B2(n_71),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_126),
.B1(n_104),
.B2(n_100),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_125),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_97),
.B1(n_71),
.B2(n_85),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_84),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_107),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_132),
.B(n_106),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_98),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_115),
.B1(n_126),
.B2(n_127),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

AOI321xp33_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_124),
.A3(n_120),
.B1(n_116),
.B2(n_111),
.C(n_69),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_128),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_137),
.C(n_139),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_133),
.C(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_138),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_142),
.A2(n_70),
.B1(n_63),
.B2(n_67),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_146),
.C(n_147),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_105),
.B(n_63),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_72),
.B1(n_4),
.B2(n_5),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_146),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_148),
.C(n_142),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_8),
.B(n_72),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_8),
.Y(n_154)
);


endmodule