module fake_jpeg_1385_n_610 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_610);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_610;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_62),
.B(n_70),
.Y(n_134)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_19),
.B(n_10),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_10),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_71),
.B(n_121),
.Y(n_158)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_79),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_35),
.A2(n_10),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_81),
.B(n_83),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_9),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_88),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_89),
.Y(n_215)
);

HAxp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_0),
.CON(n_90),
.SN(n_90)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_90),
.B(n_104),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_36),
.C(n_44),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_91),
.A2(n_25),
.B(n_31),
.Y(n_172)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_94),
.Y(n_204)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_98),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_101),
.Y(n_151)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_11),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g197 ( 
.A(n_106),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_11),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_116),
.B(n_117),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_11),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

BUFx4f_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_23),
.B(n_11),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_122),
.Y(n_191)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

BUFx4f_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_48),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_130),
.A2(n_107),
.B1(n_58),
.B2(n_52),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_68),
.A2(n_25),
.B1(n_31),
.B2(n_57),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_135),
.A2(n_155),
.B1(n_160),
.B2(n_175),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_137),
.B(n_138),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_73),
.A2(n_27),
.B1(n_23),
.B2(n_33),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_77),
.A2(n_25),
.B1(n_31),
.B2(n_57),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_27),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_171),
.B(n_179),
.Y(n_227)
);

NAND2x1_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_124),
.Y(n_229)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_85),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_41),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_88),
.B(n_41),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_82),
.B(n_43),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_189),
.B(n_14),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_190),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_120),
.A2(n_46),
.B1(n_48),
.B2(n_34),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_SL g255 ( 
.A1(n_193),
.A2(n_194),
.B(n_210),
.C(n_1),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_125),
.A2(n_46),
.B1(n_37),
.B2(n_49),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_89),
.B(n_43),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_76),
.B(n_49),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_63),
.A2(n_58),
.B1(n_52),
.B2(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_60),
.Y(n_213)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_65),
.Y(n_217)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_217),
.Y(n_280)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_219),
.Y(n_329)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_220),
.Y(n_309)
);

AO22x1_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_90),
.B1(n_114),
.B2(n_111),
.Y(n_222)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_224),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_177),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_225),
.B(n_229),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_228),
.Y(n_318)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_153),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_230),
.Y(n_295)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_232),
.Y(n_319)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_233),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_136),
.B(n_87),
.C(n_96),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_234),
.B(n_251),
.C(n_265),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_186),
.A2(n_114),
.B1(n_111),
.B2(n_98),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_235),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_140),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_236),
.B(n_259),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_237),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_186),
.A2(n_52),
.B1(n_50),
.B2(n_122),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_238),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_140),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_239),
.B(n_278),
.Y(n_304)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_240),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_244),
.A2(n_249),
.B1(n_252),
.B2(n_267),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_150),
.A2(n_50),
.B1(n_39),
.B2(n_12),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_168),
.Y(n_250)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_250),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_150),
.B(n_9),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_135),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_252)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_255),
.A2(n_152),
.B1(n_161),
.B2(n_142),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_158),
.B(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_258),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_2),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_199),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_148),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_262),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_130),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_261),
.A2(n_290),
.B1(n_153),
.B2(n_145),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_144),
.B(n_3),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_146),
.B(n_3),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_263),
.B(n_269),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_149),
.Y(n_264)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

OR2x2_ASAP7_75t_SL g265 ( 
.A(n_134),
.B(n_13),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_266),
.B(n_279),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_160),
.A2(n_5),
.B1(n_8),
.B2(n_12),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_154),
.B(n_3),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_185),
.C(n_204),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_134),
.B(n_141),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g270 ( 
.A1(n_177),
.A2(n_5),
.B1(n_12),
.B2(n_16),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_270),
.A2(n_283),
.B(n_252),
.Y(n_338)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_139),
.Y(n_271)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_187),
.Y(n_273)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_131),
.B(n_5),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_270),
.Y(n_335)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_212),
.Y(n_275)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_275),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_190),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_170),
.B(n_17),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_132),
.B(n_17),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_285),
.Y(n_308)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_178),
.Y(n_282)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

AO22x1_ASAP7_75t_L g283 ( 
.A1(n_143),
.A2(n_17),
.B1(n_18),
.B2(n_147),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_161),
.Y(n_284)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_284),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_202),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_191),
.A2(n_18),
.B(n_194),
.C(n_166),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_286),
.B(n_163),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_202),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_225),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_208),
.Y(n_288)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_129),
.Y(n_289)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_210),
.A2(n_18),
.B1(n_193),
.B2(n_196),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_129),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_292),
.Y(n_326)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_151),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_151),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_293),
.B(n_294),
.Y(n_351)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_192),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_301),
.A2(n_314),
.B1(n_340),
.B2(n_244),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_226),
.A2(n_165),
.B1(n_184),
.B2(n_142),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_315),
.A2(n_328),
.B(n_238),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_247),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_324),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_268),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_327),
.B(n_293),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_332),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_260),
.B(n_269),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_334),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_335),
.B(n_231),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_226),
.B(n_181),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_344),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_248),
.A2(n_209),
.B1(n_183),
.B2(n_215),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_337),
.A2(n_341),
.B1(n_230),
.B2(n_284),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_227),
.A2(n_159),
.B1(n_176),
.B2(n_157),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_248),
.A2(n_209),
.B1(n_215),
.B2(n_169),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_268),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_220),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_262),
.B(n_157),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_263),
.B(n_173),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_346),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_274),
.B(n_173),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_258),
.B(n_197),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_379),
.Y(n_415)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_348),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_335),
.A2(n_251),
.B(n_256),
.C(n_286),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_355),
.B(n_383),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_328),
.A2(n_229),
.B(n_255),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_356),
.A2(n_378),
.B(n_382),
.Y(n_403)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_358),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_359),
.A2(n_363),
.B1(n_395),
.B2(n_297),
.Y(n_396)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_253),
.C(n_234),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_365),
.C(n_369),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_350),
.A2(n_255),
.B1(n_243),
.B2(n_294),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_221),
.C(n_222),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_222),
.C(n_280),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_370),
.Y(n_397)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_349),
.Y(n_373)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_376),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_299),
.A2(n_283),
.B1(n_255),
.B2(n_275),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_377),
.A2(n_393),
.B1(n_327),
.B2(n_295),
.Y(n_414)
);

A2O1A1O1Ixp25_ASAP7_75t_L g378 ( 
.A1(n_299),
.A2(n_265),
.B(n_230),
.C(n_273),
.D(n_241),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_380),
.B(n_387),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_321),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_394),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_250),
.B(n_254),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_297),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_389),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_297),
.A2(n_245),
.B(n_246),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_388),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_320),
.B(n_308),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_306),
.A2(n_197),
.B1(n_214),
.B2(n_183),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_392),
.B1(n_340),
.B2(n_303),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_317),
.B(n_277),
.C(n_272),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_276),
.C(n_323),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_306),
.A2(n_214),
.B1(n_169),
.B2(n_207),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_338),
.A2(n_149),
.B1(n_207),
.B2(n_240),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_321),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_388),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_404),
.B(n_431),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_370),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_422),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_305),
.C(n_310),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_419),
.C(n_429),
.Y(n_436)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_391),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_412),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_368),
.A2(n_311),
.B1(n_342),
.B2(n_324),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_413),
.A2(n_381),
.B1(n_383),
.B2(n_357),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_414),
.A2(n_361),
.B1(n_389),
.B2(n_390),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_298),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_371),
.B(n_336),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_377),
.A2(n_345),
.B1(n_344),
.B2(n_346),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_421),
.A2(n_425),
.B1(n_393),
.B2(n_352),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_298),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_369),
.A2(n_365),
.B1(n_356),
.B2(n_367),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_384),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_325),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_305),
.C(n_304),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_379),
.C(n_384),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_367),
.B(n_310),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_361),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_432),
.B(n_442),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_403),
.A2(n_358),
.B(n_382),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_433),
.A2(n_435),
.B(n_448),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_403),
.A2(n_378),
.B(n_355),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_437),
.A2(n_447),
.B1(n_430),
.B2(n_420),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_420),
.B(n_353),
.Y(n_438)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_438),
.Y(n_472)
);

AOI32xp33_ASAP7_75t_L g439 ( 
.A1(n_400),
.A2(n_380),
.A3(n_378),
.B1(n_372),
.B2(n_376),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_440),
.B(n_443),
.C(n_462),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_406),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_386),
.C(n_323),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_395),
.Y(n_444)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_444),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_421),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_415),
.A2(n_392),
.B1(n_311),
.B2(n_394),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_415),
.A2(n_408),
.B(n_428),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_399),
.Y(n_450)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_452),
.A2(n_459),
.B1(n_416),
.B2(n_402),
.Y(n_481)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_453),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_413),
.A2(n_354),
.B(n_325),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_454),
.A2(n_424),
.B(n_406),
.Y(n_470)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_461),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_457),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_360),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_458),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_415),
.A2(n_303),
.B1(n_318),
.B2(n_373),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_417),
.B(n_333),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_224),
.Y(n_488)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_405),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_417),
.B(n_333),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_375),
.Y(n_463)
);

XNOR2x2_ASAP7_75t_SL g466 ( 
.A(n_463),
.B(n_419),
.Y(n_466)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_464),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_465),
.A2(n_467),
.B1(n_468),
.B2(n_476),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_460),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_437),
.A2(n_411),
.B1(n_427),
.B2(n_409),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_434),
.A2(n_409),
.B1(n_425),
.B2(n_414),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_470),
.A2(n_474),
.B(n_495),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_398),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_478),
.Y(n_499)
);

A2O1A1Ixp33_ASAP7_75t_SL g474 ( 
.A1(n_433),
.A2(n_452),
.B(n_434),
.C(n_439),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_493),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_448),
.A2(n_410),
.B1(n_397),
.B2(n_407),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_435),
.A2(n_432),
.B1(n_446),
.B2(n_438),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_477),
.A2(n_480),
.B1(n_486),
.B2(n_494),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_398),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_445),
.A2(n_397),
.B1(n_424),
.B2(n_416),
.Y(n_480)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_481),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_441),
.A2(n_426),
.B1(n_402),
.B2(n_429),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_312),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_488),
.Y(n_508)
);

OA22x2_ASAP7_75t_L g493 ( 
.A1(n_450),
.A2(n_426),
.B1(n_366),
.B2(n_318),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_441),
.A2(n_426),
.B1(n_339),
.B2(n_296),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_454),
.A2(n_300),
.B(n_331),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_496),
.B(n_443),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_457),
.Y(n_500)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_500),
.Y(n_529)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_489),
.Y(n_503)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_503),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_436),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_506),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_482),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_507),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_436),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_482),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_472),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_511),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_473),
.B(n_440),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_510),
.B(n_513),
.Y(n_541)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_485),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_478),
.B(n_440),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_512),
.B(n_518),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_462),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_466),
.B(n_462),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_487),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_480),
.A2(n_447),
.B1(n_442),
.B2(n_459),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_516),
.B1(n_519),
.B2(n_484),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_467),
.A2(n_463),
.B1(n_453),
.B2(n_456),
.Y(n_516)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_490),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_468),
.A2(n_444),
.B1(n_455),
.B2(n_451),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_469),
.B(n_458),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_520),
.B(n_494),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_483),
.A2(n_464),
.B1(n_461),
.B2(n_460),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_521),
.A2(n_477),
.B1(n_486),
.B2(n_483),
.Y(n_525)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_495),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_523),
.A2(n_534),
.B1(n_543),
.B2(n_508),
.Y(n_551)
);

XOR2x2_ASAP7_75t_L g547 ( 
.A(n_525),
.B(n_526),
.Y(n_547)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_527),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_479),
.C(n_488),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_536),
.C(n_538),
.Y(n_550)
);

AOI21x1_ASAP7_75t_L g533 ( 
.A1(n_517),
.A2(n_479),
.B(n_470),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_498),
.A2(n_465),
.B1(n_481),
.B2(n_474),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_535),
.B(n_540),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_499),
.B(n_513),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_542),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_499),
.B(n_474),
.Y(n_538)
);

XNOR2x1_ASAP7_75t_L g540 ( 
.A(n_517),
.B(n_474),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_514),
.B(n_493),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_502),
.A2(n_493),
.B1(n_339),
.B2(n_331),
.Y(n_543)
);

OAI221xp5_ASAP7_75t_L g544 ( 
.A1(n_531),
.A2(n_519),
.B1(n_497),
.B2(n_516),
.C(n_502),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_544),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_532),
.B(n_504),
.Y(n_545)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_545),
.Y(n_561)
);

AOI221xp5_ASAP7_75t_L g546 ( 
.A1(n_524),
.A2(n_521),
.B1(n_497),
.B2(n_501),
.C(n_515),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_546),
.A2(n_554),
.B1(n_555),
.B2(n_309),
.Y(n_568)
);

OAI221xp5_ASAP7_75t_L g548 ( 
.A1(n_529),
.A2(n_506),
.B1(n_496),
.B2(n_508),
.C(n_501),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_548),
.A2(n_525),
.B1(n_538),
.B2(n_526),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_551),
.A2(n_219),
.B1(n_228),
.B2(n_264),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_493),
.C(n_300),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_552),
.B(n_557),
.C(n_560),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_527),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_539),
.B(n_319),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_536),
.C(n_528),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_530),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_558),
.A2(n_309),
.B1(n_242),
.B2(n_257),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_312),
.C(n_343),
.Y(n_560)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_562),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_553),
.A2(n_543),
.B1(n_534),
.B2(n_540),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_563),
.A2(n_565),
.B1(n_568),
.B2(n_569),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_559),
.A2(n_542),
.B1(n_537),
.B2(n_330),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_550),
.B(n_343),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_566),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_SL g567 ( 
.A(n_549),
.B(n_330),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_573),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_570),
.B(n_572),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_560),
.B(n_322),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_556),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_551),
.A2(n_302),
.B1(n_319),
.B2(n_307),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_574),
.B(n_552),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_564),
.B(n_557),
.C(n_550),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_575),
.B(n_581),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_579),
.B(n_583),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_564),
.B(n_547),
.C(n_556),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_571),
.B(n_558),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_582),
.B(n_584),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_547),
.C(n_559),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_561),
.B(n_302),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_562),
.A2(n_271),
.B(n_322),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_585),
.A2(n_565),
.B(n_569),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_575),
.B(n_573),
.C(n_563),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_588),
.B(n_586),
.Y(n_599)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_590),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_572),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_595),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_567),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_593),
.A2(n_594),
.B(n_586),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_581),
.A2(n_307),
.B(n_289),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_578),
.Y(n_595)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_596),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_587),
.B(n_577),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_L g603 ( 
.A(n_597),
.B(n_591),
.C(n_589),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_599),
.B(n_600),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_589),
.A2(n_233),
.B1(n_282),
.B2(n_288),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_603),
.A2(n_601),
.B(n_598),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_605),
.B(n_606),
.Y(n_607)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_604),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_607),
.A2(n_602),
.B(n_600),
.Y(n_608)
);

AOI21x1_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_593),
.B(n_291),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_609),
.A2(n_292),
.B(n_232),
.Y(n_610)
);


endmodule