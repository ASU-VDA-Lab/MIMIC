module fake_jpeg_25751_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_19),
.B1(n_32),
.B2(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_40),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_43),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_54),
.B1(n_56),
.B2(n_44),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_30),
.B1(n_23),
.B2(n_24),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_20),
.B1(n_32),
.B2(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_30),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_21),
.B1(n_34),
.B2(n_25),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_58),
.B1(n_66),
.B2(n_44),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_34),
.B1(n_25),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_33),
.B1(n_28),
.B2(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_33),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_33),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_90),
.C(n_43),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_26),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.Y(n_94)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_44),
.B1(n_28),
.B2(n_33),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_26),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_62),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_107),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_67),
.A3(n_66),
.B1(n_40),
.B2(n_39),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_62),
.B(n_39),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_114),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_116),
.Y(n_120)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_40),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_53),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_49),
.C(n_47),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_125),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_80),
.B1(n_77),
.B2(n_90),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_137),
.B1(n_96),
.B2(n_93),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_73),
.A3(n_80),
.B1(n_68),
.B2(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_139),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_85),
.B1(n_62),
.B2(n_89),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_140),
.B1(n_44),
.B2(n_39),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_85),
.B1(n_82),
.B2(n_65),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_162),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_112),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_154),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_96),
.B1(n_93),
.B2(n_98),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_132),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_95),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_17),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_96),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_79),
.B(n_91),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_127),
.B(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_164),
.B1(n_167),
.B2(n_114),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_43),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_65),
.B1(n_107),
.B2(n_74),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_101),
.B1(n_74),
.B2(n_87),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_87),
.B1(n_115),
.B2(n_47),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_124),
.A2(n_123),
.B1(n_138),
.B2(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_174),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_171),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_17),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_167),
.B1(n_158),
.B2(n_144),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_165),
.B1(n_147),
.B2(n_144),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_128),
.C(n_72),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_182),
.C(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_180),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_103),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_72),
.C(n_53),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_53),
.C(n_17),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_186),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_103),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_189),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_187),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_151),
.B1(n_159),
.B2(n_28),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_197),
.B1(n_207),
.B2(n_175),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_145),
.B(n_154),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_205),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_187),
.B1(n_186),
.B2(n_181),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_183),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_149),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_208),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_143),
.C(n_156),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_204),
.C(n_181),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_143),
.C(n_157),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_155),
.Y(n_205)
);

XNOR2x2_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_178),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_173),
.C(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_224),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_173),
.C(n_34),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_202),
.B(n_25),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_203),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_191),
.B1(n_198),
.B2(n_199),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_205),
.B(n_221),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_217),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_234),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_209),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_221),
.A2(n_199),
.B1(n_207),
.B2(n_193),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_236),
.A2(n_223),
.B(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_3),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_23),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g242 ( 
.A(n_235),
.B(n_225),
.C(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_22),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_3),
.C(n_4),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_246),
.C(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_5),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_4),
.C(n_5),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_231),
.B(n_227),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_254),
.B(n_7),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_227),
.B(n_236),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_256),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_246),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_261),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_245),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_260),
.Y(n_266)
);

AOI221xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_252),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_252),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_7),
.C2(n_12),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_265),
.B1(n_258),
.B2(n_11),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_10),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_249),
.C2(n_251),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_268),
.Y(n_271)
);


endmodule