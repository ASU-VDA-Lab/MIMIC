module real_jpeg_23611_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx6_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_0),
.Y(n_120)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_4),
.A2(n_41),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_4),
.B(n_31),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_68),
.C(n_84),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_4),
.B(n_52),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_4),
.A2(n_106),
.B1(n_223),
.B2(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_6),
.A2(n_32),
.B1(n_35),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_6),
.A2(n_46),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_6),
.A2(n_46),
.B1(n_67),
.B2(n_68),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_7),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_7),
.A2(n_27),
.B1(n_32),
.B2(n_35),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_7),
.A2(n_27),
.B1(n_53),
.B2(n_54),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_7),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_8),
.A2(n_67),
.B1(n_68),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_77),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_73),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_11),
.A2(n_67),
.B1(n_68),
.B2(n_91),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_11),
.A2(n_32),
.B1(n_35),
.B2(n_91),
.Y(n_139)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_14),
.A2(n_32),
.B1(n_35),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_14),
.A2(n_57),
.B1(n_67),
.B2(n_68),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_15),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_15),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_15),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_15),
.A2(n_40),
.B1(n_67),
.B2(n_68),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_145),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_143),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_19),
.B(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_78),
.C(n_100),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_20),
.B(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_58),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_23),
.B(n_43),
.C(n_58),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_31),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_24),
.Y(n_99)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_29),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_29),
.A2(n_31),
.B1(n_39),
.B2(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_37),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_30),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_95)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_36),
.B(n_60),
.C(n_63),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g172 ( 
.A(n_32),
.B(n_61),
.CON(n_172),
.SN(n_172)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_35),
.C(n_62),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_35),
.A2(n_51),
.A3(n_54),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_41),
.Y(n_133)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_55),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_47),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_47),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_47),
.A2(n_93),
.B1(n_94),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_48),
.A2(n_52),
.B1(n_162),
.B2(n_172),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_50),
.B(n_53),
.Y(n_173)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_52),
.B(n_139),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_54),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_54),
.B(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_61),
.B(n_87),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_61),
.B(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_66),
.B(n_109),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_66),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_68),
.B1(n_84),
.B2(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_67),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_70),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_72),
.A2(n_122),
.B(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_78),
.A2(n_79),
.B1(n_100),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_92),
.C(n_95),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_80),
.A2(n_81),
.B1(n_92),
.B2(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_88),
.B(n_89),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_82),
.A2(n_125),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_82),
.A2(n_179),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_82),
.A2(n_125),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_82),
.A2(n_125),
.B1(n_178),
.B2(n_199),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_87),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_88),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_95),
.B(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_100),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_105),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_108),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_106),
.A2(n_108),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_106),
.A2(n_118),
.B(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_106),
.A2(n_214),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_141),
.B2(n_142),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_128),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_123),
.B2(n_127),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_140),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_247),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_166),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_163),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_149),
.B(n_163),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_150),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_153),
.B(n_155),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_184),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_242),
.B(n_246),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_193),
.B(n_241),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_180),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_169),
.B(n_180),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.C(n_177),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_174),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_176),
.B(n_177),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_188),
.C(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_192),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_187),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_236),
.B(n_240),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_210),
.B(n_235),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_202),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_200),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_219),
.B(n_234),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_218),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_226),
.B(n_233),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_237),
.B(n_238),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);


endmodule