module fake_netlist_5_490_n_158 (n_29, n_16, n_0, n_12, n_9, n_36, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_34, n_4, n_32, n_35, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_158);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_36;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_34;
input n_4;
input n_32;
input n_35;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_158;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_76;
wire n_87;
wire n_150;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_104;
wire n_41;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_6),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_75),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_58),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_60),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_44),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

AO21x2_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_96),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_118),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_113),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_111),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_7),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_8),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_35),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_130),
.B(n_129),
.C(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_141),
.C(n_127),
.Y(n_143)
);

OAI221xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_16),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_146),
.Y(n_147)
);

AO22x2_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_34),
.B1(n_21),
.B2(n_22),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_153),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_29),
.Y(n_157)
);

AOI211xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_158)
);


endmodule