module fake_jpeg_23879_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_7),
.B(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_6),
.B(n_7),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_15),
.B1(n_24),
.B2(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_14),
.B1(n_24),
.B2(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_14),
.B1(n_24),
.B2(n_22),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_44),
.B(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_29),
.B1(n_31),
.B2(n_15),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_49),
.B1(n_56),
.B2(n_63),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_57),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_51),
.C(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_60),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_23),
.Y(n_51)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_19),
.A3(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_23),
.C(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_67),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_17),
.B1(n_27),
.B2(n_20),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_1),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_47),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_92),
.Y(n_100)
);

XNOR2x1_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_54),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_83),
.C(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_49),
.B1(n_77),
.B2(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_56),
.B1(n_46),
.B2(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_62),
.B1(n_59),
.B2(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_2),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_92),
.B1(n_70),
.B2(n_86),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_69),
.A3(n_68),
.B1(n_79),
.B2(n_81),
.C1(n_72),
.C2(n_71),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.C(n_88),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_84),
.B(n_82),
.C(n_73),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_90),
.B1(n_87),
.B2(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_85),
.C(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_113),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_85),
.C(n_91),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_102),
.C(n_96),
.Y(n_117)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_102),
.A3(n_107),
.B1(n_101),
.B2(n_99),
.C(n_97),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_121),
.B(n_111),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_102),
.B(n_97),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_110),
.B1(n_111),
.B2(n_71),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_122),
.A2(n_123),
.B(n_125),
.C(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_16),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_3),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_117),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.C(n_9),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_130),
.B(n_9),
.Y(n_132)
);

OAI31xp33_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_5),
.A3(n_6),
.B(n_9),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_131),
.A2(n_132),
.B(n_10),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_10),
.B(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_10),
.Y(n_135)
);


endmodule