module fake_jpeg_2240_n_525 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_13),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_54),
.Y(n_158)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_55),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_48),
.Y(n_120)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_37),
.Y(n_130)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_102),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_32),
.B1(n_47),
.B2(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_104),
.A2(n_113),
.B1(n_116),
.B2(n_135),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_47),
.B1(n_32),
.B2(n_50),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_48),
.B1(n_25),
.B2(n_33),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_115),
.A2(n_31),
.B1(n_29),
.B2(n_2),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_47),
.B1(n_39),
.B2(n_19),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_19),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_138),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_130),
.B(n_150),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_62),
.B1(n_72),
.B2(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_24),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_51),
.A2(n_71),
.B1(n_58),
.B2(n_60),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_159),
.B1(n_165),
.B2(n_31),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_54),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_128),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_50),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_73),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_68),
.B(n_37),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_84),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_78),
.A2(n_22),
.B1(n_21),
.B2(n_35),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_169),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_33),
.B1(n_35),
.B2(n_77),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_171),
.A2(n_181),
.B1(n_184),
.B2(n_190),
.Y(n_268)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_192),
.C(n_202),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_175),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_194),
.Y(n_231)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_100),
.B1(n_97),
.B2(n_96),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_113),
.A2(n_92),
.B1(n_86),
.B2(n_31),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_182),
.A2(n_185),
.B1(n_115),
.B2(n_137),
.Y(n_250)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_31),
.B1(n_29),
.B2(n_2),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_127),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_196),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_0),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_199),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_112),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_1),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_207),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_105),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_229),
.B(n_132),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_112),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_108),
.B(n_1),
.Y(n_207)
);

BUFx4f_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_213),
.B(n_216),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_162),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_215),
.B(n_220),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_218),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_109),
.B(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_221),
.B(n_222),
.Y(n_281)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

INVx3_ASAP7_75t_SL g223 ( 
.A(n_128),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_224),
.Y(n_267)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_133),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_137),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_230),
.B1(n_110),
.B2(n_104),
.Y(n_232)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_208),
.B1(n_210),
.B2(n_200),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_111),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_232),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_159),
.B1(n_121),
.B2(n_129),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_233),
.A2(n_247),
.B1(n_250),
.B2(n_259),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_184),
.A2(n_139),
.B1(n_134),
.B2(n_158),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_182),
.A2(n_177),
.B1(n_176),
.B2(n_196),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_263),
.B1(n_280),
.B2(n_187),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_174),
.A2(n_139),
.B1(n_134),
.B2(n_143),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_188),
.B(n_131),
.C(n_166),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_273),
.C(n_277),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_203),
.A2(n_29),
.B1(n_5),
.B2(n_6),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_170),
.A2(n_228),
.B1(n_198),
.B2(n_186),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_274),
.B1(n_195),
.B2(n_220),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_198),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_7),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_178),
.B(n_3),
.C(n_5),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_179),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_180),
.B(n_7),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_183),
.A2(n_191),
.B1(n_208),
.B2(n_223),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_251),
.A2(n_212),
.B1(n_219),
.B2(n_201),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_284),
.A2(n_297),
.B1(n_303),
.B2(n_282),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_286),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_288),
.A2(n_293),
.B1(n_294),
.B2(n_308),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_289),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_241),
.B(n_172),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_290),
.B(n_321),
.Y(n_333)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_231),
.B(n_189),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_292),
.B(n_298),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_218),
.B1(n_199),
.B2(n_217),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_247),
.A2(n_216),
.B(n_169),
.C(n_227),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_295),
.A2(n_296),
.B(n_306),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_248),
.A2(n_230),
.B(n_224),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_227),
.B1(n_10),
.B2(n_12),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_275),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_236),
.A2(n_9),
.B(n_12),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_301),
.A2(n_269),
.B(n_263),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_268),
.A2(n_281),
.B1(n_240),
.B2(n_265),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_237),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_304),
.Y(n_363)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_243),
.A2(n_271),
.B(n_235),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_259),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_233),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_309),
.A2(n_316),
.B1(n_300),
.B2(n_287),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_15),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_310),
.B(n_313),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_16),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_322),
.Y(n_342)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_267),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_274),
.A2(n_16),
.B1(n_256),
.B2(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_258),
.Y(n_317)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_254),
.Y(n_318)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_318),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_280),
.A2(n_232),
.B1(n_264),
.B2(n_234),
.Y(n_320)
);

AO21x2_ASAP7_75t_SL g332 ( 
.A1(n_320),
.A2(n_232),
.B(n_262),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_238),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_246),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_264),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_325),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_238),
.B(n_255),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_324),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_266),
.B(n_252),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_327),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_246),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_260),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_253),
.C(n_252),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_339),
.C(n_348),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_285),
.B(n_253),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_283),
.A2(n_239),
.B(n_232),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_296),
.B(n_322),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_323),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_343),
.B(n_365),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_239),
.C(n_278),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_302),
.A2(n_234),
.B1(n_282),
.B2(n_278),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_349),
.A2(n_358),
.B1(n_288),
.B2(n_284),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_353),
.B1(n_357),
.B2(n_366),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_299),
.A2(n_261),
.B1(n_249),
.B2(n_257),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_261),
.C(n_249),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_348),
.C(n_337),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_299),
.A2(n_257),
.B1(n_245),
.B2(n_273),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_287),
.A2(n_293),
.B1(n_294),
.B2(n_313),
.Y(n_358)
);

NOR3xp33_ASAP7_75t_SL g359 ( 
.A(n_292),
.B(n_245),
.C(n_301),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_364),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_325),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_290),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_383),
.C(n_391),
.Y(n_401)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_346),
.A2(n_320),
.B1(n_314),
.B2(n_316),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_372),
.A2(n_384),
.B1(n_385),
.B2(n_396),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_298),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_373),
.B(n_380),
.Y(n_420)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_374),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_375),
.Y(n_424)
);

XNOR2x1_ASAP7_75t_L g376 ( 
.A(n_329),
.B(n_320),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_376),
.B(n_338),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_388),
.Y(n_414)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_334),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_390),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_367),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_352),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_382),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_327),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_346),
.A2(n_320),
.B1(n_300),
.B2(n_309),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_343),
.A2(n_295),
.B1(n_289),
.B2(n_312),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_342),
.Y(n_388)
);

AOI322xp5_ASAP7_75t_L g390 ( 
.A1(n_335),
.A2(n_311),
.A3(n_319),
.B1(n_326),
.B2(n_307),
.C1(n_317),
.C2(n_297),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_330),
.B(n_291),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_333),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_397),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_335),
.B(n_304),
.C(n_318),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_361),
.C(n_345),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_330),
.B(n_315),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_355),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_332),
.A2(n_286),
.B1(n_341),
.B2(n_340),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_333),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_400),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_363),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_351),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_425),
.Y(n_436)
);

AOI22x1_ASAP7_75t_L g405 ( 
.A1(n_386),
.A2(n_332),
.B1(n_358),
.B2(n_349),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_405),
.A2(n_422),
.B1(n_427),
.B2(n_389),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_382),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_406),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_386),
.A2(n_332),
.B1(n_340),
.B2(n_350),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_408),
.A2(n_372),
.B1(n_368),
.B2(n_371),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_429),
.C(n_392),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_379),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_396),
.A2(n_331),
.B1(n_353),
.B2(n_345),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_423),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_361),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_426),
.B(n_389),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_387),
.A2(n_336),
.B1(n_363),
.B2(n_360),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_356),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_388),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_376),
.C(n_394),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_414),
.Y(n_430)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_430),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_433),
.C(n_441),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_432),
.A2(n_444),
.B1(n_422),
.B2(n_405),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_429),
.B(n_391),
.C(n_373),
.Y(n_433)
);

AND2x2_ASAP7_75t_SL g435 ( 
.A(n_424),
.B(n_398),
.Y(n_435)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_438),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_439),
.B(n_442),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_409),
.Y(n_440)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_440),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_379),
.C(n_395),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_416),
.A2(n_377),
.B1(n_393),
.B2(n_400),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_450),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_385),
.Y(n_445)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_404),
.B(n_384),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_451),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_354),
.C(n_336),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_403),
.C(n_411),
.Y(n_467)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_420),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_449),
.B(n_453),
.Y(n_463)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_416),
.A2(n_359),
.B1(n_360),
.B2(n_354),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_424),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_415),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_SL g454 ( 
.A1(n_438),
.A2(n_408),
.B(n_405),
.C(n_419),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_454),
.A2(n_471),
.B(n_452),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_435),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_468),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_401),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_467),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_461),
.A2(n_437),
.B1(n_445),
.B2(n_450),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_428),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_436),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_435),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_432),
.A2(n_417),
.B1(n_407),
.B2(n_410),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_470),
.Y(n_475)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_431),
.C(n_447),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_477),
.Y(n_494)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_446),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_481),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_451),
.C(n_441),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_483),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_443),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_439),
.C(n_440),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_485),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_409),
.C(n_426),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_472),
.A2(n_418),
.B1(n_412),
.B2(n_430),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_487),
.Y(n_493)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_470),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_488),
.A2(n_462),
.B(n_471),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_427),
.B1(n_434),
.B2(n_413),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_489),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_456),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_488),
.A2(n_475),
.B1(n_460),
.B2(n_478),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_492),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_479),
.C(n_482),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_483),
.A2(n_462),
.B(n_460),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_498),
.B(n_469),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_455),
.C(n_473),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_457),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_484),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_504),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_499),
.B(n_480),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_485),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_506),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_481),
.C(n_473),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_508),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_469),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_510),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_503),
.A2(n_497),
.B1(n_496),
.B2(n_493),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_511),
.A2(n_490),
.B(n_498),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_496),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_517),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_506),
.C(n_501),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_512),
.C(n_514),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_519),
.C(n_511),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_521),
.A2(n_495),
.B(n_510),
.Y(n_522)
);

O2A1O1Ixp33_ASAP7_75t_SL g523 ( 
.A1(n_522),
.A2(n_457),
.B(n_454),
.C(n_442),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_454),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_454),
.Y(n_525)
);


endmodule