module real_jpeg_13916_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_16;

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_3),
.B(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_13),
.B1(n_22),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_27),
.B1(n_44),
.B2(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_3),
.B(n_13),
.C(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_5),
.A2(n_13),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_23),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_13),
.B1(n_22),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_6),
.A2(n_32),
.B1(n_44),
.B2(n_46),
.Y(n_73)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_60),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_39),
.B(n_59),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_28),
.B(n_38),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_19),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_16),
.Y(n_12)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_18),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_22),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_17),
.B(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_24),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_31),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_35),
.B(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_37),
.B1(n_44),
.B2(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_56),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_50),
.Y(n_74)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_46),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_83),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_64),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_82),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);


endmodule