module fake_jpeg_465_n_543 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_543);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx2_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_119),
.Y(n_132)
);

CKINVDCx9p33_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g141 ( 
.A(n_58),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_23),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_59),
.B(n_73),
.Y(n_137)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_61),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_64),
.Y(n_179)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_67),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_75),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_82),
.A2(n_11),
.B1(n_86),
.B2(n_112),
.Y(n_197)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_85),
.Y(n_135)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_86),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_87),
.B(n_94),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_92),
.B(n_99),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_93),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_34),
.B(n_15),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_15),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_97),
.B(n_100),
.Y(n_165)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_15),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_101),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_102),
.B(n_103),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_16),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_25),
.A2(n_13),
.B1(n_7),
.B2(n_8),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_106),
.A2(n_82),
.B1(n_44),
.B2(n_38),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_108),
.A2(n_115),
.B(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_109),
.B(n_114),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_20),
.B(n_13),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_50),
.B(n_2),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_32),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_123),
.Y(n_139)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_50),
.B(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_44),
.Y(n_149)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_2),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_53),
.C(n_40),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_131),
.B(n_132),
.C(n_151),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_47),
.B1(n_28),
.B2(n_40),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_140),
.A2(n_142),
.B1(n_150),
.B2(n_151),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_93),
.B1(n_57),
.B2(n_95),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_45),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_145),
.B(n_161),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_47),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_146),
.B(n_149),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_70),
.A2(n_47),
.B1(n_28),
.B2(n_40),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_62),
.A2(n_47),
.B1(n_53),
.B2(n_40),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_107),
.A2(n_20),
.B1(n_30),
.B2(n_37),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_152),
.A2(n_162),
.B1(n_171),
.B2(n_200),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_66),
.A2(n_53),
.B1(n_31),
.B2(n_37),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_154),
.A2(n_163),
.B1(n_167),
.B2(n_172),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_SL g156 ( 
.A(n_65),
.Y(n_156)
);

CKINVDCx9p33_ASAP7_75t_R g252 ( 
.A(n_156),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_79),
.B(n_36),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_111),
.A2(n_30),
.B1(n_53),
.B2(n_31),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_68),
.A2(n_31),
.B1(n_49),
.B2(n_46),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_31),
.B1(n_49),
.B2(n_46),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_71),
.A2(n_32),
.B1(n_45),
.B2(n_27),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_67),
.A2(n_44),
.B1(n_38),
.B2(n_27),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_175),
.A2(n_178),
.B1(n_195),
.B2(n_197),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_67),
.A2(n_38),
.B1(n_52),
.B2(n_32),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_7),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_183),
.B(n_186),
.Y(n_280)
);

NAND2xp67_ASAP7_75t_SL g184 ( 
.A(n_122),
.B(n_52),
.Y(n_184)
);

OR2x2_ASAP7_75t_SL g240 ( 
.A(n_184),
.B(n_131),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_88),
.B(n_7),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_77),
.B(n_8),
.Y(n_188)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_188),
.B(n_192),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_84),
.B(n_8),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_85),
.A2(n_52),
.B1(n_9),
.B2(n_10),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_193),
.A2(n_135),
.B1(n_191),
.B2(n_159),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_83),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_89),
.B(n_9),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_120),
.A2(n_11),
.B1(n_91),
.B2(n_110),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_64),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_141),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_110),
.A2(n_11),
.B1(n_90),
.B2(n_108),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_108),
.A2(n_11),
.B1(n_113),
.B2(n_121),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_205),
.A2(n_210),
.B1(n_212),
.B2(n_145),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_58),
.A2(n_55),
.B1(n_104),
.B2(n_56),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_209),
.A2(n_211),
.B1(n_203),
.B2(n_175),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_113),
.A2(n_121),
.B1(n_116),
.B2(n_24),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_58),
.A2(n_55),
.B1(n_104),
.B2(n_56),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_113),
.A2(n_121),
.B1(n_116),
.B2(n_24),
.Y(n_212)
);

BUFx4f_ASAP7_75t_SL g218 ( 
.A(n_141),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_218),
.Y(n_327)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_129),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_129),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_223),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_160),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_224),
.B(n_225),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_146),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_226),
.B(n_261),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_132),
.B(n_142),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_227),
.A2(n_262),
.B(n_255),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_228),
.B(n_237),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_229),
.Y(n_304)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_141),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_230),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_137),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_233),
.B(n_235),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_234),
.B(n_248),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_194),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_184),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_150),
.A2(n_140),
.B1(n_178),
.B2(n_143),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_239),
.A2(n_244),
.B1(n_247),
.B2(n_254),
.Y(n_308)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_242),
.A2(n_246),
.B1(n_275),
.B2(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_139),
.B(n_147),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_243),
.B(n_259),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_133),
.A2(n_138),
.B1(n_148),
.B2(n_169),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_177),
.A2(n_209),
.B1(n_211),
.B2(n_195),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_179),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_128),
.Y(n_250)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_128),
.B(n_174),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_251),
.B(n_255),
.C(n_240),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_179),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_253),
.B(n_258),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_127),
.A2(n_215),
.B1(n_136),
.B2(n_191),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_130),
.B(n_136),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_135),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_155),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_153),
.B(n_190),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_189),
.B(n_158),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_264),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_172),
.B(n_206),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_130),
.B(n_168),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_189),
.B(n_202),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_155),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_269),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_202),
.B(n_199),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_213),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_278),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_273),
.B1(n_237),
.B2(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_197),
.A2(n_159),
.B1(n_213),
.B2(n_176),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_127),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_277),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_215),
.A2(n_197),
.B1(n_181),
.B2(n_134),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_157),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_134),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_181),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_187),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_187),
.B(n_207),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_207),
.B(n_180),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_129),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_156),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_287),
.Y(n_319)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_288),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_204),
.B(n_165),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_289),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_158),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_156),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_252),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_295),
.A2(n_312),
.B1(n_221),
.B2(n_229),
.Y(n_377)
);

OAI32xp33_ASAP7_75t_L g296 ( 
.A1(n_226),
.A2(n_228),
.A3(n_232),
.B1(n_261),
.B2(n_284),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_320),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g355 ( 
.A1(n_303),
.A2(n_331),
.B(n_285),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_232),
.B(n_266),
.C(n_280),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_305),
.B(n_337),
.C(n_303),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_227),
.B(n_290),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_330),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_265),
.A2(n_263),
.B1(n_245),
.B2(n_273),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_257),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_270),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_262),
.A2(n_267),
.B(n_246),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_322),
.A2(n_218),
.B(n_276),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_217),
.B(n_255),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_332),
.Y(n_363)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_239),
.B(n_265),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_267),
.A2(n_275),
.B1(n_254),
.B2(n_258),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_248),
.B(n_253),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_272),
.B(n_236),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_336),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_244),
.B(n_278),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_251),
.B(n_281),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_294),
.B(n_251),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_340),
.B(n_341),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_332),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_344),
.B(n_347),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_323),
.B(n_250),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_345),
.B(n_354),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_282),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_346),
.B(n_372),
.C(n_376),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_317),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_308),
.A2(n_271),
.B1(n_231),
.B2(n_268),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_349),
.A2(n_359),
.B1(n_360),
.B2(n_377),
.Y(n_412)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_322),
.A2(n_292),
.B(n_287),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_352),
.A2(n_374),
.B(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_333),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_355),
.A2(n_361),
.B(n_373),
.Y(n_386)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_313),
.Y(n_356)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

A2O1A1Ixp33_ASAP7_75t_SL g358 ( 
.A1(n_312),
.A2(n_252),
.B(n_218),
.C(n_230),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_358),
.A2(n_316),
.B(n_361),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_308),
.A2(n_274),
.B1(n_219),
.B2(n_220),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_330),
.A2(n_288),
.B1(n_286),
.B2(n_229),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_366),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_297),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_371),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_249),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_369),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_370),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_297),
.B(n_277),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_279),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_315),
.A2(n_241),
.B(n_242),
.Y(n_374)
);

AOI32xp33_ASAP7_75t_L g375 ( 
.A1(n_307),
.A2(n_256),
.A3(n_238),
.B1(n_291),
.B2(n_221),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_379),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_293),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_296),
.B(n_324),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_305),
.B(n_293),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_349),
.A2(n_295),
.B1(n_314),
.B2(n_319),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_383),
.Y(n_436)
);

NOR2x1_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_324),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_385),
.A2(n_388),
.B(n_400),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_387),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_359),
.A2(n_319),
.B1(n_325),
.B2(n_338),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_306),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_396),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_342),
.B(n_339),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_352),
.A2(n_311),
.B(n_306),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_365),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_408),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_377),
.A2(n_302),
.B1(n_329),
.B2(n_337),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_403),
.A2(n_348),
.B1(n_358),
.B2(n_362),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_326),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_367),
.C(n_376),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_301),
.B(n_327),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_321),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_357),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_343),
.A2(n_334),
.B(n_300),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_357),
.Y(n_421)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_414),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_403),
.A2(n_360),
.B1(n_350),
.B2(n_363),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_416),
.A2(n_435),
.B1(n_439),
.B2(n_440),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_406),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_434),
.Y(n_446)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_393),
.Y(n_419)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_419),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_409),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_425),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_299),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_432),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_389),
.B(n_371),
.Y(n_427)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_346),
.Y(n_428)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_428),
.Y(n_457)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_394),
.Y(n_429)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

BUFx12_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_430),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_431),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_298),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_437),
.C(n_390),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_343),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_411),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_372),
.C(n_363),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_398),
.B(n_370),
.Y(n_438)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_438),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_356),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_394),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_441),
.A2(n_442),
.B1(n_443),
.B2(n_391),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_353),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_396),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_416),
.A2(n_443),
.B1(n_435),
.B2(n_436),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_445),
.A2(n_450),
.B1(n_418),
.B2(n_452),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_436),
.A2(n_413),
.B1(n_412),
.B2(n_402),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_454),
.C(n_455),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_381),
.C(n_390),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_385),
.C(n_400),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_385),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_461),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_386),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_386),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_466),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_428),
.C(n_380),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_465),
.C(n_469),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_380),
.C(n_382),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_392),
.Y(n_466)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_392),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_467),
.B(n_424),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_471),
.B(n_477),
.Y(n_500)
);

OAI321xp33_ASAP7_75t_L g472 ( 
.A1(n_453),
.A2(n_421),
.A3(n_423),
.B1(n_439),
.B2(n_425),
.C(n_427),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_472),
.A2(n_474),
.B1(n_480),
.B2(n_485),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_466),
.B(n_398),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_473),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_447),
.A2(n_441),
.B1(n_418),
.B2(n_423),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_382),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_399),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_482),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_422),
.C(n_408),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_483),
.C(n_455),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_405),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_446),
.B(n_454),
.C(n_461),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_458),
.A2(n_412),
.B1(n_442),
.B2(n_387),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_484),
.A2(n_487),
.B1(n_450),
.B2(n_459),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_453),
.B(n_440),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_486),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_458),
.A2(n_414),
.B1(n_429),
.B2(n_419),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_457),
.B(n_397),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_449),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_445),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_493),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_492),
.B(n_495),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_446),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_465),
.C(n_464),
.Y(n_495)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_499),
.A2(n_501),
.B1(n_480),
.B2(n_474),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_476),
.A2(n_462),
.B1(n_448),
.B2(n_456),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_502),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_503),
.B(n_407),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_476),
.A2(n_397),
.B1(n_407),
.B2(n_358),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_504),
.B(n_486),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_508),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_499),
.A2(n_484),
.B(n_472),
.Y(n_506)
);

OAI21x1_ASAP7_75t_SL g522 ( 
.A1(n_506),
.A2(n_510),
.B(n_496),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_475),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_490),
.A2(n_488),
.B(n_481),
.Y(n_510)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_500),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_512),
.B(n_493),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_516),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_501),
.A2(n_470),
.B(n_483),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_514),
.A2(n_492),
.B(n_470),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_515),
.B(n_498),
.Y(n_517)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_517),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_502),
.Y(n_518)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_518),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_478),
.B(n_507),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_495),
.Y(n_521)
);

AO21x1_ASAP7_75t_L g532 ( 
.A1(n_521),
.A2(n_522),
.B(n_525),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_506),
.A2(n_497),
.B1(n_491),
.B2(n_410),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_517),
.C(n_524),
.Y(n_528)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_518),
.Y(n_526)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_526),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_528),
.B(n_530),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_520),
.A2(n_511),
.B(n_510),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_529),
.B(n_505),
.Y(n_533)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_533),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_532),
.B(n_491),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_535),
.B(n_526),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_538),
.A2(n_536),
.B(n_351),
.Y(n_541)
);

AOI322xp5_ASAP7_75t_L g539 ( 
.A1(n_534),
.A2(n_531),
.A3(n_527),
.B1(n_430),
.B2(n_410),
.C1(n_478),
.C2(n_304),
.Y(n_539)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_539),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_541),
.A2(n_537),
.B(n_338),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_540),
.Y(n_543)
);


endmodule