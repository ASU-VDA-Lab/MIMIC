module fake_netlist_6_4475_n_1089 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1089);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1089;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_842;
wire n_720;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_844;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_816;
wire n_743;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_1082;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_6),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_77),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_136),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_12),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_18),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_21),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_41),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_47),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_72),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_108),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_70),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_103),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_170),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_35),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_36),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_105),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_104),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_94),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_150),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_119),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_106),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_133),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_155),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_11),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_145),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_83),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_120),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_5),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_101),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_179),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_54),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_31),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_109),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_21),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_164),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_91),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_59),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_97),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_95),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_84),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_51),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_74),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_29),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_25),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_18),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_98),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_57),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_174),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_121),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_71),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_157),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_73),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_163),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_213),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g279 ( 
.A(n_218),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_215),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_262),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g284 ( 
.A(n_209),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_246),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_274),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_206),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_220),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_238),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_225),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_274),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_226),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_238),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

INVx4_ASAP7_75t_R g310 ( 
.A(n_256),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_233),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_239),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_224),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_243),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_266),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_257),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_304),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_279),
.A2(n_243),
.B1(n_264),
.B2(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_301),
.A2(n_261),
.B1(n_270),
.B2(n_268),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

CKINVDCx6p67_ASAP7_75t_R g331 ( 
.A(n_321),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_207),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_210),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_271),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_282),
.A2(n_267),
.B1(n_263),
.B2(n_259),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_258),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

AOI22x1_ASAP7_75t_SL g350 ( 
.A1(n_306),
.A2(n_255),
.B1(n_252),
.B2(n_250),
.Y(n_350)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

BUFx8_ASAP7_75t_L g354 ( 
.A(n_277),
.Y(n_354)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_313),
.A2(n_316),
.B(n_280),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_288),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_306),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_277),
.B(n_288),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_280),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_211),
.Y(n_365)
);

OAI21x1_ASAP7_75t_L g366 ( 
.A1(n_289),
.A2(n_231),
.B(n_221),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_286),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_289),
.B(n_292),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_212),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_284),
.A2(n_249),
.B1(n_247),
.B2(n_245),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_281),
.Y(n_373)
);

BUFx12f_ASAP7_75t_L g374 ( 
.A(n_281),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_275),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_374),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_333),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_374),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_331),
.Y(n_383)
);

INVxp33_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_323),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_323),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_361),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_331),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_350),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_348),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_354),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_354),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_330),
.B(n_307),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_354),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_285),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_R g398 ( 
.A(n_359),
.B(n_312),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_360),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_R g401 ( 
.A(n_359),
.B(n_312),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_373),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_365),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_343),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_337),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_337),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_341),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_351),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_324),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_351),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_R g416 ( 
.A(n_369),
.B(n_318),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_329),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_342),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_346),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_328),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_340),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_345),
.B(n_290),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_352),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_357),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_375),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_368),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_339),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_349),
.B(n_290),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_363),
.B(n_284),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_347),
.B(n_222),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_349),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_349),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_349),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_370),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_370),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_440),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_443),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_408),
.B(n_223),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_444),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_410),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_L g455 ( 
.A1(n_403),
.A2(n_287),
.B1(n_295),
.B2(n_314),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_384),
.B(n_283),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_347),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_406),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_404),
.B(n_367),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_429),
.B(n_227),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_413),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_397),
.B(n_228),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_295),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_415),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_347),
.Y(n_467)
);

INVx3_ASAP7_75t_R g468 ( 
.A(n_381),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_430),
.B(n_229),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_431),
.B(n_230),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_370),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_426),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_428),
.B(n_237),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

OAI22xp33_ASAP7_75t_L g486 ( 
.A1(n_392),
.A2(n_314),
.B1(n_292),
.B2(n_244),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_292),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_366),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_417),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_332),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_419),
.B(n_332),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_425),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_445),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_401),
.B(n_364),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_419),
.Y(n_503)
);

BUFx6f_ASAP7_75t_SL g504 ( 
.A(n_394),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_434),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_383),
.Y(n_506)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_382),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_420),
.B(n_240),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_434),
.B(n_364),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_434),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_434),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_411),
.B(n_366),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_390),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_399),
.B(n_364),
.Y(n_515)
);

INVx4_ASAP7_75t_SL g516 ( 
.A(n_389),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_421),
.B(n_310),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_416),
.B(n_353),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_418),
.B(n_353),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_386),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_387),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_395),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_396),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_R g527 ( 
.A(n_388),
.B(n_22),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_391),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_447),
.Y(n_529)
);

AO22x2_ASAP7_75t_L g530 ( 
.A1(n_525),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_453),
.B(n_0),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_513),
.A2(n_358),
.B1(n_336),
.B2(n_335),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_485),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_460),
.Y(n_535)
);

AOI211xp5_ASAP7_75t_L g536 ( 
.A1(n_455),
.A2(n_358),
.B(n_336),
.C(n_335),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_469),
.Y(n_537)
);

BUFx6f_ASAP7_75t_SL g538 ( 
.A(n_454),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_452),
.B(n_1),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_513),
.A2(n_520),
.B1(n_493),
.B2(n_492),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_456),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_471),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_477),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_458),
.B(n_338),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_494),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_454),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_489),
.A2(n_338),
.B1(n_4),
.B2(n_5),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_459),
.B(n_23),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_462),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_464),
.B(n_338),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_457),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_465),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_448),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_482),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_478),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_522),
.A2(n_450),
.B1(n_517),
.B2(n_497),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_482),
.B(n_24),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_508),
.B(n_3),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_490),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_469),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_490),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_479),
.B(n_26),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_467),
.B(n_3),
.Y(n_568)
);

OR2x6_ASAP7_75t_SL g569 ( 
.A(n_526),
.B(n_7),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_515),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_461),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_491),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_466),
.Y(n_575)
);

AO22x2_ASAP7_75t_L g576 ( 
.A1(n_522),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_27),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_502),
.B(n_470),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_474),
.B(n_8),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_451),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_473),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_473),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_512),
.B(n_476),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_511),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_501),
.B(n_9),
.Y(n_588)
);

OR2x2_ASAP7_75t_SL g589 ( 
.A(n_468),
.B(n_10),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_503),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_487),
.B(n_10),
.Y(n_592)
);

BUFx6f_ASAP7_75t_SL g593 ( 
.A(n_507),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_546),
.A2(n_472),
.B(n_481),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_563),
.B(n_449),
.C(n_483),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_579),
.B(n_585),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_554),
.B(n_514),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_537),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_540),
.A2(n_472),
.B(n_481),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_552),
.A2(n_472),
.B(n_481),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_548),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_529),
.A2(n_500),
.B(n_484),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_532),
.B(n_486),
.Y(n_603)
);

OR2x6_ASAP7_75t_SL g604 ( 
.A(n_575),
.B(n_504),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_574),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_547),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_580),
.B(n_523),
.Y(n_608)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_568),
.A2(n_588),
.B(n_571),
.C(n_539),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_529),
.A2(n_500),
.B(n_484),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_537),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_570),
.B(n_521),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_543),
.A2(n_544),
.B1(n_545),
.B2(n_573),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_531),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_574),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_553),
.A2(n_489),
.B(n_487),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_558),
.B(n_488),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_567),
.A2(n_560),
.B1(n_577),
.B2(n_561),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_555),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_531),
.A2(n_500),
.B(n_484),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_557),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_535),
.B(n_519),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_542),
.B(n_519),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_572),
.B(n_523),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_564),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_555),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_590),
.A2(n_505),
.B(n_503),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_533),
.A2(n_487),
.B(n_463),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_591),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_555),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_566),
.A2(n_487),
.B(n_509),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_541),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_569),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_582),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_582),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_590),
.A2(n_505),
.B(n_496),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_565),
.A2(n_505),
.B(n_496),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_565),
.A2(n_496),
.B(n_518),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_551),
.B(n_523),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_565),
.A2(n_559),
.B(n_556),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_584),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_584),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_587),
.A2(n_496),
.B(n_524),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_567),
.B(n_524),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_586),
.A2(n_495),
.B(n_30),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_577),
.B(n_495),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_586),
.A2(n_495),
.B(n_32),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_581),
.A2(n_583),
.B(n_534),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_534),
.A2(n_495),
.B(n_33),
.Y(n_651)
);

INVxp33_ASAP7_75t_SL g652 ( 
.A(n_541),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_560),
.A2(n_527),
.B1(n_504),
.B2(n_506),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_562),
.A2(n_34),
.B(n_28),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_624),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_596),
.B(n_572),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_606),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_SL g658 ( 
.A1(n_629),
.A2(n_609),
.B(n_616),
.C(n_632),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_614),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_645),
.A2(n_562),
.B(n_592),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_603),
.B(n_558),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_618),
.A2(n_549),
.B1(n_550),
.B2(n_576),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_597),
.B(n_550),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_621),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_594),
.A2(n_536),
.B(n_576),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_607),
.B(n_530),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_613),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_608),
.A2(n_528),
.B(n_530),
.C(n_589),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_637),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_630),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_516),
.Y(n_672)
);

OAI221xp5_ASAP7_75t_L g673 ( 
.A1(n_595),
.A2(n_507),
.B1(n_538),
.B2(n_593),
.C(n_516),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_613),
.B(n_11),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_612),
.B(n_12),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_646),
.B(n_538),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_617),
.B(n_593),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_624),
.B(n_37),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_638),
.A2(n_124),
.B(n_204),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_602),
.A2(n_122),
.B(n_203),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_623),
.B(n_13),
.Y(n_681)
);

BUFx8_ASAP7_75t_SL g682 ( 
.A(n_601),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_636),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_610),
.A2(n_620),
.B(n_600),
.Y(n_684)
);

AO22x1_ASAP7_75t_L g685 ( 
.A1(n_652),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_598),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_618),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_626),
.B(n_16),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_634),
.B(n_17),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_633),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_644),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_R g692 ( 
.A(n_605),
.B(n_38),
.Y(n_692)
);

OAI22x1_ASAP7_75t_L g693 ( 
.A1(n_653),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_635),
.B(n_19),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_625),
.A2(n_39),
.B(n_40),
.C(n_42),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_622),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_648),
.A2(n_48),
.B(n_49),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_641),
.B(n_643),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_604),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_642),
.B(n_50),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_605),
.B(n_52),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_611),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_598),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_SL g704 ( 
.A1(n_611),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_651),
.A2(n_58),
.B(n_60),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_619),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_619),
.B(n_627),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_627),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_631),
.B(n_61),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_640),
.B(n_62),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_671),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_682),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_655),
.Y(n_714)
);

BUFx12f_ASAP7_75t_L g715 ( 
.A(n_655),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_659),
.Y(n_716)
);

BUFx12f_ASAP7_75t_L g717 ( 
.A(n_655),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_683),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_699),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_709),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_663),
.Y(n_721)
);

INVx6_ASAP7_75t_L g722 ( 
.A(n_672),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_709),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_691),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_657),
.Y(n_725)
);

BUFx2_ASAP7_75t_SL g726 ( 
.A(n_703),
.Y(n_726)
);

BUFx4f_ASAP7_75t_SL g727 ( 
.A(n_677),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_656),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_709),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_706),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_698),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_676),
.Y(n_732)
);

BUFx2_ASAP7_75t_SL g733 ( 
.A(n_703),
.Y(n_733)
);

BUFx2_ASAP7_75t_SL g734 ( 
.A(n_702),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_668),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_664),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_686),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_666),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_690),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_686),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_670),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_667),
.B(n_654),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_708),
.B(n_599),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_708),
.Y(n_744)
);

CKINVDCx16_ASAP7_75t_R g745 ( 
.A(n_678),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_692),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_673),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_706),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_694),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_674),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_707),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_661),
.B(n_650),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_711),
.B(n_660),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_710),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_675),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_688),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_681),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_701),
.B(n_639),
.Y(n_758)
);

BUFx2_ASAP7_75t_SL g759 ( 
.A(n_665),
.Y(n_759)
);

INVx3_ASAP7_75t_SL g760 ( 
.A(n_693),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_679),
.B(n_628),
.Y(n_761)
);

BUFx4_ASAP7_75t_SL g762 ( 
.A(n_685),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_689),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_700),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_704),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_687),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_662),
.Y(n_767)
);

NAND2x1p5_ASAP7_75t_L g768 ( 
.A(n_697),
.B(n_647),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_704),
.Y(n_769)
);

INVx3_ASAP7_75t_SL g770 ( 
.A(n_669),
.Y(n_770)
);

BUFx10_ASAP7_75t_L g771 ( 
.A(n_695),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_696),
.Y(n_772)
);

INVx6_ASAP7_75t_L g773 ( 
.A(n_680),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_658),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_684),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_705),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_659),
.Y(n_777)
);

INVx6_ASAP7_75t_SL g778 ( 
.A(n_682),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_752),
.A2(n_649),
.B(n_64),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_728),
.B(n_63),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_751),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_757),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_731),
.B(n_68),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_725),
.Y(n_784)
);

OAI21x1_ASAP7_75t_SL g785 ( 
.A1(n_767),
.A2(n_69),
.B(n_75),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_716),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_721),
.B(n_76),
.Y(n_787)
);

AOI221xp5_ASAP7_75t_L g788 ( 
.A1(n_766),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_714),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_712),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_769),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_753),
.A2(n_87),
.B(n_88),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_739),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_770),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_722),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_761),
.A2(n_96),
.B(n_99),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_755),
.A2(n_100),
.B1(n_102),
.B2(n_107),
.C(n_110),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_765),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_737),
.B(n_114),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_735),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_739),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_735),
.Y(n_802)
);

INVx3_ASAP7_75t_R g803 ( 
.A(n_778),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_718),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_715),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_718),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_768),
.A2(n_115),
.B(n_116),
.Y(n_807)
);

BUFx8_ASAP7_75t_L g808 ( 
.A(n_717),
.Y(n_808)
);

AOI221xp5_ASAP7_75t_L g809 ( 
.A1(n_759),
.A2(n_117),
.B1(n_118),
.B2(n_125),
.C(n_126),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_724),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_760),
.A2(n_127),
.B(n_128),
.C(n_129),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_750),
.B(n_130),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_738),
.Y(n_813)
);

OAI222xp33_ASAP7_75t_L g814 ( 
.A1(n_745),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.C1(n_135),
.C2(n_137),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_741),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_775),
.A2(n_138),
.B(n_139),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_750),
.B(n_140),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_724),
.Y(n_818)
);

BUFx4f_ASAP7_75t_SL g819 ( 
.A(n_778),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_732),
.B(n_141),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_737),
.B(n_142),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_777),
.Y(n_822)
);

NAND2x1p5_ASAP7_75t_L g823 ( 
.A(n_737),
.B(n_143),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_714),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_747),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_714),
.Y(n_826)
);

AO21x2_ASAP7_75t_L g827 ( 
.A1(n_775),
.A2(n_149),
.B(n_152),
.Y(n_827)
);

BUFx10_ASAP7_75t_L g828 ( 
.A(n_746),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_L g829 ( 
.A(n_772),
.B(n_153),
.C(n_154),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_736),
.B(n_763),
.Y(n_830)
);

AO31x2_ASAP7_75t_L g831 ( 
.A1(n_772),
.A2(n_156),
.A3(n_158),
.B(n_159),
.Y(n_831)
);

OAI21x1_ASAP7_75t_SL g832 ( 
.A1(n_756),
.A2(n_161),
.B(n_162),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_729),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_806),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_800),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_830),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_806),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_815),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_786),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_800),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_802),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_SL g842 ( 
.A1(n_829),
.A2(n_745),
.B1(n_771),
.B2(n_774),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_783),
.A2(n_758),
.B(n_742),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_804),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_810),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_819),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_818),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_822),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_784),
.Y(n_849)
);

BUFx2_ASAP7_75t_R g850 ( 
.A(n_805),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_813),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_790),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_793),
.B(n_754),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_796),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_801),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_781),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_833),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_831),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_833),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_831),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_827),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_833),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_807),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_792),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_816),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_812),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_789),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_817),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_789),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_789),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_832),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_787),
.B(n_774),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_785),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_824),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_SL g875 ( 
.A1(n_779),
.A2(n_771),
.B1(n_774),
.B2(n_764),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_811),
.A2(n_763),
.B(n_758),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_799),
.A2(n_730),
.B(n_748),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_795),
.B(n_739),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_R g879 ( 
.A(n_868),
.B(n_820),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_836),
.B(n_749),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_846),
.Y(n_881)
);

NOR2x1p5_ASAP7_75t_L g882 ( 
.A(n_868),
.B(n_713),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_856),
.B(n_855),
.Y(n_883)
);

INVxp33_ASAP7_75t_L g884 ( 
.A(n_878),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_834),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_857),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_R g887 ( 
.A(n_846),
.B(n_808),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_834),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_R g889 ( 
.A(n_872),
.B(n_780),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_837),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_866),
.B(n_754),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_862),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_R g893 ( 
.A(n_843),
.B(n_808),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_856),
.B(n_719),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_872),
.B(n_754),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_837),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_842),
.A2(n_875),
.B1(n_825),
.B2(n_782),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_852),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_853),
.B(n_828),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_873),
.B(n_776),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_850),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_851),
.B(n_849),
.Y(n_902)
);

AND2x4_ASAP7_75t_SL g903 ( 
.A(n_853),
.B(n_859),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_857),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_853),
.B(n_828),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_835),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_874),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_847),
.B(n_826),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_849),
.B(n_824),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_878),
.B(n_722),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_849),
.B(n_743),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_867),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_885),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_906),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_884),
.B(n_840),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_897),
.A2(n_873),
.B1(n_871),
.B2(n_876),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_885),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_883),
.B(n_840),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_903),
.B(n_841),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_888),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_886),
.B(n_841),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_881),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_888),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_890),
.B(n_839),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_890),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_899),
.B(n_803),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_896),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_896),
.Y(n_928)
);

NAND2x1_ASAP7_75t_L g929 ( 
.A(n_900),
.B(n_839),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_900),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_886),
.B(n_845),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_912),
.B(n_907),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_907),
.B(n_845),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_894),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_889),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_929),
.A2(n_858),
.B(n_860),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_914),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_920),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_924),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_935),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_913),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_928),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_932),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_924),
.Y(n_944)
);

OAI22xp33_ASAP7_75t_L g945 ( 
.A1(n_934),
.A2(n_879),
.B1(n_889),
.B2(n_930),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_917),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_929),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_930),
.Y(n_948)
);

OAI21xp33_ASAP7_75t_L g949 ( 
.A1(n_916),
.A2(n_893),
.B(n_911),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_923),
.A2(n_925),
.B(n_927),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_923),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_SL g952 ( 
.A1(n_926),
.A2(n_814),
.B(n_794),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_948),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_945),
.A2(n_882),
.B1(n_904),
.B2(n_898),
.Y(n_954)
);

OA21x2_ASAP7_75t_L g955 ( 
.A1(n_940),
.A2(n_932),
.B(n_922),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_944),
.B(n_891),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_939),
.B(n_908),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_937),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_943),
.B(n_905),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_941),
.Y(n_960)
);

AOI221xp5_ASAP7_75t_L g961 ( 
.A1(n_945),
.A2(n_880),
.B1(n_915),
.B2(n_902),
.C(n_895),
.Y(n_961)
);

INVx5_ASAP7_75t_SL g962 ( 
.A(n_947),
.Y(n_962)
);

OAI221xp5_ASAP7_75t_L g963 ( 
.A1(n_949),
.A2(n_879),
.B1(n_895),
.B2(n_922),
.C(n_901),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_946),
.B(n_915),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_960),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_955),
.B(n_947),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_953),
.B(n_941),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_958),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_959),
.B(n_947),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_957),
.B(n_942),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_962),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_947),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_962),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_965),
.B(n_971),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_967),
.B(n_956),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_965),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_973),
.B(n_961),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_966),
.A2(n_954),
.B1(n_963),
.B2(n_952),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_969),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_968),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_979),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_974),
.B(n_969),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_975),
.B(n_970),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_977),
.B(n_972),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_976),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_978),
.B(n_972),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_980),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_979),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_974),
.B(n_942),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_979),
.B(n_887),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_976),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_983),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_988),
.B(n_938),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_990),
.B(n_887),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_991),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_988),
.B(n_938),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_982),
.B(n_918),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_981),
.B(n_950),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_991),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_986),
.B(n_918),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_992),
.B(n_984),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_994),
.B(n_985),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_993),
.B(n_989),
.Y(n_1003)
);

OAI221xp5_ASAP7_75t_L g1004 ( 
.A1(n_998),
.A2(n_987),
.B1(n_797),
.B2(n_791),
.C(n_809),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_1000),
.B(n_910),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_997),
.B(n_951),
.Y(n_1006)
);

AOI211xp5_ASAP7_75t_L g1007 ( 
.A1(n_996),
.A2(n_798),
.B(n_762),
.C(n_788),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_996),
.B(n_931),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_1002),
.B(n_995),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1001),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1008),
.Y(n_1012)
);

AO22x1_ASAP7_75t_L g1013 ( 
.A1(n_1005),
.A2(n_999),
.B1(n_900),
.B2(n_919),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1011),
.B(n_1006),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1010),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1012),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1009),
.B(n_1004),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1013),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_SL g1019 ( 
.A1(n_1011),
.A2(n_823),
.B(n_821),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_1015),
.A2(n_1007),
.B(n_877),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_1016),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_L g1022 ( 
.A(n_1014),
.B(n_734),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_931),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1018),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1021),
.B(n_1019),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1022),
.A2(n_871),
.B(n_744),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_SL g1027 ( 
.A(n_1024),
.B(n_893),
.C(n_727),
.Y(n_1027)
);

AOI211xp5_ASAP7_75t_L g1028 ( 
.A1(n_1020),
.A2(n_723),
.B(n_729),
.C(n_870),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_1023),
.A2(n_861),
.B(n_877),
.C(n_936),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_L g1030 ( 
.A(n_1025),
.B(n_720),
.C(n_909),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1028),
.B(n_933),
.Y(n_1031)
);

AOI221x1_ASAP7_75t_L g1032 ( 
.A1(n_1027),
.A2(n_1026),
.B1(n_1029),
.B2(n_726),
.C(n_733),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_SL g1033 ( 
.A(n_1025),
.B(n_729),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1027),
.B(n_720),
.Y(n_1034)
);

OAI211xp5_ASAP7_75t_L g1035 ( 
.A1(n_1025),
.A2(n_740),
.B(n_874),
.C(n_730),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_1027),
.A2(n_861),
.B(n_903),
.C(n_869),
.Y(n_1036)
);

OAI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_1027),
.A2(n_892),
.B(n_919),
.Y(n_1037)
);

AOI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_1034),
.A2(n_892),
.B1(n_864),
.B2(n_876),
.C(n_862),
.Y(n_1038)
);

NOR2x1p5_ASAP7_75t_L g1039 ( 
.A(n_1031),
.B(n_748),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1030),
.B(n_892),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_SL g1041 ( 
.A(n_1036),
.B(n_165),
.C(n_167),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1037),
.B(n_921),
.Y(n_1042)
);

OAI221xp5_ASAP7_75t_L g1043 ( 
.A1(n_1033),
.A2(n_773),
.B1(n_864),
.B2(n_854),
.C(n_863),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_740),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1032),
.Y(n_1045)
);

OAI211xp5_ASAP7_75t_L g1046 ( 
.A1(n_1032),
.A2(n_867),
.B(n_862),
.C(n_869),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1042),
.B(n_921),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1045),
.A2(n_900),
.B1(n_892),
.B2(n_919),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_1040),
.B(n_876),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_1046),
.B(n_933),
.Y(n_1050)
);

NAND5xp2_ASAP7_75t_L g1051 ( 
.A(n_1041),
.B(n_843),
.C(n_838),
.D(n_171),
.E(n_172),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_1039),
.B(n_869),
.Y(n_1052)
);

NOR2x1_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_1043),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1038),
.B(n_900),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1045),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1045),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_1039),
.Y(n_1057)
);

NAND2x1_ASAP7_75t_L g1058 ( 
.A(n_1041),
.B(n_862),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_1055),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1056),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_1053),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_SL g1062 ( 
.A(n_1057),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_1052),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_1058),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1051),
.A2(n_865),
.B(n_863),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_1047),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1061),
.B(n_1050),
.Y(n_1067)
);

XOR2xp5_ASAP7_75t_L g1068 ( 
.A(n_1066),
.B(n_1054),
.Y(n_1068)
);

AOI211xp5_ASAP7_75t_SL g1069 ( 
.A1(n_1064),
.A2(n_1049),
.B(n_1048),
.C(n_173),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_1060),
.A2(n_168),
.B(n_169),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1062),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1059),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_SL g1073 ( 
.A1(n_1063),
.A2(n_862),
.B1(n_773),
.B2(n_854),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_1070),
.Y(n_1074)
);

OAI221xp5_ASAP7_75t_L g1075 ( 
.A1(n_1067),
.A2(n_1065),
.B1(n_863),
.B2(n_854),
.C(n_865),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1071),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1074),
.Y(n_1077)
);

XNOR2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1077),
.B(n_1068),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_1076),
.B1(n_1072),
.B2(n_1075),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1079),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_1069),
.B(n_1073),
.C(n_177),
.Y(n_1081)
);

AOI222xp33_ASAP7_75t_SL g1082 ( 
.A1(n_1080),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.C1(n_180),
.C2(n_182),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1081),
.A2(n_743),
.B1(n_844),
.B2(n_848),
.Y(n_1083)
);

AOI221xp5_ASAP7_75t_R g1084 ( 
.A1(n_1082),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.C(n_188),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1085),
.A2(n_192),
.B(n_193),
.Y(n_1086)
);

AOI22x1_ASAP7_75t_L g1087 ( 
.A1(n_1084),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_1087)
);

NAND4xp25_ASAP7_75t_L g1088 ( 
.A(n_1086),
.B(n_1087),
.C(n_198),
.D(n_199),
.Y(n_1088)
);

AOI211xp5_ASAP7_75t_L g1089 ( 
.A1(n_1088),
.A2(n_197),
.B(n_200),
.C(n_202),
.Y(n_1089)
);


endmodule