module fake_jpeg_24744_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_62),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_46),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_57),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_56),
.B1(n_60),
.B2(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx12f_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_16),
.B1(n_27),
.B2(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_17),
.B1(n_26),
.B2(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_65),
.Y(n_95)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_72),
.B1(n_77),
.B2(n_83),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_32),
.B1(n_31),
.B2(n_36),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_78),
.B1(n_82),
.B2(n_45),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_33),
.C(n_37),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_52),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_41),
.B1(n_37),
.B2(n_17),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_53),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_15),
.B1(n_21),
.B2(n_23),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_41),
.B1(n_37),
.B2(n_28),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_50),
.B1(n_62),
.B2(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_97),
.B1(n_104),
.B2(n_81),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_56),
.B1(n_49),
.B2(n_48),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_67),
.B1(n_65),
.B2(n_83),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_98),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_42),
.B(n_57),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_74),
.B(n_75),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_61),
.B1(n_48),
.B2(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_102),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_66),
.B1(n_63),
.B2(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_24),
.B(n_25),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_120),
.B1(n_28),
.B2(n_22),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_67),
.B1(n_74),
.B2(n_44),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_108),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_121),
.Y(n_130)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_84),
.B(n_97),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_83),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_88),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_101),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_148),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_84),
.B1(n_102),
.B2(n_85),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_138),
.B1(n_147),
.B2(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_139),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_127),
.A2(n_104),
.B(n_95),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_123),
.B(n_128),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_137),
.B(n_124),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_103),
.B1(n_90),
.B2(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_106),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_148),
.C(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_109),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_44),
.B1(n_41),
.B2(n_23),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_44),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_149),
.Y(n_155)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_156),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_121),
.B(n_114),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_138),
.Y(n_188)
);

AOI211xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_111),
.B(n_116),
.C(n_118),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_162),
.B1(n_164),
.B2(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_165),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_134),
.A2(n_118),
.B1(n_120),
.B2(n_107),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_114),
.B(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_147),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_117),
.B1(n_112),
.B2(n_126),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_171),
.B1(n_143),
.B2(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_140),
.C(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_117),
.B1(n_112),
.B2(n_109),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_173),
.B1(n_190),
.B2(n_55),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_137),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_180),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_145),
.C(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_129),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_55),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_143),
.Y(n_189)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_162),
.B1(n_157),
.B2(n_151),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_194),
.B1(n_201),
.B2(n_7),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_157),
.B1(n_168),
.B2(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_163),
.B1(n_167),
.B2(n_151),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_160),
.C(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_198),
.C(n_185),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_1),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_55),
.C(n_21),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_15),
.B1(n_28),
.B2(n_3),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_1),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_55),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_190),
.B(n_185),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_211),
.B(n_208),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_186),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_207),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_210),
.C(n_211),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_214),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_182),
.C(n_175),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_184),
.C(n_55),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_28),
.C(n_2),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_7),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_218),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_202),
.B1(n_193),
.B2(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_191),
.B(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_214),
.C(n_8),
.Y(n_230)
);

AOI221xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_192),
.B1(n_8),
.B2(n_9),
.C(n_14),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_229),
.B(n_234),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_235),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_6),
.Y(n_231)
);

OAI21x1_ASAP7_75t_SL g237 ( 
.A1(n_231),
.A2(n_233),
.B(n_11),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_6),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_6),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_9),
.B(n_13),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_231),
.A3(n_229),
.B1(n_224),
.B2(n_10),
.C1(n_5),
.C2(n_13),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_10),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_232),
.A2(n_224),
.B(n_223),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_241),
.B(n_242),
.Y(n_245)
);

NAND2x1_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_238),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_5),
.B1(n_13),
.B2(n_10),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_14),
.B(n_2),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_239),
.B(n_14),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_1),
.B(n_2),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_245),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_251),
.B1(n_248),
.B2(n_3),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_2),
.C(n_3),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_4),
.Y(n_254)
);


endmodule