module fake_netlist_5_1475_n_39 (n_8, n_4, n_5, n_7, n_0, n_2, n_3, n_6, n_1, n_39);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_2;
input n_3;
input n_6;
input n_1;

output n_39;

wire n_29;
wire n_16;
wire n_12;
wire n_9;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_10;
wire n_24;
wire n_28;
wire n_21;
wire n_34;
wire n_38;
wire n_32;
wire n_35;
wire n_11;
wire n_17;
wire n_19;
wire n_37;
wire n_15;
wire n_26;
wire n_30;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_20;

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx5p33_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

AND3x2_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.C(n_2),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx3_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_9),
.C(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

NAND4xp25_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_18),
.C(n_19),
.D(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

AOI221xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_19),
.B1(n_20),
.B2(n_15),
.C(n_16),
.Y(n_27)
);

NOR2x1_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AND3x1_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_20),
.C(n_16),
.Y(n_30)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NAND4xp25_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_28),
.C(n_3),
.D(n_5),
.Y(n_33)
);

AOI322xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_1),
.C2(n_8),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_31),
.Y(n_35)
);

AO22x2_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_31),
.B1(n_7),
.B2(n_8),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_37),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_35),
.B1(n_36),
.B2(n_33),
.Y(n_39)
);


endmodule