module fake_jpeg_21374_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_6),
.B(n_10),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_44),
.B1(n_16),
.B2(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_24),
.C(n_14),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_14),
.B1(n_27),
.B2(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_54),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_33),
.B(n_35),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_30),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_49),
.C(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_22),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_24),
.B1(n_20),
.B2(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_43),
.B1(n_25),
.B2(n_21),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_45),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_56),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_54),
.B1(n_59),
.B2(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_85),
.C(n_15),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_58),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_92),
.B(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_77),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_15),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_57),
.B1(n_21),
.B2(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_75),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_57),
.B(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_93),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_79),
.B(n_73),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_104),
.B(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_102),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_17),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_90),
.C(n_81),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_110),
.C(n_17),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_86),
.Y(n_109)
);

NAND4xp25_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_7),
.C(n_10),
.D(n_11),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_92),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_98),
.A3(n_101),
.B1(n_97),
.B2(n_103),
.C1(n_84),
.C2(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_111),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_107),
.C(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_110),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_12),
.B(n_3),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_122),
.A2(n_118),
.B1(n_107),
.B2(n_112),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_117),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_127),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_1),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_129),
.A2(n_121),
.B1(n_17),
.B2(n_12),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_130),
.B(n_131),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);


endmodule