module fake_aes_5673_n_34 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_6), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_1), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_2), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_7), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_10), .B1(n_13), .B2(n_12), .Y(n_16) );
O2A1O1Ixp5_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_0), .B(n_1), .C(n_2), .Y(n_17) );
O2A1O1Ixp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_0), .B(n_1), .C(n_2), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_20) );
AOI22xp33_ASAP7_75t_SL g21 ( .A1(n_16), .A2(n_10), .B1(n_9), .B2(n_14), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_16), .B(n_15), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AOI211xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_19), .B(n_21), .C(n_18), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
NAND4xp25_ASAP7_75t_L g28 ( .A(n_26), .B(n_25), .C(n_17), .D(n_24), .Y(n_28) );
AND3x2_ASAP7_75t_L g29 ( .A(n_27), .B(n_8), .C(n_26), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_29), .Y(n_30) );
INVx2_ASAP7_75t_SL g31 ( .A(n_28), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_8), .B1(n_27), .B2(n_31), .Y(n_33) );
AOI22xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_34) );
endmodule