module fake_jpeg_17478_n_382 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_40),
.B(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_21),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_46),
.B(n_54),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_29),
.B(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_63),
.Y(n_74)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_29),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_66),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_32),
.B(n_28),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_34),
.B(n_30),
.C(n_23),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_17),
.B1(n_31),
.B2(n_33),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_69),
.A2(n_73),
.B1(n_78),
.B2(n_112),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_70),
.A2(n_81),
.B1(n_87),
.B2(n_92),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_13),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_72),
.B(n_11),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_31),
.B1(n_22),
.B2(n_34),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_31),
.B1(n_23),
.B2(n_34),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_77),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_63),
.B1(n_22),
.B2(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_80),
.B(n_97),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_23),
.B1(n_35),
.B2(n_25),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_30),
.B1(n_36),
.B2(n_35),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_88),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_36),
.B1(n_35),
.B2(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_26),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_36),
.B1(n_35),
.B2(n_25),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_24),
.B1(n_25),
.B2(n_14),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_106),
.B1(n_111),
.B2(n_113),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_16),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_10),
.B(n_0),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_102),
.B(n_105),
.Y(n_154)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_27),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_24),
.B1(n_14),
.B2(n_16),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_45),
.A2(n_24),
.B1(n_16),
.B2(n_14),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_48),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_60),
.A2(n_27),
.B1(n_26),
.B2(n_5),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_61),
.B1(n_6),
.B2(n_9),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_26),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_12),
.B1(n_2),
.B2(n_6),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_125),
.B1(n_153),
.B2(n_89),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_123),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_124),
.B(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_12),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_133),
.A2(n_139),
.B1(n_134),
.B2(n_122),
.Y(n_197)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_61),
.B1(n_52),
.B2(n_44),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_134),
.A2(n_161),
.B1(n_109),
.B2(n_116),
.Y(n_185)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_91),
.B(n_26),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_137),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_74),
.B(n_6),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_44),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_9),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_151),
.Y(n_177)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

BUFx24_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_44),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_150),
.A2(n_163),
.B1(n_164),
.B2(n_125),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_82),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_68),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_75),
.B(n_12),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_159),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_85),
.B(n_109),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_114),
.Y(n_158)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_84),
.A2(n_0),
.B1(n_117),
.B2(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_68),
.A2(n_104),
.B1(n_103),
.B2(n_89),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_0),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_82),
.B(n_0),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_166),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_95),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_204),
.B1(n_147),
.B2(n_160),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_191),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_SL g237 ( 
.A(n_182),
.B(n_194),
.C(n_177),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_193),
.B1(n_197),
.B2(n_198),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_116),
.B(n_95),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_90),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_90),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_195),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_127),
.A2(n_98),
.B1(n_128),
.B2(n_143),
.Y(n_193)
);

AO21x2_ASAP7_75t_L g194 ( 
.A1(n_134),
.A2(n_98),
.B(n_150),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_202),
.B1(n_208),
.B2(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_126),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_148),
.C(n_143),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_207),
.C(n_186),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_133),
.A2(n_129),
.B1(n_152),
.B2(n_159),
.Y(n_202)
);

OAI22x1_ASAP7_75t_L g203 ( 
.A1(n_122),
.A2(n_131),
.B1(n_158),
.B2(n_141),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_188),
.B1(n_210),
.B2(n_181),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_131),
.A2(n_168),
.B1(n_167),
.B2(n_135),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_149),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_132),
.A2(n_155),
.B1(n_162),
.B2(n_158),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_160),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_120),
.B(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_191),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_120),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_206),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_160),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_219),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_222),
.B1(n_223),
.B2(n_230),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_147),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_228),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_193),
.B1(n_198),
.B2(n_176),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_224),
.B(n_234),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_227),
.B(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_229),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_170),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_185),
.B1(n_202),
.B2(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_179),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_247),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_170),
.C(n_174),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_246),
.C(n_224),
.Y(n_270)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_235),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_238),
.B1(n_242),
.B2(n_249),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_205),
.B1(n_211),
.B2(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_240),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_171),
.B(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_189),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_206),
.B1(n_178),
.B2(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_178),
.B(n_200),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_245),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_188),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_244),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_175),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_175),
.B(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_190),
.B(n_213),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_199),
.A2(n_194),
.B1(n_172),
.B2(n_197),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_201),
.A2(n_194),
.B1(n_172),
.B2(n_197),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_252),
.B1(n_215),
.B2(n_227),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_187),
.A2(n_194),
.B1(n_193),
.B2(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_177),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_254),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_220),
.A2(n_236),
.B1(n_225),
.B2(n_252),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_266),
.B1(n_275),
.B2(n_269),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_226),
.B(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_282),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_216),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_273),
.B(n_277),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_225),
.A2(n_230),
.B(n_249),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_285),
.B1(n_273),
.B2(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_227),
.A2(n_221),
.B(n_223),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_221),
.A2(n_251),
.B(n_238),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_232),
.B(n_229),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_218),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_233),
.A2(n_217),
.B(n_250),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_286),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_219),
.A2(n_234),
.B(n_225),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_216),
.A2(n_186),
.B(n_234),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_291),
.A2(n_294),
.B1(n_309),
.B2(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_261),
.B1(n_269),
.B2(n_266),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_284),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_295),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_257),
.B(n_272),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_260),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_297),
.A2(n_303),
.B(n_308),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_299),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_276),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_300),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_260),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_264),
.C(n_270),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_259),
.Y(n_305)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_255),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_274),
.A2(n_261),
.B1(n_258),
.B2(n_271),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_261),
.A2(n_278),
.B1(n_277),
.B2(n_280),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_262),
.B(n_257),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_263),
.C(n_283),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_261),
.A2(n_285),
.B1(n_286),
.B2(n_256),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_256),
.Y(n_316)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_316),
.A2(n_301),
.B1(n_290),
.B2(n_288),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

NOR3xp33_ASAP7_75t_SL g319 ( 
.A(n_294),
.B(n_264),
.C(n_255),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_320),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_298),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_289),
.C(n_307),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_307),
.C(n_306),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_314),
.C(n_312),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_332),
.C(n_301),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_311),
.C(n_292),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_327),
.Y(n_334)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_296),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_336),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_309),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_339),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_310),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_343),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_333),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_349),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_310),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_333),
.A2(n_288),
.B(n_290),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_345),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_308),
.B(n_303),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_347),
.A2(n_348),
.B(n_324),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_297),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_299),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_348),
.Y(n_356)
);

AOI221xp5_ASAP7_75t_L g359 ( 
.A1(n_337),
.A2(n_342),
.B1(n_347),
.B2(n_323),
.C(n_345),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_359),
.B(n_361),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_346),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_340),
.C(n_343),
.Y(n_364)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_349),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_365),
.A2(n_367),
.B(n_355),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_351),
.A2(n_322),
.B1(n_329),
.B2(n_325),
.Y(n_366)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_366),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_339),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_367),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_363),
.A2(n_356),
.B1(n_322),
.B2(n_361),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_370),
.A2(n_353),
.B1(n_354),
.B2(n_360),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_350),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_373),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_357),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_369),
.C(n_376),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_374),
.C(n_362),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_364),
.C(n_358),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_328),
.C(n_327),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_352),
.Y(n_382)
);


endmodule