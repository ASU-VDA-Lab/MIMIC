module fake_jpeg_20472_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_40),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_22),
.B1(n_18),
.B2(n_25),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_33),
.B1(n_34),
.B2(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_73),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_65),
.B(n_69),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_39),
.B1(n_37),
.B2(n_21),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_33),
.B1(n_34),
.B2(n_23),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_70),
.B1(n_75),
.B2(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_15),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_23),
.B1(n_15),
.B2(n_31),
.Y(n_70)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_23),
.B1(n_31),
.B2(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_48),
.B1(n_27),
.B2(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_84),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_27),
.Y(n_106)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_92),
.B(n_95),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_101),
.B1(n_102),
.B2(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_65),
.B(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_108),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_27),
.B1(n_20),
.B2(n_36),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_67),
.B1(n_70),
.B2(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_76),
.B1(n_82),
.B2(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_19),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_114),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_57),
.A2(n_27),
.B1(n_20),
.B2(n_9),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_19),
.B1(n_16),
.B2(n_27),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_115),
.B(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_120),
.Y(n_144)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_122),
.Y(n_146)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_131),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_82),
.B(n_72),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_133),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_128),
.Y(n_148)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_89),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_134),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_71),
.B(n_57),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_13),
.B(n_14),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_71),
.B(n_79),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_93),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_61),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_60),
.A3(n_107),
.B1(n_98),
.B2(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_164),
.B(n_158),
.Y(n_187)
);

AO21x2_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_101),
.B(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_109),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_169),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_138),
.B1(n_141),
.B2(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_170),
.B1(n_173),
.B2(n_86),
.Y(n_190)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_106),
.C(n_110),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_87),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_87),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_86),
.B1(n_72),
.B2(n_58),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_98),
.C(n_60),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_64),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_138),
.B1(n_129),
.B2(n_125),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_163),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_64),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_56),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_86),
.B1(n_104),
.B2(n_59),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_197),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_125),
.B1(n_118),
.B2(n_135),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_177),
.A2(n_192),
.B1(n_201),
.B2(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_128),
.Y(n_186)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_190),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_130),
.B(n_120),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_196),
.B(n_206),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_104),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_104),
.B1(n_97),
.B2(n_59),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_97),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_195),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_56),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_9),
.B(n_14),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_146),
.B(n_9),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_203),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_149),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_97),
.B1(n_19),
.B2(n_16),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_14),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_12),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_16),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_143),
.A2(n_0),
.B(n_1),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_211),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_167),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_215),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_172),
.CI(n_168),
.CON(n_211),
.SN(n_211)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_198),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_223),
.C(n_206),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_157),
.C(n_145),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_188),
.C(n_182),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_159),
.C(n_147),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_202),
.C(n_205),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_190),
.B1(n_178),
.B2(n_195),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_196),
.A2(n_149),
.B1(n_147),
.B2(n_156),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_149),
.C(n_11),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_201),
.C(n_203),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_200),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_232),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_180),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_235),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_214),
.A2(n_181),
.B1(n_202),
.B2(n_178),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_195),
.B1(n_182),
.B2(n_184),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_239),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_149),
.B1(n_187),
.B2(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_227),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_244),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_226),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_212),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_189),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_233),
.C(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_218),
.B1(n_212),
.B2(n_228),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_251),
.B1(n_234),
.B2(n_240),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_228),
.B1(n_215),
.B2(n_213),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_208),
.B(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_256),
.C(n_243),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_229),
.C(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_11),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_211),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_258),
.A2(n_232),
.B1(n_231),
.B2(n_227),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_271),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_278),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_239),
.B1(n_243),
.B2(n_224),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_251),
.B1(n_261),
.B2(n_6),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_224),
.B1(n_179),
.B2(n_11),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_277),
.B1(n_249),
.B2(n_262),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_255),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_179),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_274),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_10),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_10),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_5),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_0),
.B(n_1),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_1),
.B(n_2),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_273),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_254),
.C(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_287),
.C(n_278),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_289),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_4),
.C(n_5),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_266),
.A2(n_4),
.B(n_5),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_7),
.B(n_8),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_291),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_273),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_279),
.A2(n_280),
.B(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_295),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_276),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_296),
.B(n_297),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_5),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_303),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_296),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_302),
.A3(n_306),
.B1(n_295),
.B2(n_294),
.C1(n_300),
.C2(n_282),
.Y(n_308)
);

XNOR2x2_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_282),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_309),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_310),
.B(n_7),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_7),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_7),
.Y(n_313)
);


endmodule