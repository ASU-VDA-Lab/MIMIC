module real_jpeg_14038_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_33;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_53;
wire n_18;
wire n_22;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_27;
wire n_19;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_3),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_13),
.C(n_23),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_16),
.B1(n_32),
.B2(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_3),
.B(n_49),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_41),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_29),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_26),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_20),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_11),
.B1(n_46),
.B2(n_53),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_17),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_18),
.Y(n_19)
);

AO22x1_ASAP7_75t_SL g22 ( 
.A1(n_13),
.A2(n_14),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

INVx5_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_35),
.B(n_38),
.Y(n_34)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_24),
.B1(n_32),
.B2(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

OA22x2_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_37),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_54),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);


endmodule