module fake_jpeg_25898_n_59 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

INVx11_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_10),
.B1(n_23),
.B2(n_20),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_30),
.B1(n_32),
.B2(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_43),
.B1(n_1),
.B2(n_4),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_5),
.B(n_6),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_51)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_47),
.C(n_9),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_53),
.B(n_51),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_45),
.C(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_8),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_15),
.B(n_16),
.Y(n_57)
);

OAI21x1_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_17),
.B(n_18),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);


endmodule