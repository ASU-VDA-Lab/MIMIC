module fake_aes_1706_n_672 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_672);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_672;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_30), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_43), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_64), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_69), .Y(n_79) );
INVx2_ASAP7_75t_SL g80 ( .A(n_47), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_12), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_22), .Y(n_82) );
BUFx2_ASAP7_75t_L g83 ( .A(n_56), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_36), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_20), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_27), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_74), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_37), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_23), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_72), .Y(n_94) );
INVx3_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
BUFx2_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_33), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_26), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_49), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_54), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_48), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_14), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_17), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_59), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_44), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_11), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_39), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_38), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_29), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_0), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_66), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_32), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_99), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_83), .B(n_1), .Y(n_125) );
INVx2_ASAP7_75t_SL g126 ( .A(n_83), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_96), .B(n_1), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_95), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_76), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_99), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_99), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_96), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_115), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_115), .B(n_4), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_100), .B(n_4), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_117), .B(n_5), .Y(n_141) );
NOR3xp33_ASAP7_75t_L g142 ( .A(n_81), .B(n_5), .C(n_6), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_79), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_78), .B(n_6), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_80), .B(n_115), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_82), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_87), .B(n_7), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_122), .B(n_8), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_113), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_88), .A2(n_42), .B(n_71), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_90), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_90), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_91), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
NAND2x1p5_ASAP7_75t_L g164 ( .A(n_138), .B(n_121), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
BUFx4f_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_135), .B(n_87), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_127), .B(n_103), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_125), .B(n_105), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_127), .B(n_103), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_154), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_154), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_126), .B(n_107), .Y(n_174) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_125), .B(n_121), .Y(n_175) );
OR2x6_ASAP7_75t_L g176 ( .A(n_125), .B(n_120), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_123), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_126), .A2(n_120), .B1(n_85), .B2(n_118), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_125), .B(n_109), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_159), .B(n_85), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_123), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_139), .Y(n_190) );
BUFx10_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
BUFx10_ASAP7_75t_L g192 ( .A(n_124), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_145), .A2(n_108), .B1(n_118), .B2(n_114), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_130), .B(n_119), .Y(n_196) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_130), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_147), .B(n_105), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_141), .A2(n_114), .B1(n_106), .B2(n_116), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_128), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_131), .B(n_119), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_146), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_129), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_123), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_129), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_131), .B(n_106), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_140), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_123), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_160), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_132), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_123), .Y(n_215) );
AO22x2_ASAP7_75t_L g216 ( .A1(n_142), .A2(n_112), .B1(n_111), .B2(n_110), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_132), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_136), .B(n_112), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_136), .B(n_109), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_143), .B(n_111), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_123), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_143), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_198), .B(n_141), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_198), .B(n_144), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_191), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_191), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_177), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_175), .A2(n_144), .B1(n_162), .B2(n_161), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_194), .A2(n_161), .B(n_148), .C(n_149), .Y(n_231) );
INVx4_ASAP7_75t_L g232 ( .A(n_192), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_177), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_192), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_198), .B(n_148), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_167), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_175), .B(n_149), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_172), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_167), .A2(n_162), .B(n_152), .C(n_153), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_196), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_196), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_195), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_174), .B(n_152), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_208), .Y(n_246) );
OAI22xp5_ASAP7_75t_SL g247 ( .A1(n_190), .A2(n_86), .B1(n_104), .B2(n_158), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_212), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_172), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_176), .A2(n_153), .B1(n_93), .B2(n_89), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_179), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_212), .Y(n_252) );
INVxp33_ASAP7_75t_SL g253 ( .A(n_199), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_183), .Y(n_254) );
OR2x2_ASAP7_75t_SL g255 ( .A(n_185), .B(n_158), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_173), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_173), .B(n_168), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_176), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_169), .B(n_150), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_176), .B(n_150), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_167), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_169), .B(n_155), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_171), .B(n_207), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_183), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_189), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_168), .B(n_155), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_164), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_164), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_176), .B(n_156), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_219), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_164), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_170), .B(n_156), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
NOR2xp67_ASAP7_75t_L g276 ( .A(n_180), .B(n_157), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_197), .B(n_102), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_171), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_219), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_207), .Y(n_280) );
INVxp67_ASAP7_75t_L g281 ( .A(n_201), .Y(n_281) );
CKINVDCx6p67_ASAP7_75t_R g282 ( .A(n_170), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_189), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_200), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_226), .B(n_170), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_270), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_228), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_256), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_226), .B(n_207), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_280), .Y(n_291) );
BUFx4f_ASAP7_75t_L g292 ( .A(n_282), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_270), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_259), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_281), .B(n_197), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_270), .Y(n_296) );
BUFx8_ASAP7_75t_L g297 ( .A(n_270), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_230), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_223), .B(n_197), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_273), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_233), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_226), .B(n_181), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_232), .B(n_181), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_273), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_253), .A2(n_216), .B1(n_165), .B2(n_166), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_229), .A2(n_188), .B1(n_187), .B2(n_184), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_253), .B(n_182), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_230), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_232), .B(n_214), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_233), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_230), .Y(n_313) );
CKINVDCx6p67_ASAP7_75t_R g314 ( .A(n_271), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_245), .B(n_217), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_257), .Y(n_317) );
OR2x6_ASAP7_75t_L g318 ( .A(n_271), .B(n_216), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_237), .B(n_282), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_273), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_273), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_237), .A2(n_216), .B1(n_222), .B2(n_218), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_249), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_230), .Y(n_324) );
HAxp5_ASAP7_75t_L g325 ( .A(n_249), .B(n_216), .CON(n_325), .SN(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_271), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_238), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_260), .A2(n_218), .B1(n_213), .B2(n_211), .Y(n_328) );
BUFx12f_ASAP7_75t_L g329 ( .A(n_271), .Y(n_329) );
AOI21x1_ASAP7_75t_L g330 ( .A1(n_277), .A2(n_220), .B(n_202), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_261), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_245), .B(n_204), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_294), .B(n_240), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_290), .B(n_268), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_309), .A2(n_278), .B1(n_258), .B2(n_260), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_329), .A2(n_247), .B1(n_268), .B2(n_263), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_303), .B(n_241), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_285), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_318), .A2(n_260), .B1(n_242), .B2(n_236), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_285), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_288), .A2(n_239), .B(n_276), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_318), .A2(n_239), .B1(n_235), .B2(n_224), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_318), .A2(n_236), .B1(n_261), .B2(n_274), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_318), .A2(n_236), .B1(n_261), .B2(n_274), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_329), .A2(n_267), .B1(n_254), .B2(n_265), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_290), .B(n_225), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_290), .B(n_225), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_307), .A2(n_250), .B1(n_279), .B2(n_275), .Y(n_350) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_297), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_297), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_301), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_315), .A2(n_255), .B1(n_272), .B2(n_264), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_298), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_317), .B(n_243), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_301), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_327), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_298), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_312), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_312), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_298), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_308), .A2(n_231), .B1(n_157), .B2(n_209), .C(n_203), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_333), .B(n_289), .Y(n_364) );
INVx4_ASAP7_75t_L g365 ( .A(n_351), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_336), .A2(n_327), .B1(n_323), .B2(n_302), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_358), .B(n_295), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_304), .B1(n_302), .B2(n_322), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_351), .A2(n_314), .B1(n_292), .B2(n_326), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_351), .A2(n_302), .B1(n_304), .B2(n_314), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_335), .A2(n_299), .B1(n_292), .B2(n_328), .C(n_332), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_356), .Y(n_372) );
AO31x2_ASAP7_75t_L g373 ( .A1(n_354), .A2(n_291), .A3(n_102), .B(n_101), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_339), .A2(n_326), .B1(n_292), .B2(n_304), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_346), .A2(n_277), .B(n_311), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_333), .B(n_319), .Y(n_376) );
OAI211xp5_ASAP7_75t_L g377 ( .A1(n_346), .A2(n_316), .B(n_325), .C(n_319), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_352), .A2(n_306), .B1(n_325), .B2(n_286), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_352), .A2(n_311), .B1(n_306), .B2(n_286), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_363), .B(n_331), .C(n_99), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_311), .B1(n_286), .B2(n_261), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_310), .B1(n_313), .B2(n_298), .Y(n_382) );
CKINVDCx6p67_ASAP7_75t_R g383 ( .A(n_333), .Y(n_383) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_349), .A2(n_110), .B(n_92), .C(n_97), .Y(n_384) );
AO31x2_ASAP7_75t_L g385 ( .A1(n_354), .A2(n_91), .A3(n_92), .B(n_97), .Y(n_385) );
AO31x2_ASAP7_75t_L g386 ( .A1(n_342), .A2(n_98), .A3(n_101), .B(n_193), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_342), .A2(n_284), .B1(n_331), .B2(n_269), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_356), .A2(n_284), .B1(n_331), .B2(n_269), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_337), .A2(n_300), .B1(n_293), .B2(n_305), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_337), .A2(n_234), .B1(n_227), .B2(n_293), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_372), .B(n_337), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_383), .B(n_338), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_378), .A2(n_356), .B1(n_334), .B2(n_347), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_364), .Y(n_394) );
OAI33xp33_ASAP7_75t_L g395 ( .A1(n_384), .A2(n_98), .A3(n_338), .B1(n_348), .B2(n_357), .B3(n_361), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_386), .Y(n_396) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_387), .A2(n_341), .B(n_330), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_377), .B(n_350), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_386), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_350), .B1(n_363), .B2(n_343), .C(n_345), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_370), .A2(n_344), .B1(n_361), .B2(n_360), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_365), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_376), .B(n_340), .Y(n_403) );
OA21x2_ASAP7_75t_L g404 ( .A1(n_380), .A2(n_341), .B(n_361), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_385), .B(n_340), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_374), .A2(n_347), .B1(n_334), .B2(n_360), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_373), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_334), .B1(n_347), .B2(n_340), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_385), .B(n_344), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_373), .B(n_344), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_389), .Y(n_413) );
OAI31xp33_ASAP7_75t_L g414 ( .A1(n_369), .A2(n_347), .A3(n_334), .B(n_353), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_371), .A2(n_334), .B1(n_347), .B2(n_357), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_375), .B(n_360), .C(n_357), .Y(n_416) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_390), .A2(n_353), .B(n_300), .C(n_320), .Y(n_417) );
NAND2x1p5_ASAP7_75t_SL g418 ( .A(n_382), .B(n_355), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
AOI222xp33_ASAP7_75t_SL g420 ( .A1(n_367), .A2(n_9), .B1(n_10), .B2(n_11), .C1(n_12), .C2(n_13), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_379), .B(n_353), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_381), .B(n_287), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_393), .A2(n_355), .B1(n_362), .B2(n_359), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
BUFx2_ASAP7_75t_SL g427 ( .A(n_392), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_406), .B(n_410), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_391), .B(n_200), .Y(n_429) );
INVx2_ASAP7_75t_SL g430 ( .A(n_394), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_394), .B(n_403), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_392), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_400), .A2(n_284), .B1(n_200), .B2(n_206), .C(n_287), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_400), .A2(n_287), .B1(n_320), .B2(n_305), .Y(n_436) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_398), .A2(n_362), .B1(n_359), .B2(n_355), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_403), .B(n_206), .Y(n_438) );
OAI31xp33_ASAP7_75t_L g439 ( .A1(n_414), .A2(n_206), .A3(n_296), .B(n_362), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_414), .B(n_362), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_398), .B(n_359), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_422), .B(n_359), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_419), .B(n_10), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
INVx5_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_408), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_407), .A2(n_296), .B1(n_321), .B2(n_324), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_421), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_408), .Y(n_451) );
AOI21xp5_ASAP7_75t_SL g452 ( .A1(n_417), .A2(n_313), .B(n_310), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_421), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_399), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_399), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_415), .A2(n_409), .B1(n_413), .B2(n_422), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_396), .B(n_15), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_413), .B(n_193), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_396), .B(n_99), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_405), .B(n_158), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_405), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
OAI21xp33_ASAP7_75t_SL g464 ( .A1(n_411), .A2(n_202), .B(n_269), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_411), .B(n_158), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_411), .B(n_15), .Y(n_466) );
OAI322xp33_ASAP7_75t_L g467 ( .A1(n_420), .A2(n_133), .A3(n_134), .B1(n_163), .B2(n_215), .C1(n_251), .C2(n_283), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_399), .B(n_313), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_424), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_401), .A2(n_310), .B(n_313), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_423), .B(n_283), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_424), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_426), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_435), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_446), .B(n_416), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_431), .B(n_418), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_432), .B(n_416), .Y(n_479) );
OR2x6_ASAP7_75t_L g480 ( .A(n_427), .B(n_418), .Y(n_480) );
NOR3xp33_ASAP7_75t_SL g481 ( .A(n_467), .B(n_456), .C(n_429), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_447), .B(n_418), .Y(n_482) );
XOR2x2_ASAP7_75t_L g483 ( .A(n_432), .B(n_420), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_457), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_428), .B(n_397), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_455), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_457), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_428), .B(n_397), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_459), .A2(n_133), .B(n_134), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_441), .B(n_397), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_450), .B(n_397), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_427), .B(n_404), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_433), .B(n_395), .C(n_246), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_455), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_430), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_450), .B(n_404), .Y(n_496) );
AOI32xp33_ASAP7_75t_L g497 ( .A1(n_430), .A2(n_395), .A3(n_246), .B1(n_244), .B2(n_251), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_445), .B(n_404), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_434), .B(n_404), .Y(n_499) );
AOI21x1_ASAP7_75t_L g500 ( .A1(n_459), .A2(n_266), .B(n_244), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_445), .Y(n_501) );
NAND4xp25_ASAP7_75t_SL g502 ( .A(n_439), .B(n_16), .C(n_18), .D(n_19), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_453), .B(n_163), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_462), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_444), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_448), .B(n_163), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_451), .B(n_163), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_459), .B(n_454), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_461), .B(n_163), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_454), .B(n_163), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_134), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_463), .B(n_134), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_469), .B(n_134), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_473), .B(n_134), .Y(n_514) );
AND2x2_ASAP7_75t_SL g515 ( .A(n_466), .B(n_310), .Y(n_515) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_472), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_447), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_466), .B(n_133), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_473), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_468), .B(n_442), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_460), .Y(n_521) );
AND4x1_ASAP7_75t_L g522 ( .A(n_447), .B(n_21), .C(n_24), .D(n_25), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_447), .B(n_133), .C(n_178), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_468), .B(n_133), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_447), .B(n_133), .Y(n_525) );
AOI31xp67_ASAP7_75t_SL g526 ( .A1(n_438), .A2(n_28), .A3(n_31), .B(n_34), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_443), .B(n_266), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_468), .B(n_40), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_458), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_471), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_508), .B(n_440), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_504), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_517), .B(n_464), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_495), .B(n_440), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_520), .B(n_437), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_475), .B(n_449), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_516), .B(n_460), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_505), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_508), .B(n_470), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_477), .B(n_425), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_530), .B(n_436), .Y(n_543) );
NAND2xp33_ASAP7_75t_SL g544 ( .A(n_482), .B(n_452), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_520), .B(n_465), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_494), .Y(n_546) );
OAI31xp67_ASAP7_75t_L g547 ( .A1(n_483), .A2(n_215), .A3(n_452), .B(n_51), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_480), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_494), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_474), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_484), .Y(n_551) );
NOR2xp33_ASAP7_75t_R g552 ( .A(n_502), .B(n_45), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_487), .B(n_465), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_485), .B(n_46), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_485), .B(n_52), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_509), .Y(n_556) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_482), .B(n_246), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_501), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_529), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_488), .B(n_53), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_512), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_480), .B(n_55), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_519), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_478), .B(n_57), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_521), .B(n_58), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_515), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_488), .B(n_61), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_479), .B(n_63), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_521), .B(n_65), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_483), .B(n_67), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_490), .B(n_68), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_519), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_490), .B(n_499), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_480), .B(n_70), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_506), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_506), .Y(n_577) );
NAND2x1_ASAP7_75t_L g578 ( .A(n_480), .B(n_210), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_476), .B(n_75), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_503), .B(n_252), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_493), .A2(n_248), .B1(n_252), .B2(n_205), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_551), .B(n_476), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_571), .B(n_498), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_532), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_558), .B(n_476), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_540), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_561), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_561), .Y(n_588) );
AOI322xp5_ASAP7_75t_L g589 ( .A1(n_574), .A2(n_481), .A3(n_491), .B1(n_496), .B2(n_515), .C1(n_492), .C2(n_489), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_550), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_545), .B(n_491), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_559), .B(n_503), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_534), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_536), .B(n_522), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_534), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_556), .B(n_496), .Y(n_596) );
NOR2x1_ASAP7_75t_SL g597 ( .A(n_533), .B(n_500), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_556), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_567), .B(n_507), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_544), .B(n_528), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_553), .B(n_507), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_537), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_562), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_546), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_546), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_542), .B(n_513), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_542), .Y(n_608) );
OAI32xp33_ASAP7_75t_L g609 ( .A1(n_544), .A2(n_525), .A3(n_526), .B1(n_523), .B2(n_518), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_576), .B(n_577), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_549), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_563), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_531), .B(n_511), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_539), .B(n_514), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_538), .B(n_524), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g617 ( .A1(n_547), .A2(n_497), .B(n_528), .Y(n_617) );
OAI321xp33_ASAP7_75t_L g618 ( .A1(n_535), .A2(n_524), .A3(n_511), .B1(n_513), .B2(n_527), .C(n_526), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_578), .B(n_528), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_581), .A2(n_510), .B1(n_514), .B2(n_248), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_531), .B(n_514), .Y(n_621) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_538), .B(n_510), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g623 ( .A(n_552), .B(n_510), .C(n_186), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_562), .B(n_178), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_563), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g626 ( .A(n_581), .B(n_178), .C(n_186), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_543), .A2(n_178), .B1(n_186), .B2(n_205), .C(n_210), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_569), .B(n_186), .C(n_205), .Y(n_628) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_575), .B(n_221), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_569), .A2(n_205), .B1(n_210), .B2(n_221), .C(n_566), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_533), .A2(n_210), .B(n_221), .Y(n_631) );
AOI211xp5_ASAP7_75t_SL g632 ( .A1(n_548), .A2(n_221), .B(n_575), .C(n_568), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_557), .B(n_579), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g634 ( .A1(n_552), .A2(n_554), .B(n_555), .C(n_579), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_573), .B(n_541), .Y(n_635) );
NOR3x1_ASAP7_75t_L g636 ( .A(n_564), .B(n_560), .C(n_572), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_573), .B(n_541), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_548), .B(n_580), .Y(n_638) );
AO21x1_ASAP7_75t_L g639 ( .A1(n_634), .A2(n_601), .B(n_617), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_634), .A2(n_601), .B1(n_604), .B2(n_594), .Y(n_640) );
OAI211xp5_ASAP7_75t_SL g641 ( .A1(n_589), .A2(n_608), .B(n_632), .C(n_598), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_583), .A2(n_616), .B1(n_622), .B2(n_623), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_587), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_587), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_609), .A2(n_618), .B(n_597), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_590), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_584), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_586), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_619), .A2(n_616), .B(n_629), .C(n_633), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_588), .A2(n_583), .B1(n_635), .B2(n_607), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_638), .A2(n_614), .B1(n_637), .B2(n_596), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_646), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_SL g653 ( .A1(n_640), .A2(n_630), .B(n_631), .C(n_615), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_639), .B(n_582), .Y(n_654) );
NAND2x1_ASAP7_75t_L g655 ( .A(n_643), .B(n_591), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_645), .A2(n_628), .B(n_626), .C(n_592), .Y(n_656) );
AOI221x1_ASAP7_75t_L g657 ( .A1(n_640), .A2(n_626), .B1(n_585), .B2(n_620), .C(n_611), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_647), .Y(n_658) );
AOI322xp5_ASAP7_75t_L g659 ( .A1(n_642), .A2(n_591), .A3(n_614), .B1(n_602), .B2(n_621), .C1(n_599), .C2(n_606), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_654), .A2(n_641), .B1(n_650), .B2(n_649), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_659), .B(n_648), .Y(n_661) );
AND4x1_ASAP7_75t_L g662 ( .A(n_657), .B(n_636), .C(n_624), .D(n_651), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_656), .A2(n_644), .B1(n_615), .B2(n_610), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_661), .A2(n_653), .B1(n_658), .B2(n_652), .C(n_655), .Y(n_664) );
AND3x2_ASAP7_75t_L g665 ( .A(n_662), .B(n_603), .C(n_625), .Y(n_665) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_660), .B(n_627), .C(n_570), .D(n_565), .Y(n_666) );
INVx4_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
NAND3x1_ASAP7_75t_L g668 ( .A(n_664), .B(n_663), .C(n_600), .Y(n_668) );
XNOR2xp5_ASAP7_75t_L g669 ( .A(n_668), .B(n_666), .Y(n_669) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_669), .A2(n_667), .B(n_605), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_612), .B1(n_613), .B2(n_593), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_593), .B(n_595), .Y(n_672) );
endmodule