module fake_jpeg_26703_n_94 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_33),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_16),
.B(n_23),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_27),
.B(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_23),
.B1(n_20),
.B2(n_24),
.Y(n_39)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_9),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_57),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_35),
.C(n_27),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_41),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_35),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_67),
.C(n_12),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_18),
.B1(n_12),
.B2(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_53),
.B1(n_55),
.B2(n_50),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_15),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_69),
.B1(n_8),
.B2(n_6),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_74),
.C(n_65),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_52),
.C(n_11),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_78),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_60),
.B1(n_67),
.B2(n_16),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_77),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_11),
.C(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_80),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_70),
.B(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_1),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_80),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_86),
.C(n_87),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_11),
.C(n_3),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_83),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_92),
.B(n_5),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_87),
.C(n_4),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_5),
.Y(n_94)
);


endmodule