module fake_jpeg_27499_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx11_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx9p33_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_23),
.B1(n_29),
.B2(n_17),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_53),
.B1(n_56),
.B2(n_35),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_23),
.B1(n_17),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_50),
.B1(n_57),
.B2(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_36),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_21),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_25),
.B1(n_21),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_21),
.B1(n_30),
.B2(n_28),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_24),
.B1(n_16),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_69),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_40),
.B(n_41),
.C(n_38),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_82),
.B(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_64),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_36),
.B1(n_35),
.B2(n_38),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_65),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_40),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_72),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_34),
.B1(n_38),
.B2(n_37),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_76),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_36),
.B1(n_21),
.B2(n_16),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_86),
.B1(n_47),
.B2(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_53),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_33),
.Y(n_80)
);

NOR2x1_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_43),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_85),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_30),
.B(n_27),
.C(n_18),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_36),
.C(n_27),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_88),
.C(n_45),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_35),
.B1(n_18),
.B2(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_43),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_35),
.B1(n_32),
.B2(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_43),
.B(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_48),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_32),
.C(n_35),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_102),
.B1(n_66),
.B2(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_93),
.B(n_101),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_75),
.B(n_77),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_45),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_74),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_67),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_112),
.Y(n_120)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_47),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_116),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_69),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_71),
.B1(n_77),
.B2(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_126),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_72),
.C(n_83),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_60),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_64),
.B(n_82),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_80),
.B(n_73),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_127),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_81),
.B1(n_67),
.B2(n_47),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_85),
.A3(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_112),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_58),
.B1(n_66),
.B2(n_4),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_89),
.B1(n_108),
.B2(n_100),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_135),
.B1(n_113),
.B2(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_7),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_102),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_142),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_97),
.B1(n_107),
.B2(n_104),
.C(n_110),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_9),
.Y(n_175)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_100),
.B1(n_109),
.B2(n_91),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_156),
.A2(n_158),
.B1(n_131),
.B2(n_118),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_103),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_103),
.B1(n_11),
.B2(n_12),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_160),
.B(n_9),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_177),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_127),
.C(n_119),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_167),
.C(n_151),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_123),
.B(n_115),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_155),
.B(n_147),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_123),
.C(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_140),
.A2(n_117),
.B1(n_124),
.B2(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_144),
.B1(n_158),
.B2(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_174),
.B1(n_159),
.B2(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_176),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_117),
.B1(n_136),
.B2(n_12),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_188),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_183),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_156),
.B1(n_152),
.B2(n_142),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_184),
.B(n_186),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_192),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_147),
.C(n_143),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_178),
.C(n_166),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_198),
.C(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_172),
.C(n_173),
.Y(n_198)
);

OAI31xp33_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_177),
.A3(n_168),
.B(n_161),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_171),
.B1(n_197),
.B2(n_193),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_170),
.C(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_11),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_188),
.B1(n_161),
.B2(n_182),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_210),
.B1(n_194),
.B2(n_202),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_209),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_168),
.B1(n_184),
.B2(n_182),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_180),
.C(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_13),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_220),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_209),
.C(n_211),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_206),
.B(n_204),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_217),
.C(n_213),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_13),
.B(n_14),
.C(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_215),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_194),
.B(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_223),
.B(n_14),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_14),
.Y(n_230)
);


endmodule