module fake_jpeg_5263_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_46),
.B(n_47),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_33),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_51),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_26),
.B1(n_32),
.B2(n_17),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_19),
.B1(n_25),
.B2(n_18),
.Y(n_85)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_70),
.Y(n_93)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_25),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_25),
.A3(n_40),
.B1(n_42),
.B2(n_28),
.Y(n_78)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_32),
.B1(n_26),
.B2(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_32),
.B1(n_26),
.B2(n_38),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_33),
.C(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_84),
.B1(n_94),
.B2(n_66),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_24),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_87),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_29),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_51),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_29),
.B1(n_19),
.B2(n_13),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_64),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_18),
.B1(n_20),
.B2(n_25),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_66),
.B1(n_67),
.B2(n_58),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_102),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_48),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_111),
.C(n_106),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_108),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_51),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_65),
.B(n_47),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_122),
.B(n_57),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_65),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_47),
.C(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_59),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_120),
.B1(n_57),
.B2(n_72),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_87),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_79),
.C(n_95),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_92),
.B(n_75),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_78),
.B1(n_85),
.B2(n_74),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_131),
.B1(n_147),
.B2(n_150),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_75),
.B(n_83),
.C(n_73),
.Y(n_137)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_83),
.B1(n_54),
.B2(n_50),
.Y(n_141)
);

OR2x4_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_83),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_16),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_84),
.B1(n_94),
.B2(n_90),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_81),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_87),
.B1(n_88),
.B2(n_72),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_53),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_53),
.C(n_81),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_107),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_154),
.B(n_163),
.Y(n_206)
);

OAI22x1_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_108),
.B1(n_100),
.B2(n_109),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_16),
.B1(n_28),
.B2(n_23),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_179),
.B(n_146),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_98),
.B1(n_97),
.B2(n_71),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_164),
.B1(n_169),
.B2(n_175),
.Y(n_188)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_97),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_96),
.B1(n_70),
.B2(n_57),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_139),
.C(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_157),
.C(n_155),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_137),
.C(n_134),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_110),
.B1(n_99),
.B2(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_46),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_174),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_56),
.B1(n_77),
.B2(n_18),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_102),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_63),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_63),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_182),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_186),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_189),
.C(n_193),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_185),
.B(n_203),
.CI(n_175),
.CON(n_225),
.SN(n_225)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_194),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_127),
.C(n_132),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_165),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_144),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_198),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_129),
.B1(n_132),
.B2(n_137),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_159),
.B1(n_202),
.B2(n_198),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_129),
.A3(n_143),
.B1(n_126),
.B2(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_135),
.B1(n_125),
.B2(n_20),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_153),
.B1(n_163),
.B2(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_16),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_18),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_179),
.B(n_154),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_202),
.B1(n_180),
.B2(n_182),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_214),
.B1(n_229),
.B2(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_165),
.B1(n_153),
.B2(n_158),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_253)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_152),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_232),
.B1(n_20),
.B2(n_27),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_188),
.A2(n_159),
.B1(n_164),
.B2(n_161),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_184),
.C(n_193),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_238),
.C(n_239),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_195),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_249),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_189),
.C(n_224),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_185),
.C(n_200),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_230),
.B(n_207),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_243),
.B1(n_221),
.B2(n_233),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_196),
.C(n_206),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_190),
.C(n_63),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_16),
.C(n_20),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_250),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_27),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_28),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_223),
.C(n_218),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_0),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_253),
.B1(n_208),
.B2(n_207),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_225),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_259),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_218),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_231),
.B1(n_225),
.B2(n_215),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_269),
.B1(n_14),
.B2(n_13),
.Y(n_283)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_213),
.B1(n_211),
.B2(n_220),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_267),
.Y(n_287)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_271),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_244),
.C(n_249),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_246),
.B(n_15),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_238),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_274),
.A2(n_272),
.B(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_276),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_235),
.C(n_250),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_1),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_14),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_23),
.C(n_28),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_11),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_296),
.B(n_299),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_265),
.B1(n_261),
.B2(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_269),
.B1(n_264),
.B2(n_266),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_264),
.B1(n_2),
.B2(n_3),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_302),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_1),
.B(n_2),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_300),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_12),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_12),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_1),
.B(n_2),
.Y(n_301)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_4),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_280),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_308),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_278),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_277),
.Y(n_309)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_274),
.A3(n_275),
.B1(n_276),
.B2(n_11),
.C1(n_28),
.C2(n_9),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_300),
.B(n_8),
.Y(n_322)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_301),
.B(n_5),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_4),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_4),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_290),
.B(n_295),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_315),
.Y(n_324)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_305),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_322),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_295),
.B1(n_294),
.B2(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_313),
.C(n_304),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_325),
.A2(n_326),
.B(n_318),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_310),
.B(n_305),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_320),
.Y(n_329)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_330),
.A3(n_324),
.B1(n_323),
.B2(n_327),
.C1(n_9),
.C2(n_7),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_7),
.C(n_9),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_10),
.Y(n_333)
);


endmodule