module fake_jpeg_32079_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_28),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_0),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_57),
.B1(n_69),
.B2(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_85),
.B1(n_56),
.B2(n_55),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_62),
.B1(n_65),
.B2(n_46),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_68),
.B1(n_61),
.B2(n_67),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_84),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_92),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_48),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_69),
.B1(n_54),
.B2(n_65),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_101),
.B1(n_25),
.B2(n_41),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_51),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_62),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_103),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_53),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_49),
.CI(n_3),
.CON(n_106),
.SN(n_106)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_2),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_5),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_3),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_114),
.B(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_23),
.C(n_40),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_37),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_4),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_120),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_9),
.Y(n_124)
);

NOR4xp25_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_126),
.C(n_34),
.D(n_36),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_13),
.B(n_17),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_136),
.B(n_112),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_18),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_32),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_132),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_113),
.C(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_142),
.B(n_130),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_139),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_129),
.C(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_129),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_131),
.C(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_135),
.Y(n_152)
);


endmodule