module fake_aes_10095_n_667 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_667);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_667;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g89 ( .A(n_77), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_33), .Y(n_90) );
OR2x2_ASAP7_75t_L g91 ( .A(n_74), .B(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_31), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_76), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_36), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_85), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_30), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_80), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_10), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_50), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_64), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_88), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_55), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_2), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_44), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_79), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_1), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_78), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_37), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_53), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_17), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_56), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_16), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_40), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_28), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_54), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_65), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_59), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_9), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_11), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_60), .Y(n_127) );
INVxp67_ASAP7_75t_SL g128 ( .A(n_86), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_57), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_4), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_115), .B(n_0), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_130), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_132) );
NOR2x1_ASAP7_75t_L g133 ( .A(n_114), .B(n_3), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_130), .B(n_3), .Y(n_134) );
CKINVDCx11_ASAP7_75t_R g135 ( .A(n_94), .Y(n_135) );
CKINVDCx8_ASAP7_75t_R g136 ( .A(n_94), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_102), .B(n_5), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_115), .B(n_5), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_114), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_92), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_101), .Y(n_142) );
INVx4_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_108), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_101), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_92), .B(n_6), .Y(n_147) );
INVxp67_ASAP7_75t_L g148 ( .A(n_99), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_99), .B(n_7), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_100), .B(n_8), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_100), .B(n_9), .Y(n_153) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_96), .A2(n_41), .B(n_84), .Y(n_154) );
NAND2xp33_ASAP7_75t_SL g155 ( .A(n_91), .B(n_10), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_97), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_110), .B(n_11), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_101), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_143), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_143), .Y(n_160) );
OR2x2_ASAP7_75t_L g161 ( .A(n_134), .B(n_125), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_143), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_136), .B(n_90), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_139), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_148), .B(n_93), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_136), .B(n_98), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_155), .A2(n_126), .B1(n_110), .B2(n_117), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_140), .B(n_95), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_151), .A2(n_117), .B1(n_126), .B2(n_113), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_151), .B(n_91), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_140), .B(n_106), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_149), .B(n_107), .Y(n_180) );
NAND2xp33_ASAP7_75t_L g181 ( .A(n_149), .B(n_118), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_150), .B(n_121), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_152), .B(n_129), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_137), .B(n_105), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_153), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_137), .B(n_127), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_134), .B(n_150), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_159), .A2(n_154), .B(n_156), .Y(n_193) );
AND2x4_ASAP7_75t_SL g194 ( .A(n_165), .B(n_144), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_192), .B(n_133), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_192), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_166), .B(n_135), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_166), .B(n_156), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_177), .A2(n_138), .B1(n_131), .B2(n_133), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_177), .A2(n_157), .B1(n_147), .B2(n_113), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_191), .B(n_147), .Y(n_205) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_171), .B(n_157), .C(n_132), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_172), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_161), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_184), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_159), .A2(n_154), .B(n_122), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_172), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_177), .B(n_113), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_191), .B(n_111), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_167), .B(n_128), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_173), .B(n_97), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_185), .B(n_103), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_185), .B(n_103), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_162), .Y(n_218) );
OR2x6_ASAP7_75t_L g219 ( .A(n_184), .B(n_132), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_190), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_179), .B(n_180), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_161), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_184), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_184), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_174), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_185), .A2(n_113), .B1(n_141), .B2(n_109), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_162), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_162), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_186), .B(n_113), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_174), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_186), .A2(n_141), .B1(n_124), .B2(n_104), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_176), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_183), .B(n_104), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_162), .B(n_122), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_176), .B(n_123), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_227), .A2(n_190), .B(n_189), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_197), .B(n_169), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_197), .B(n_196), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_231), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_227), .A2(n_189), .B(n_188), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_199), .B(n_178), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_232), .A2(n_188), .B(n_187), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_196), .B(n_178), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_195), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_231), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_196), .B(n_164), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_195), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_194), .B(n_182), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_232), .A2(n_187), .B(n_182), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_200), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_220), .A2(n_163), .B(n_160), .Y(n_253) );
BUFx4f_ASAP7_75t_L g254 ( .A(n_219), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_234), .A2(n_163), .B(n_160), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_205), .A2(n_181), .B(n_175), .C(n_123), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_194), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
BUFx4f_ASAP7_75t_L g260 ( .A(n_219), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_199), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_199), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_193), .A2(n_154), .B(n_120), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_202), .A2(n_120), .B(n_109), .C(n_112), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_199), .B(n_101), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_219), .B(n_112), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_211), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_208), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_204), .B(n_113), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g270 ( .A1(n_219), .A2(n_116), .B1(n_119), .B2(n_124), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_209), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_216), .A2(n_116), .B1(n_119), .B2(n_129), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_208), .Y(n_274) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_210), .A2(n_158), .B(n_146), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_212), .A2(n_127), .B1(n_101), .B2(n_158), .Y(n_276) );
CKINVDCx8_ASAP7_75t_R g277 ( .A(n_198), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_217), .A2(n_158), .B(n_146), .C(n_14), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_237), .A2(n_146), .B(n_101), .Y(n_279) );
OAI22xp5_ASAP7_75t_SL g280 ( .A1(n_222), .A2(n_12), .B1(n_13), .B2(n_15), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_203), .A2(n_142), .B(n_43), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_254), .A2(n_228), .B1(n_212), .B2(n_215), .Y(n_282) );
CKINVDCx6p67_ASAP7_75t_R g283 ( .A(n_266), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_240), .B(n_209), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_252), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_268), .A2(n_222), .B1(n_206), .B2(n_233), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_223), .B(n_213), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_246), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_261), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_275), .A2(n_226), .B(n_236), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_263), .A2(n_226), .B(n_235), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_254), .A2(n_214), .B1(n_223), .B2(n_221), .Y(n_292) );
OAI22x1_ASAP7_75t_L g293 ( .A1(n_274), .A2(n_12), .B1(n_15), .B2(n_16), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_239), .B(n_224), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_238), .A2(n_224), .B(n_209), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_240), .B(n_224), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_242), .A2(n_244), .B(n_251), .Y(n_297) );
OR2x6_ASAP7_75t_L g298 ( .A(n_257), .B(n_229), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_SL g299 ( .A1(n_264), .A2(n_229), .B(n_48), .C(n_87), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_261), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_278), .A2(n_230), .B(n_225), .C(n_218), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_246), .Y(n_302) );
AOI222xp33_ASAP7_75t_L g303 ( .A1(n_280), .A2(n_142), .B1(n_18), .B2(n_19), .C1(n_20), .C2(n_17), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_261), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_260), .A2(n_142), .B1(n_225), .B2(n_218), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_260), .A2(n_142), .B1(n_225), .B2(n_218), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_249), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_243), .A2(n_230), .B(n_225), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_248), .A2(n_230), .B1(n_225), .B2(n_218), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_243), .A2(n_255), .B(n_249), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_259), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_266), .B(n_230), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g314 ( .A1(n_264), .A2(n_47), .B(n_83), .C(n_82), .Y(n_314) );
BUFx2_ASAP7_75t_SL g315 ( .A(n_277), .Y(n_315) );
AOI221xp5_ASAP7_75t_SL g316 ( .A1(n_273), .A2(n_256), .B1(n_269), .B2(n_247), .C(n_241), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_261), .B(n_230), .Y(n_317) );
OA21x2_ASAP7_75t_L g318 ( .A1(n_301), .A2(n_281), .B(n_279), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_311), .A2(n_265), .B(n_267), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_316), .A2(n_265), .B(n_276), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_285), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_286), .B(n_248), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_297), .A2(n_245), .B(n_262), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_294), .A2(n_270), .B(n_272), .C(n_250), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_304), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_312), .B(n_270), .Y(n_326) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_289), .B(n_271), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
OA21x2_ASAP7_75t_L g329 ( .A1(n_290), .A2(n_276), .B(n_142), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_291), .A2(n_272), .B(n_271), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_271), .B(n_262), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_282), .A2(n_271), .B(n_262), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_308), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_282), .B(n_262), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_287), .A2(n_218), .B(n_142), .C(n_20), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_303), .A2(n_18), .B1(n_19), .B2(n_21), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_289), .B(n_46), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_291), .A2(n_45), .B(n_75), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_296), .Y(n_342) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_295), .A2(n_42), .B(n_71), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_284), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_317), .A2(n_39), .B(n_69), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_292), .A2(n_38), .B(n_68), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_317), .A2(n_35), .B(n_67), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_330), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_332), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_321), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_328), .B(n_335), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_334), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_326), .B(n_298), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
BUFx5_ASAP7_75t_L g357 ( .A(n_337), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_329), .Y(n_359) );
OAI322xp33_ASAP7_75t_L g360 ( .A1(n_322), .A2(n_292), .A3(n_303), .B1(n_293), .B2(n_306), .C1(n_307), .C2(n_310), .Y(n_360) );
NAND3xp33_ASAP7_75t_L g361 ( .A(n_338), .B(n_314), .C(n_299), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_340), .B(n_306), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_331), .A2(n_307), .B(n_309), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_336), .Y(n_364) );
OA21x2_ASAP7_75t_L g365 ( .A1(n_323), .A2(n_284), .B(n_313), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_337), .B(n_298), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_335), .B(n_300), .Y(n_367) );
OA21x2_ASAP7_75t_L g368 ( .A1(n_319), .A2(n_313), .B(n_300), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_332), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_342), .B(n_305), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_329), .Y(n_372) );
AOI21x1_ASAP7_75t_L g373 ( .A1(n_318), .A2(n_298), .B(n_305), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_342), .B(n_315), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_339), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_375), .B(n_325), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_350), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_375), .B(n_325), .Y(n_382) );
INVx4_ASAP7_75t_L g383 ( .A(n_362), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_348), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_353), .B(n_333), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_357), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_358), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_356), .B(n_347), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_356), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_351), .B(n_352), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_375), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_357), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_355), .B(n_324), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_357), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_357), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_355), .B(n_344), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_351), .B(n_344), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_357), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_352), .B(n_320), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_364), .B(n_320), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_357), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_364), .B(n_320), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_357), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_366), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_357), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_357), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_357), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_358), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_366), .B(n_320), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_383), .B(n_373), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_391), .B(n_354), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_393), .B(n_365), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_393), .B(n_365), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_395), .B(n_365), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_391), .B(n_354), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_395), .B(n_365), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
INVx4_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_377), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_383), .B(n_373), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_379), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_381), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_398), .B(n_374), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_383), .B(n_356), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_404), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_405), .B(n_365), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_386), .A2(n_362), .B(n_361), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_388), .B(n_359), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
AOI21xp33_ASAP7_75t_SL g434 ( .A1(n_396), .A2(n_349), .B(n_370), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_377), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_404), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_396), .B(n_359), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_380), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_399), .B(n_359), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_399), .B(n_372), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_402), .B(n_372), .Y(n_442) );
NAND4xp25_ASAP7_75t_L g443 ( .A(n_394), .B(n_374), .C(n_376), .D(n_367), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_378), .Y(n_444) );
NOR2x1p5_ASAP7_75t_L g445 ( .A(n_383), .B(n_372), .Y(n_445) );
NOR4xp25_ASAP7_75t_SL g446 ( .A(n_402), .B(n_360), .C(n_362), .D(n_340), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_404), .B(n_367), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_380), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_398), .B(n_371), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_380), .B(n_371), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_408), .B(n_368), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_406), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_378), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_405), .B(n_368), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_382), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_408), .B(n_369), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_382), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_383), .B(n_356), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_382), .B(n_371), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_406), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_385), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_439), .B(n_407), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_419), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_413), .B(n_392), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_439), .B(n_407), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_448), .B(n_407), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_419), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_448), .B(n_397), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_456), .B(n_392), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_456), .B(n_410), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_462), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_420), .B(n_390), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_458), .B(n_410), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_458), .B(n_424), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_425), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_425), .B(n_409), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_430), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_420), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_434), .B(n_360), .C(n_361), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_430), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_437), .B(n_409), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_413), .B(n_397), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_443), .B(n_394), .C(n_397), .D(n_411), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_417), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_417), .B(n_426), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_451), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_460), .Y(n_491) );
NOR2x1_ASAP7_75t_L g492 ( .A(n_420), .B(n_362), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_447), .B(n_403), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_420), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_450), .B(n_385), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_434), .B(n_394), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_432), .B(n_403), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_447), .B(n_385), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_432), .Y(n_500) );
OR2x6_ASAP7_75t_L g501 ( .A(n_445), .B(n_362), .Y(n_501) );
OAI211xp5_ASAP7_75t_L g502 ( .A1(n_431), .A2(n_411), .B(n_346), .C(n_401), .Y(n_502) );
OAI21xp33_ASAP7_75t_L g503 ( .A1(n_414), .A2(n_400), .B(n_401), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_436), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_438), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_428), .B(n_403), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_438), .B(n_401), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_440), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_428), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_452), .B(n_400), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_453), .Y(n_511) );
NAND2xp33_ASAP7_75t_SL g512 ( .A(n_445), .B(n_400), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_436), .B(n_345), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_440), .Y(n_514) );
NOR2xp33_ASAP7_75t_SL g515 ( .A(n_453), .B(n_340), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_452), .B(n_387), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_387), .Y(n_517) );
NOR2x1_ASAP7_75t_SL g518 ( .A(n_461), .B(n_387), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_441), .B(n_384), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_441), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_442), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_442), .B(n_384), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_489), .B(n_429), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_488), .B(n_418), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_477), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_477), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_464), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_486), .A2(n_415), .B1(n_418), .B2(n_414), .Y(n_530) );
AOI21xp33_ASAP7_75t_SL g531 ( .A1(n_482), .A2(n_429), .B(n_415), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_490), .B(n_416), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_499), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_491), .B(n_416), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_506), .B(n_455), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_469), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_509), .Y(n_537) );
OAI32xp33_ASAP7_75t_L g538 ( .A1(n_512), .A2(n_436), .A3(n_449), .B1(n_455), .B2(n_457), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_505), .B(n_412), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_473), .B(n_421), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_518), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_474), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_470), .B(n_421), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g544 ( .A1(n_496), .A2(n_412), .B(n_422), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_478), .Y(n_545) );
AND4x1_ASAP7_75t_L g546 ( .A(n_492), .B(n_446), .C(n_341), .D(n_22), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_500), .B(n_421), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_508), .B(n_422), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_480), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_483), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_514), .B(n_520), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_485), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_517), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_471), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_511), .A2(n_436), .B(n_449), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_521), .B(n_449), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_510), .B(n_454), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_510), .B(n_422), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_516), .Y(n_560) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_504), .B(n_412), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_516), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_497), .B(n_449), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_504), .B(n_412), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_497), .B(n_433), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_498), .B(n_422), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_501), .B(n_459), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_507), .B(n_433), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_501), .A2(n_446), .B1(n_369), .B2(n_454), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_493), .B(n_459), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_471), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_501), .B(n_459), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_498), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_495), .B(n_433), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g575 ( .A(n_481), .B(n_494), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_561), .A2(n_515), .B(n_476), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_537), .B(n_472), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_531), .A2(n_503), .B1(n_502), .B2(n_472), .C(n_476), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_526), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_527), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_524), .Y(n_581) );
AOI21xp33_ASAP7_75t_SL g582 ( .A1(n_561), .A2(n_475), .B(n_513), .Y(n_582) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_541), .A2(n_475), .B(n_513), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_555), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_571), .B(n_468), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_529), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_536), .Y(n_587) );
XNOR2xp5_ASAP7_75t_L g588 ( .A(n_553), .B(n_467), .Y(n_588) );
OAI32xp33_ASAP7_75t_L g589 ( .A1(n_541), .A2(n_522), .A3(n_519), .B1(n_484), .B2(n_479), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_564), .B(n_519), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_542), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_545), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_573), .A2(n_484), .B1(n_479), .B2(n_522), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_557), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_563), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_R g596 ( .A1(n_523), .A2(n_454), .B(n_444), .C(n_435), .Y(n_596) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_573), .A2(n_463), .B1(n_369), .B2(n_444), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_549), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_550), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_530), .A2(n_459), .B1(n_427), .B2(n_435), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_552), .Y(n_601) );
CKINVDCx8_ASAP7_75t_R g602 ( .A(n_564), .Y(n_602) );
INVxp67_ASAP7_75t_SL g603 ( .A(n_575), .Y(n_603) );
OAI22xp33_ASAP7_75t_SL g604 ( .A1(n_566), .A2(n_427), .B1(n_389), .B2(n_435), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_539), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_559), .B(n_570), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_533), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_551), .Y(n_608) );
NOR3xp33_ASAP7_75t_SL g609 ( .A(n_569), .B(n_538), .C(n_566), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_551), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_565), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_578), .A2(n_530), .B1(n_544), .B2(n_572), .Y(n_612) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_602), .A2(n_556), .B(n_557), .C(n_573), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_603), .A2(n_564), .B(n_547), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_600), .A2(n_572), .B1(n_567), .B2(n_559), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g617 ( .A1(n_582), .A2(n_546), .B(n_572), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_604), .A2(n_567), .B(n_548), .C(n_539), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_596), .A2(n_528), .B1(n_548), .B2(n_525), .C(n_532), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_603), .A2(n_567), .B(n_570), .C(n_535), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_589), .A2(n_558), .B(n_534), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_593), .A2(n_535), .B1(n_560), .B2(n_562), .C(n_554), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_593), .A2(n_560), .B1(n_562), .B2(n_554), .C(n_574), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_594), .A2(n_543), .B1(n_565), .B2(n_568), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_594), .A2(n_568), .B1(n_540), .B2(n_427), .Y(n_625) );
NAND4xp75_ASAP7_75t_L g626 ( .A(n_609), .B(n_368), .C(n_363), .D(n_343), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_580), .Y(n_627) );
OAI321xp33_ASAP7_75t_L g628 ( .A1(n_581), .A2(n_444), .A3(n_384), .B1(n_378), .B2(n_369), .C(n_363), .Y(n_628) );
NOR4xp25_ASAP7_75t_L g629 ( .A(n_581), .B(n_390), .C(n_23), .D(n_368), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_607), .A2(n_427), .B1(n_390), .B2(n_389), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_576), .A2(n_389), .B1(n_369), .B2(n_390), .Y(n_631) );
OAI21xp33_ASAP7_75t_SL g632 ( .A1(n_590), .A2(n_345), .B(n_347), .Y(n_632) );
AOI31xp33_ASAP7_75t_SL g633 ( .A1(n_588), .A2(n_25), .A3(n_26), .B(n_27), .Y(n_633) );
NAND3x1_ASAP7_75t_L g634 ( .A(n_614), .B(n_577), .C(n_609), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_612), .B(n_583), .C(n_585), .D(n_611), .Y(n_635) );
OAI21xp33_ASAP7_75t_L g636 ( .A1(n_615), .A2(n_584), .B(n_592), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_622), .A2(n_586), .B1(n_587), .B2(n_591), .C(n_601), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_616), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_623), .A2(n_598), .B1(n_599), .B2(n_597), .C(n_610), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_617), .A2(n_608), .B(n_595), .C(n_606), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_621), .A2(n_597), .B1(n_605), .B2(n_371), .C(n_389), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_613), .B(n_390), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_620), .A2(n_327), .B(n_389), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g644 ( .A1(n_618), .A2(n_29), .B(n_32), .C(n_34), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_629), .A2(n_368), .B(n_343), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_627), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_637), .B(n_619), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_640), .A2(n_631), .B1(n_625), .B2(n_632), .C(n_633), .Y(n_648) );
NAND4xp25_ASAP7_75t_SL g649 ( .A(n_641), .B(n_631), .C(n_624), .D(n_626), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_639), .B(n_630), .C(n_628), .Y(n_650) );
OR5x1_ASAP7_75t_L g651 ( .A(n_635), .B(n_49), .C(n_51), .D(n_52), .E(n_58), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_636), .B(n_356), .Y(n_652) );
AOI211x1_ASAP7_75t_L g653 ( .A1(n_634), .A2(n_62), .B(n_63), .C(n_66), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_647), .B(n_638), .Y(n_654) );
NAND2x1p5_ASAP7_75t_SL g655 ( .A(n_653), .B(n_644), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_650), .B(n_646), .Y(n_656) );
NAND4xp75_ASAP7_75t_L g657 ( .A(n_652), .B(n_642), .C(n_643), .D(n_645), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_656), .B(n_649), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_654), .B(n_648), .C(n_655), .D(n_651), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_657), .Y(n_660) );
XOR2x1_ASAP7_75t_L g661 ( .A(n_660), .B(n_657), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_658), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_659), .B1(n_356), .B2(n_327), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_661), .B(n_81), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_343), .B(n_318), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_343), .B(n_318), .Y(n_666) );
AOI21xp33_ASAP7_75t_SL g667 ( .A1(n_666), .A2(n_318), .B(n_369), .Y(n_667) );
endmodule