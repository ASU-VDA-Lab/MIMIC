module fake_jpeg_17561_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_12),
.B(n_11),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_SL g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_10),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_61),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_53),
.B1(n_47),
.B2(n_46),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_66),
.B1(n_71),
.B2(n_6),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_51),
.B1(n_54),
.B2(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_74),
.B1(n_43),
.B2(n_17),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_50),
.B1(n_51),
.B2(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_2),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_54),
.B1(n_48),
.B2(n_5),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_80),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_88),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_7),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_8),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_91),
.B1(n_75),
.B2(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_64),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_81),
.B1(n_86),
.B2(n_76),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_87),
.B1(n_95),
.B2(n_94),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_108),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_100),
.B1(n_99),
.B2(n_85),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_92),
.B1(n_97),
.B2(n_79),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_111),
.B1(n_109),
.B2(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_82),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_117),
.B1(n_78),
.B2(n_23),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_114),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_120),
.B(n_118),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_119),
.C(n_115),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_26),
.B(n_27),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_28),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_29),
.C(n_30),
.Y(n_126)
);

AOI21x1_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_31),
.B(n_33),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_38),
.B(n_37),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_36),
.Y(n_129)
);


endmodule