module fake_jpeg_13261_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_10),
.B(n_16),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_6),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_20),
.B(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.C(n_72),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_0),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_50),
.Y(n_77)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_52),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_18),
.C(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_63),
.B1(n_45),
.B2(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_91),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_59),
.B(n_58),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_97),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_49),
.Y(n_92)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_4),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_95),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_98),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_61),
.B(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_1),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_2),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_117),
.B(n_33),
.Y(n_128)
);

NOR4xp25_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_29),
.C(n_39),
.D(n_38),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_43),
.C(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_118),
.B(n_121),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_107),
.B1(n_106),
.B2(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_12),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_17),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_125),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_21),
.B(n_30),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_31),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.C(n_35),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_132),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_110),
.B1(n_112),
.B2(n_115),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_124),
.C(n_122),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_136),
.A2(n_138),
.B(n_129),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_123),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_137),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.C(n_135),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_119),
.Y(n_145)
);


endmodule