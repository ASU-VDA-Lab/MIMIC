module fake_jpeg_23614_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g77 ( 
.A(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_9),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_63),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_31),
.B1(n_36),
.B2(n_29),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_55),
.B(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_31),
.B1(n_25),
.B2(n_36),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_29),
.B1(n_31),
.B2(n_23),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_26),
.B(n_34),
.C(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_59),
.B(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_25),
.B1(n_36),
.B2(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_30),
.B1(n_23),
.B2(n_32),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_69),
.B(n_21),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_30),
.B1(n_23),
.B2(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_22),
.B1(n_37),
.B2(n_27),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_72),
.B1(n_46),
.B2(n_48),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_27),
.B1(n_37),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_19),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_46),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_37),
.B1(n_27),
.B2(n_20),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_20),
.B1(n_24),
.B2(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_89),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_80),
.A2(n_95),
.B1(n_78),
.B2(n_50),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_98),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_48),
.C(n_43),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_63),
.C(n_51),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_48),
.CI(n_41),
.CON(n_89),
.SN(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_45),
.B1(n_40),
.B2(n_24),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_116),
.B1(n_78),
.B2(n_57),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_101),
.B(n_2),
.Y(n_147)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_97),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_35),
.B1(n_45),
.B2(n_40),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_104),
.B1(n_107),
.B2(n_71),
.Y(n_125)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_41),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_100),
.B(n_109),
.Y(n_148)
);

OR2x4_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_43),
.Y(n_102)
);

FAx1_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_3),
.CI(n_4),
.CON(n_149),
.SN(n_149)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_35),
.B1(n_45),
.B2(n_38),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_18),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_34),
.B1(n_24),
.B2(n_26),
.Y(n_107)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_18),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_115),
.Y(n_129)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_34),
.B1(n_26),
.B2(n_41),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_77),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_139),
.C(n_140),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_50),
.B1(n_60),
.B2(n_57),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_118),
.A2(n_114),
.B1(n_110),
.B2(n_97),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_133),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_72),
.B1(n_69),
.B2(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_43),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_43),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_0),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_106),
.B(n_113),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_43),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_79),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_91),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_80),
.A2(n_42),
.B1(n_1),
.B2(n_3),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_146),
.C(n_128),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_42),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_103),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_42),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_87),
.B(n_116),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_99),
.B(n_103),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_145),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_93),
.B(n_87),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_164),
.B(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_159),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_98),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_167),
.B(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

XOR2x1_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_3),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_137),
.B(n_104),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_4),
.Y(n_199)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_89),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_99),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_89),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_117),
.B(n_108),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_127),
.A3(n_149),
.B1(n_147),
.B2(n_126),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_107),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_130),
.B1(n_100),
.B2(n_121),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_130),
.B1(n_88),
.B2(n_82),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_190),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_118),
.B1(n_135),
.B2(n_88),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_185),
.B1(n_197),
.B2(n_177),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_135),
.B1(n_124),
.B2(n_136),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_204),
.B1(n_205),
.B2(n_165),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_120),
.B(n_122),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_208),
.B(n_176),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_194),
.B(n_200),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_123),
.B(n_91),
.C(n_141),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_153),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_111),
.B1(n_91),
.B2(n_6),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_161),
.C(n_170),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_156),
.C(n_150),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_5),
.B(n_6),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_172),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_212),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_153),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_232),
.C(n_191),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_215),
.B1(n_218),
.B2(n_184),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_225),
.Y(n_236)
);

BUFx12_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_222),
.Y(n_241)
);

BUFx12f_ASAP7_75t_SL g220 ( 
.A(n_208),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_220),
.A2(n_223),
.B1(n_229),
.B2(n_163),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_166),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_152),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_179),
.B1(n_174),
.B2(n_159),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_228),
.B1(n_210),
.B2(n_183),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_231),
.C(n_182),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_179),
.B1(n_174),
.B2(n_157),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_171),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_174),
.C(n_158),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_238),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_204),
.B1(n_188),
.B2(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_216),
.B(n_187),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_244),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_193),
.C(n_158),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_217),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_188),
.B1(n_202),
.B2(n_205),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_193),
.B1(n_202),
.B2(n_194),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_248),
.B1(n_194),
.B2(n_212),
.Y(n_257)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_216),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_225),
.B(n_167),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_194),
.B1(n_175),
.B2(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_245),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_227),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_253),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_162),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_261),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_262),
.B(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_260),
.A2(n_263),
.B1(n_186),
.B2(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_241),
.B(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_154),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_219),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_194),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_219),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_242),
.C(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_278),
.C(n_224),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_275),
.B(n_273),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_233),
.B1(n_239),
.B2(n_234),
.Y(n_273)
);

AO22x1_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_276),
.B1(n_265),
.B2(n_252),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_237),
.B1(n_230),
.B2(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_236),
.C(n_224),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_274),
.A2(n_259),
.B1(n_256),
.B2(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_283),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_10),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_271),
.A2(n_257),
.B(n_259),
.C(n_258),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_284),
.B(n_10),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_269),
.B1(n_277),
.B2(n_272),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_251),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_260),
.B1(n_278),
.B2(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_293),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_8),
.B(n_9),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_281),
.B(n_12),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_11),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_17),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_281),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_297),
.A2(n_293),
.B1(n_290),
.B2(n_13),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_SL g302 ( 
.A1(n_299),
.A2(n_300),
.B(n_294),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.Y(n_304)
);

NAND4xp25_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_298),
.C(n_296),
.D(n_15),
.Y(n_303)
);

OAI221xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.C(n_17),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_11),
.Y(n_306)
);


endmodule