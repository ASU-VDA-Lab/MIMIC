module real_jpeg_25279_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_0),
.B(n_48),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_0),
.B(n_68),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_0),
.B(n_50),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_0),
.B(n_32),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_0),
.B(n_27),
.Y(n_244)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_7),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_7),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_7),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_7),
.B(n_32),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_7),
.B(n_53),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_8),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_50),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_8),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_48),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_10),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_10),
.B(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_68),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_10),
.B(n_272),
.Y(n_271)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_12),
.B(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_12),
.B(n_68),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_12),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_12),
.B(n_32),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_12),
.B(n_53),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_12),
.B(n_50),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_13),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_13),
.B(n_32),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_13),
.B(n_53),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_36),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_13),
.B(n_50),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_13),
.B(n_48),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_13),
.B(n_68),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_14),
.B(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_14),
.B(n_50),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_14),
.B(n_48),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_14),
.B(n_53),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_14),
.B(n_32),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_14),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_14),
.B(n_68),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_14),
.B(n_27),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_15),
.B(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_15),
.B(n_32),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_15),
.B(n_53),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_16),
.B(n_53),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_16),
.B(n_50),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_16),
.B(n_32),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_186),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_16),
.B(n_48),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_16),
.B(n_68),
.Y(n_273)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_17),
.Y(n_115)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_17),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_151),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.C(n_91),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_21),
.B(n_79),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_22),
.B(n_56),
.C(n_73),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_46),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_23),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_29),
.C(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_26),
.B(n_62),
.Y(n_126)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_29),
.A2(n_39),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_29),
.B(n_81),
.C(n_84),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_30),
.B(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_31),
.B(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_34),
.A2(n_38),
.B1(n_41),
.B2(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_37),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_41),
.C(n_42),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_40),
.B(n_46),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_41),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_42),
.A2(n_43),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_45),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_45),
.B(n_216),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_46),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.CI(n_52),
.CON(n_46),
.SN(n_46)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_49),
.C(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_53),
.Y(n_217)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_73),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_67),
.C(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_58),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_64),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_64),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_71),
.B1(n_77),
.B2(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_67),
.B(n_76),
.C(n_78),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_86),
.C(n_87),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_84),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_87),
.Y(n_333)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.CI(n_90),
.CON(n_87),
.SN(n_87)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_91),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_105),
.C(n_109),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_92),
.B(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_101),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_93),
.B(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_95),
.B(n_101),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_98),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_105),
.B(n_109),
.Y(n_326)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_117),
.C(n_118),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_110),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_110),
.B(n_315),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.CI(n_116),
.CON(n_110),
.SN(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_117),
.B(n_118),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_134),
.B2(n_135),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_128),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_328),
.C(n_329),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_318),
.C(n_319),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_304),
.C(n_305),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_282),
.C(n_283),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_251),
.C(n_252),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_226),
.C(n_227),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_188),
.C(n_199),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_172),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_167),
.C(n_172),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_165),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_162),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_168),
.B(n_170),
.C(n_171),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_180),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_173),
.B(n_181),
.C(n_182),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_177),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_187),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_198),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_193),
.B1(n_198),
.B2(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_222),
.C(n_223),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_208),
.C(n_213),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_206),
.C(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_214)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.C(n_218),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_240),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_241),
.C(n_250),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_235),
.C(n_236),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_234),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_236),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.CI(n_239),
.CON(n_236),
.SN(n_236)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_250),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_248),
.B2(n_249),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_244),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_267),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_256),
.C(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_263),
.C(n_266),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_258),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.CI(n_261),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_275),
.C(n_280),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_275),
.B1(n_280),
.B2(n_281),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_270),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_273),
.B(n_274),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_273),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_301),
.C(n_302),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_275),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_278),
.C(n_279),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_297),
.B2(n_303),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_298),
.C(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_295),
.C(n_296),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_316),
.B2(n_317),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_310),
.C(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_322),
.C(n_327),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_327),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);


endmodule