module fake_jpeg_24778_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_9),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_0),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_13),
.B(n_17),
.C(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_27),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_10),
.B1(n_19),
.B2(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_7),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_15),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_10),
.B1(n_17),
.B2(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_7),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_27),
.B(n_26),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_49),
.C(n_46),
.Y(n_53)
);

AO22x2_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_29),
.B1(n_32),
.B2(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_39),
.B1(n_40),
.B2(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_42),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_59),
.B1(n_41),
.B2(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_39),
.C(n_36),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_50),
.C(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_45),
.B1(n_48),
.B2(n_46),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_64),
.B1(n_54),
.B2(n_57),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_47),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_63),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_67),
.CON(n_70),
.SN(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_71),
.Y(n_74)
);


endmodule