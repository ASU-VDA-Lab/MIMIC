module real_jpeg_29459_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_202;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g60 ( 
.A(n_0),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_1),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_9),
.B1(n_24),
.B2(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_4),
.A2(n_28),
.B1(n_41),
.B2(n_43),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_4),
.A2(n_28),
.B1(n_58),
.B2(n_59),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_41),
.B1(n_43),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_74)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_9),
.B1(n_24),
.B2(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_8),
.A2(n_31),
.B1(n_41),
.B2(n_43),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_8),
.A2(n_9),
.B(n_23),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_8),
.A2(n_31),
.B1(n_58),
.B2(n_59),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_8),
.B(n_21),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_8),
.A2(n_10),
.B(n_41),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_8),
.A2(n_55),
.B(n_59),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_8),
.B(n_40),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_9),
.A2(n_11),
.B1(n_24),
.B2(n_39),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_9),
.A2(n_10),
.B1(n_24),
.B2(n_42),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_9),
.A2(n_31),
.B(n_160),
.C(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_99)
);

XNOR2x2_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_109),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_107),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_15),
.B(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_71),
.B1(n_72),
.B2(n_89),
.Y(n_15)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_63),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_34),
.B2(n_35),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_18),
.A2(n_19),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_18),
.A2(n_19),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_18),
.B(n_222),
.C(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_19),
.B(n_106),
.C(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_29),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_32),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_21),
.A2(n_30),
.B1(n_32),
.B2(n_104),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_22),
.A2(n_27),
.B(n_31),
.C(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_30),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_31),
.A2(n_41),
.B(n_56),
.C(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_31),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_31),
.B(n_57),
.Y(n_198)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B(n_44),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_40),
.B(n_47),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_68),
.B(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_52),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_57),
.B1(n_84),
.B2(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_65),
.B(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_58),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_66),
.A2(n_103),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_66),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_66),
.B(n_150),
.C(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_66),
.A2(n_117),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_69),
.B(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_80),
.B(n_85),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_85),
.B1(n_86),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_73),
.A2(n_81),
.B1(n_93),
.B2(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_77),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_76),
.B(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_100),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_81),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_83),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.C(n_95),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_91),
.B(n_94),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_95),
.A2(n_96),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.C(n_105),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_97),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_98),
.A2(n_101),
.B1(n_175),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_98),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_123),
.B(n_140),
.Y(n_150)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_101),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_101),
.A2(n_175),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_101),
.B(n_122),
.C(n_185),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_101),
.B(n_166),
.C(n_174),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_103),
.B(n_117),
.C(n_118),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_116),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_106),
.B1(n_128),
.B2(n_129),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_134),
.C(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_105),
.A2(n_106),
.B1(n_133),
.B2(n_134),
.Y(n_205)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_242),
.B(n_247),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_230),
.B(n_241),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_153),
.B(n_214),
.C(n_229),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_143),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_113),
.B(n_143),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_125),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_114),
.B(n_126),
.C(n_132),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_122),
.A2(n_148),
.B1(n_183),
.B2(n_186),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_122),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_198),
.Y(n_199)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_134),
.B1(n_180),
.B2(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_133),
.B(n_138),
.Y(n_222)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_134),
.B(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_144),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_149),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_213),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_208),
.B(n_212),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_176),
.B(n_207),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_157),
.B(n_165),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_171),
.B2(n_172),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_168),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_202),
.B(n_206),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_187),
.B(n_201),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_182),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B(n_200),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_197),
.B(n_199),
.Y(n_191)
);

INVx5_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_227),
.B2(n_228),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_221),
.C(n_228),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_227),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_232),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_238),
.C(n_240),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);


endmodule