module fake_jpeg_21472_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_60),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_86),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_23),
.B1(n_49),
.B2(n_44),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_0),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_65),
.Y(n_102)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_52),
.B1(n_64),
.B2(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_99),
.B1(n_68),
.B2(n_75),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_66),
.Y(n_116)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_77),
.B1(n_76),
.B2(n_59),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_67),
.B1(n_66),
.B2(n_77),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_95),
.B1(n_58),
.B2(n_76),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_75),
.B1(n_68),
.B2(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_70),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_110),
.B1(n_57),
.B2(n_103),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_106),
.B1(n_108),
.B2(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_130),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_133),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_139),
.B1(n_8),
.B2(n_11),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_72),
.B1(n_56),
.B2(n_59),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_65),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_136),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_24),
.C(n_42),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_143),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_20),
.B1(n_41),
.B2(n_40),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_140),
.B(n_141),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_8),
.B(n_10),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_27),
.B1(n_39),
.B2(n_37),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_18),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_28),
.C(n_51),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_153),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_25),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_150),
.Y(n_158)
);

XOR2x1_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_154),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_146),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_147),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_161),
.B(n_147),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_158),
.C(n_160),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_166),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_162),
.C(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_32),
.B(n_35),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_30),
.B(n_34),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_15),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_16),
.B(n_148),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_121),
.B(n_13),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_121),
.Y(n_178)
);


endmodule