module fake_jpeg_22482_n_234 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_23),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_27),
.B1(n_19),
.B2(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_32),
.B1(n_33),
.B2(n_15),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_27),
.B1(n_24),
.B2(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_21),
.B1(n_15),
.B2(n_18),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_22),
.C(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_24),
.B1(n_34),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_62),
.B1(n_52),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_64),
.B1(n_68),
.B2(n_48),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_66),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_0),
.B(n_1),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_34),
.B(n_29),
.C(n_30),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_76),
.B1(n_70),
.B2(n_74),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_23),
.B1(n_22),
.B2(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_23),
.B1(n_22),
.B2(n_17),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_47),
.B1(n_31),
.B2(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_85),
.B1(n_60),
.B2(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_84),
.Y(n_118)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_55),
.B1(n_51),
.B2(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_91),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_50),
.B(n_55),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_67),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_93),
.Y(n_116)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_97),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_0),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_10),
.C(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_53),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_112),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_90),
.C(n_82),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_78),
.C(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_69),
.B1(n_42),
.B2(n_58),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_69),
.B1(n_97),
.B2(n_79),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_117),
.B1(n_25),
.B2(n_16),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_127),
.C(n_130),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_67),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_99),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_99),
.C(n_86),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_13),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_140),
.B(n_104),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_83),
.C(n_46),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_122),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_73),
.B(n_65),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_107),
.B(n_113),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_58),
.B1(n_65),
.B2(n_87),
.Y(n_136)
);

OAI22x1_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_87),
.B1(n_107),
.B2(n_100),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_138),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_25),
.C(n_16),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_26),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_144),
.B(n_149),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_134),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_119),
.A3(n_106),
.B1(n_105),
.B2(n_100),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_158),
.B1(n_139),
.B2(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_153),
.B1(n_156),
.B2(n_3),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_16),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_26),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_127),
.C(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_164),
.C(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_160),
.B1(n_144),
.B2(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_139),
.C(n_131),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_26),
.B1(n_1),
.B2(n_3),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_26),
.C(n_1),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_171),
.C(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_2),
.C(n_3),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_2),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_154),
.B1(n_143),
.B2(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_147),
.Y(n_184)
);

XOR2x2_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_174),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_149),
.B1(n_155),
.B2(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_4),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_167),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_168),
.C(n_162),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_7),
.C(n_8),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_171),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_SL g203 ( 
.A(n_195),
.B(n_196),
.C(n_199),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_170),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_187),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_5),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_183),
.C(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_8),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_180),
.B1(n_177),
.B2(n_179),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_207),
.B1(n_198),
.B2(n_193),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_177),
.B1(n_185),
.B2(n_181),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_182),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_8),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_182),
.B(n_183),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_195),
.B(n_10),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_217),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_216),
.C(n_204),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_202),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_208),
.B(n_209),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_213),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_225),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_226),
.C(n_220),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_206),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_230),
.B(n_219),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_12),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_12),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_12),
.Y(n_234)
);


endmodule