module real_jpeg_28067_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_325, n_11, n_14, n_7, n_3, n_5, n_4, n_324, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_325;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_324;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_0),
.A2(n_62),
.B1(n_63),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_0),
.A2(n_32),
.B(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_0),
.B(n_67),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_0),
.A2(n_35),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_0),
.B(n_35),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_0),
.B(n_91),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_0),
.A2(n_102),
.B1(n_104),
.B2(n_174),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_0),
.A2(n_31),
.B(n_190),
.Y(n_189)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_2),
.A2(n_42),
.B1(n_62),
.B2(n_63),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_42),
.B1(n_53),
.B2(n_55),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_42),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_53),
.B1(n_55),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_84),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_84),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_84),
.Y(n_294)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_47),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_5),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_5),
.A2(n_47),
.B1(n_62),
.B2(n_63),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_7),
.A2(n_53),
.B1(n_55),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_7),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_127),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_127),
.Y(n_297)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_9),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_9),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_10),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_40),
.B1(n_53),
.B2(n_55),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_53),
.B1(n_55),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_11),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_106),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_106),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_106),
.Y(n_317)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_13),
.A2(n_53),
.B1(n_55),
.B2(n_73),
.Y(n_174)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_17),
.A2(n_53),
.B1(n_55),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_17),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_17),
.A2(n_35),
.B1(n_36),
.B2(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_17),
.A2(n_62),
.B1(n_63),
.B2(n_82),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_305),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_274),
.A3(n_301),
.B1(n_303),
.B2(n_304),
.C(n_324),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_225),
.A3(n_263),
.B1(n_268),
.B2(n_273),
.C(n_325),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_119),
.C(n_138),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_95),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_23),
.B(n_95),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_74),
.C(n_85),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_24),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_60),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_26),
.B(n_44),
.C(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_27)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_28),
.A2(n_34),
.B1(n_41),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_28),
.A2(n_34),
.B1(n_89),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_28),
.A2(n_34),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_28),
.A2(n_34),
.B(n_313),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_29),
.A2(n_31),
.A3(n_36),
.B1(n_191),
.B2(n_199),
.Y(n_198)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_31),
.A2(n_32),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_32),
.B(n_70),
.Y(n_191)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_35),
.A2(n_51),
.A3(n_55),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_35),
.B(n_37),
.Y(n_199)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_39),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B1(n_57),
.B2(n_59),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_48),
.A2(n_59),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_48),
.A2(n_59),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_50),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_49),
.A2(n_50),
.B1(n_100),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_49),
.A2(n_50),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_49),
.A2(n_50),
.B1(n_148),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_49),
.A2(n_50),
.B1(n_238),
.B2(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_49),
.A2(n_50),
.B(n_250),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_50),
.B(n_70),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_52),
.B(n_53),
.Y(n_152)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_53),
.B(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_57),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_60)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_67),
.B1(n_114),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_61),
.A2(n_67),
.B1(n_134),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_61),
.A2(n_67),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_65),
.Y(n_66)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_68),
.B(n_70),
.C(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_70),
.B(n_104),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_74),
.A2(n_85),
.B1(n_86),
.B2(n_223),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_74),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_77),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_78),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_79),
.Y(n_175)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_94),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_87),
.B(n_210),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_91),
.B1(n_117),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_90),
.A2(n_91),
.B1(n_136),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_90),
.A2(n_91),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_90),
.A2(n_91),
.B1(n_283),
.B2(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_92),
.B(n_94),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_93),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_108),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_107),
.C(n_108),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_101),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_104),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_102),
.A2(n_167),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_102),
.A2(n_104),
.B1(n_162),
.B2(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_102),
.A2(n_104),
.B(n_126),
.Y(n_240)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_118),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_115),
.C(n_118),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_111),
.A2(n_112),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_111),
.A2(n_112),
.B1(n_257),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_111),
.A2(n_112),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g269 ( 
.A1(n_120),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_121),
.B(n_122),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_137),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_124),
.B(n_130),
.C(n_137),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_125),
.B(n_128),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_129),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_131),
.B(n_133),
.C(n_135),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_219),
.B(n_224),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_205),
.B(n_218),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_184),
.B(n_204),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_163),
.B(n_183),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_153),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_158),
.C(n_160),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_171),
.B(n_182),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_170),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_181),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_186),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_197),
.B1(n_202),
.B2(n_203),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_188),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_196),
.C(n_203),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_200),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_214),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_242),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_242),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.C(n_241),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_233),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_227),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.CI(n_232),
.CON(n_227),
.SN(n_227)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_229),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_239),
.B2(n_240),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_234),
.B(n_240),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_240),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_239),
.A2(n_255),
.B(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_261),
.B2(n_262),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_245),
.B(n_252),
.C(n_262),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_249),
.B(n_251),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_249),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_248),
.Y(n_282)
);

FAx1_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_276),
.CI(n_288),
.CON(n_275),
.SN(n_275)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_264),
.A2(n_269),
.B(n_272),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_289),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_275),
.B(n_302),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_289),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_287),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_278),
.B1(n_291),
.B2(n_299),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_281),
.C(n_286),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_299),
.C(n_300),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_284),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_286),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_292),
.C(n_296),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_300),
.Y(n_289)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_294),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_296),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_297),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_320),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_318),
.B2(n_319),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);


endmodule