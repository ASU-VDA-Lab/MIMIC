module fake_jpeg_28123_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_24),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_0),
.B(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_3),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_25),
.B1(n_17),
.B2(n_23),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_26),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_41),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_13),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_24),
.C(n_20),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.C(n_38),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_24),
.C(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_37),
.B1(n_38),
.B2(n_32),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_52),
.B1(n_54),
.B2(n_21),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_37),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_53),
.C(n_54),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_12),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_61),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_17),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_31),
.B1(n_15),
.B2(n_11),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_31),
.B1(n_11),
.B2(n_7),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_65),
.Y(n_67)
);

AOI221xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_65)
);

NAND4xp25_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_5),
.C(n_25),
.D(n_26),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_68),
.A2(n_64),
.B(n_66),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_67),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_70),
.Y(n_71)
);


endmodule