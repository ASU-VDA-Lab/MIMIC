module fake_jpeg_12502_n_531 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_531);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_57),
.B(n_93),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_76),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_18),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_79),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_90),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_27),
.C(n_40),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_36),
.C(n_43),
.Y(n_145)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_96),
.Y(n_108)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_28),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_20),
.B(n_17),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_20),
.B(n_17),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_97),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_100),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_25),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_39),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_20),
.B1(n_45),
.B2(n_44),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_112),
.A2(n_125),
.B1(n_19),
.B2(n_40),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_14),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_124),
.B(n_151),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_65),
.A2(n_25),
.B1(n_45),
.B2(n_44),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_66),
.B1(n_59),
.B2(n_62),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_38),
.B1(n_24),
.B2(n_29),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_36),
.B1(n_45),
.B2(n_44),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_130),
.A2(n_139),
.B1(n_147),
.B2(n_149),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_36),
.B1(n_43),
.B2(n_25),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_39),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_38),
.C(n_24),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_69),
.A2(n_26),
.B1(n_43),
.B2(n_30),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_76),
.A2(n_30),
.B1(n_26),
.B2(n_41),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_81),
.B(n_15),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_64),
.B(n_16),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_152),
.B(n_158),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_77),
.A2(n_26),
.B1(n_30),
.B2(n_41),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_160),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_79),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_101),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_53),
.B(n_14),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_54),
.B(n_16),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_161),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_96),
.A2(n_38),
.B1(n_29),
.B2(n_34),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_80),
.B(n_16),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_163),
.B(n_168),
.Y(n_229)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_100),
.B1(n_99),
.B2(n_74),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_165),
.A2(n_180),
.B1(n_185),
.B2(n_200),
.Y(n_250)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_85),
.B1(n_39),
.B2(n_41),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_167),
.A2(n_197),
.B1(n_148),
.B2(n_136),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_169),
.B(n_174),
.Y(n_222)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_172),
.A2(n_144),
.B(n_118),
.Y(n_259)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_101),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_40),
.B1(n_24),
.B2(n_29),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_108),
.A2(n_47),
.B(n_42),
.C(n_19),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_176),
.A2(n_115),
.B(n_117),
.C(n_131),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_178),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_179),
.B(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_183),
.B(n_190),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_105),
.B(n_82),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_108),
.A2(n_34),
.B1(n_19),
.B2(n_42),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_127),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_111),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_192),
.B(n_193),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_82),
.Y(n_193)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

BUFx2_ASAP7_75t_SL g255 ( 
.A(n_195),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_71),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_199),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_103),
.A2(n_34),
.B1(n_47),
.B2(n_3),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_113),
.B(n_71),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_135),
.A2(n_61),
.B1(n_47),
.B2(n_3),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_120),
.B(n_61),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_205),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_109),
.A2(n_47),
.B1(n_1),
.B2(n_3),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_207),
.B1(n_187),
.B2(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_109),
.B(n_0),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_117),
.B(n_1),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_127),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_106),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_214),
.B1(n_133),
.B2(n_141),
.Y(n_237)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_142),
.B(n_4),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_110),
.Y(n_217)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_146),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_113),
.B(n_5),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_6),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_110),
.B(n_13),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_220),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_221),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_223),
.B(n_227),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_243),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_148),
.B1(n_136),
.B2(n_133),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_235),
.A2(n_237),
.B1(n_247),
.B2(n_264),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_263),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_169),
.A2(n_114),
.B(n_115),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_176),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_188),
.A2(n_156),
.B1(n_129),
.B2(n_141),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_138),
.B(n_8),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_260),
.B(n_169),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_168),
.A2(n_194),
.B1(n_201),
.B2(n_184),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_214),
.A2(n_156),
.B1(n_129),
.B2(n_107),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_177),
.B(n_114),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_269),
.B(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_177),
.B(n_115),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_286),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_279),
.B(n_282),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_229),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_303),
.C(n_318),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_247),
.A2(n_165),
.B1(n_200),
.B2(n_179),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_281),
.A2(n_312),
.B1(n_316),
.B2(n_321),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_206),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_238),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_283),
.B(n_287),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_234),
.A2(n_190),
.B1(n_209),
.B2(n_218),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_250),
.A2(n_219),
.B1(n_194),
.B2(n_203),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_285),
.A2(n_297),
.B1(n_309),
.B2(n_224),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_220),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_189),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_288),
.B(n_289),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_232),
.B(n_215),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_220),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_296),
.Y(n_330)
);

OA22x2_ASAP7_75t_L g291 ( 
.A1(n_250),
.A2(n_176),
.B1(n_166),
.B2(n_170),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g357 ( 
.A1(n_291),
.A2(n_262),
.B(n_249),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_210),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_294),
.Y(n_351)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_234),
.A2(n_176),
.B1(n_213),
.B2(n_164),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_232),
.B(n_208),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_300),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_225),
.B(n_226),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_225),
.B(n_204),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_306),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_230),
.B(n_212),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_217),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_305),
.C(n_307),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_171),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_226),
.B(n_198),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_230),
.B(n_176),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_231),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_310),
.C(n_315),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_235),
.A2(n_191),
.B1(n_178),
.B2(n_118),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_231),
.B(n_107),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_223),
.A2(n_191),
.B1(n_178),
.B2(n_132),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_116),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_116),
.B1(n_144),
.B2(n_138),
.Y(n_316)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_255),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_138),
.C(n_7),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_319),
.A2(n_262),
.B(n_261),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_320),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_268),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_300),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_323),
.B(n_329),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_292),
.A2(n_259),
.B(n_227),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_324),
.A2(n_337),
.B(n_357),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_327),
.A2(n_331),
.B1(n_339),
.B2(n_342),
.Y(n_383)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_227),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_328),
.B(n_344),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_302),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_276),
.A2(n_270),
.B1(n_272),
.B2(n_228),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_239),
.B(n_241),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_276),
.A2(n_228),
.B1(n_251),
.B2(n_256),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_276),
.A2(n_251),
.B1(n_241),
.B2(n_254),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_277),
.Y(n_343)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_248),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_347),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_306),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_353),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_280),
.B(n_265),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_349),
.Y(n_375)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_295),
.Y(n_352)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_274),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_281),
.A2(n_239),
.B1(n_254),
.B2(n_233),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_354),
.A2(n_314),
.B1(n_309),
.B2(n_297),
.Y(n_365)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_249),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_290),
.B(n_265),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_358),
.A2(n_360),
.B(n_319),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_365),
.A2(n_378),
.B1(n_393),
.B2(n_359),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_327),
.A2(n_278),
.B1(n_292),
.B2(n_275),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_367),
.A2(n_384),
.B1(n_354),
.B2(n_348),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_298),
.C(n_292),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_372),
.C(n_376),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_350),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_379),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_338),
.B(n_289),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_370),
.B(n_374),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_285),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_326),
.B(n_279),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_303),
.C(n_307),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_328),
.A2(n_291),
.B1(n_278),
.B2(n_274),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_359),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_291),
.B1(n_318),
.B2(n_311),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_335),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_286),
.C(n_291),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_385),
.C(n_388),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_353),
.A2(n_312),
.B1(n_316),
.B2(n_310),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_311),
.C(n_293),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_363),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_391),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_321),
.Y(n_388)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_331),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_340),
.A2(n_320),
.B1(n_233),
.B2(n_271),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_360),
.A2(n_324),
.B(n_358),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_337),
.A2(n_357),
.B(n_359),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_395),
.A2(n_322),
.B(n_334),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_236),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_397),
.C(n_325),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_332),
.B(n_236),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_339),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_398),
.B(n_356),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_380),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_407),
.Y(n_441)
);

AO22x1_ASAP7_75t_SL g401 ( 
.A1(n_371),
.A2(n_357),
.B1(n_323),
.B2(n_329),
.Y(n_401)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_401),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_408),
.A2(n_416),
.B1(n_406),
.B2(n_365),
.Y(n_437)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_409),
.Y(n_443)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_361),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_413),
.A2(n_375),
.B1(n_388),
.B2(n_377),
.Y(n_434)
);

OAI32xp33_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_341),
.A3(n_351),
.B1(n_355),
.B2(n_347),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_423),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_367),
.A2(n_383),
.B1(n_384),
.B2(n_366),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_342),
.C(n_325),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_419),
.C(n_424),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_392),
.B(n_336),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_429),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_368),
.B(n_343),
.C(n_336),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_364),
.B(n_346),
.Y(n_420)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_372),
.B(n_345),
.Y(n_421)
);

XNOR2x1_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_382),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_334),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_422),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_333),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_373),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_389),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_333),
.C(n_352),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_427),
.B(n_385),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_397),
.B(n_322),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_451),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_414),
.Y(n_431)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_454),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_434),
.A2(n_436),
.B1(n_452),
.B2(n_453),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_409),
.A2(n_377),
.B1(n_378),
.B2(n_371),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_437),
.A2(n_445),
.B1(n_446),
.B2(n_402),
.Y(n_459)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_387),
.Y(n_442)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_416),
.A2(n_395),
.B1(n_393),
.B2(n_377),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_408),
.A2(n_394),
.B1(n_381),
.B2(n_374),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_399),
.Y(n_450)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_450),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_399),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_419),
.B(n_261),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_233),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_242),
.Y(n_455)
);

INVx11_ASAP7_75t_L g456 ( 
.A(n_455),
.Y(n_456)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_458),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_459),
.A2(n_470),
.B1(n_472),
.B2(n_436),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_405),
.C(n_410),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_463),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_435),
.A2(n_428),
.B(n_402),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_410),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_471),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_405),
.C(n_417),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_466),
.B(n_473),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_428),
.B(n_423),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_474),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_437),
.A2(n_403),
.B1(n_401),
.B2(n_426),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_421),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_445),
.A2(n_443),
.B1(n_448),
.B2(n_449),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_415),
.C(n_401),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_443),
.A2(n_415),
.B1(n_422),
.B2(n_361),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_317),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_440),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_479),
.A2(n_473),
.B1(n_456),
.B2(n_476),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_460),
.C(n_466),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_480),
.B(n_483),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_468),
.B(n_441),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_463),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_448),
.C(n_449),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_485),
.B(n_486),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_432),
.C(n_447),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_475),
.Y(n_487)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_487),
.Y(n_504)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_8),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_SL g489 ( 
.A(n_456),
.B(n_439),
.C(n_442),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_489),
.A2(n_474),
.B(n_471),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_432),
.C(n_447),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_491),
.C(n_485),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_438),
.C(n_439),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_490),
.A2(n_462),
.B1(n_472),
.B2(n_470),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_494),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_491),
.A2(n_469),
.B1(n_464),
.B2(n_467),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_495),
.B(n_497),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_500),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_499),
.A2(n_501),
.B(n_506),
.Y(n_510)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_481),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_492),
.A2(n_320),
.B(n_317),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_486),
.A2(n_242),
.B1(n_271),
.B2(n_9),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_503),
.C(n_10),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_6),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_480),
.C(n_478),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_508),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_496),
.A2(n_481),
.B(n_482),
.Y(n_511)
);

OAI211xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_513),
.B(n_514),
.C(n_504),
.Y(n_521)
);

NOR2x1_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_498),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_512),
.A2(n_505),
.B(n_502),
.Y(n_519)
);

NAND2x1_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_10),
.Y(n_513)
);

O2A1O1Ixp33_ASAP7_75t_SL g514 ( 
.A1(n_493),
.A2(n_10),
.B(n_11),
.C(n_500),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_501),
.C(n_503),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_506),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_517),
.A2(n_519),
.B(n_522),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_521),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_509),
.C(n_507),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_520),
.B(n_514),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_526),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_507),
.C(n_510),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_523),
.A2(n_525),
.B(n_512),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_528),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_527),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_530),
.Y(n_531)
);


endmodule