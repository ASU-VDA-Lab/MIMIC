module real_jpeg_14347_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_45),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_45),
.B1(n_62),
.B2(n_63),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_71),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_65),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_11),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_12),
.B(n_135),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_99),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_63),
.C(n_82),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_12),
.B(n_35),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_12),
.A2(n_66),
.B(n_163),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_27),
.B(n_34),
.C(n_190),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_99),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_13),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_79),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_79),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_15),
.A2(n_29),
.B1(n_43),
.B2(n_44),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_15),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_197)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_121),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_87),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_21),
.A2(n_22),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_41),
.B2(n_54),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_54),
.C(n_55),
.Y(n_120)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_26),
.A2(n_30),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_44),
.A3(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_30),
.A2(n_38),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_31),
.B(n_39),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_33),
.A2(n_36),
.B(n_99),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_36),
.A2(n_37),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_37),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_48),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_44),
.A2(n_50),
.B(n_99),
.C(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_46),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_61),
.A2(n_66),
.B1(n_72),
.B2(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_68),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_63),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_62),
.B(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_72),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_66),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_67),
.A2(n_68),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_67),
.B(n_164),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_68),
.B(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_72),
.A2(n_169),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_72),
.B(n_99),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_72),
.A2(n_137),
.B(n_177),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_73),
.B(n_87),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_77),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_85),
.B1(n_86),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_80),
.A2(n_86),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_84),
.A2(n_90),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_84),
.B(n_99),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_91),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.C(n_95),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_92),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_94),
.B(n_118),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_96),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_120),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_119),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_141),
.B(n_221),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_138),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_125),
.B(n_138),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_131),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_129),
.B(n_131),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.C(n_136),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_132),
.B(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_136),
.Y(n_207)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_216),
.B(n_220),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_201),
.B(n_215),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_185),
.B(n_200),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_165),
.B(n_184),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_154),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_148),
.B1(n_152),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B(n_151),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_149),
.A2(n_151),
.B(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_162),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_173),
.B(n_183),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_171),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_178),
.B(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_187),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_195),
.C(n_199),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_191),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_192)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_203),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_211),
.C(n_213),
.Y(n_217)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);


endmodule