module fake_netlist_6_1571_n_2662 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2662);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2662;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1674;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_2247;
wire n_544;
wire n_1711;
wire n_1078;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_2356;
wire n_1143;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_2480;
wire n_641;
wire n_1300;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_405;
wire n_2660;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_659;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1967;
wire n_1193;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_423;
wire n_1865;
wire n_586;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_595;
wire n_1767;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1627;
wire n_1295;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_1932;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_1714;
wire n_872;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_1817;
wire n_926;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_526;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_2482;
wire n_1507;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1475;
wire n_1774;
wire n_716;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_2354;
wire n_623;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1837;
wire n_600;
wire n_964;
wire n_831;
wire n_2218;
wire n_1314;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2617;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_1243;
wire n_848;
wire n_2249;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_2049;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1818;
wire n_1108;
wire n_710;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_411;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_1548;
wire n_799;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_786;
wire n_706;
wire n_1962;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_1476;
wire n_841;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_601;
wire n_2385;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1848;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_2584;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_1303;
wire n_761;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_611;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_2265;
wire n_2615;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_771;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_455;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_2600;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_629;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g391 ( 
.A(n_91),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_271),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_47),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_386),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_210),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_97),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_109),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_185),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_108),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_148),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_311),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_336),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_385),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_81),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_314),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_306),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_99),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_359),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_349),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_44),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_275),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_61),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_252),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_388),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_310),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_347),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_213),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_65),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_380),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_325),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_254),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_116),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_17),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_363),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_250),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_265),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_59),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_52),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_277),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_202),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_227),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_149),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_362),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_16),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_115),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_211),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_291),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_366),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_286),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_269),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_186),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_103),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_315),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_203),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_215),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_338),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_323),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_46),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_263),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_116),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_320),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_117),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_80),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_272),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_305),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_160),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_337),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_14),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_185),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_276),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_30),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_110),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_318),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_236),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_260),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_15),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_356),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_117),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_295),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_54),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_208),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_375),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_346),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_361),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_378),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_21),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_285),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_226),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_274),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_91),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_47),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_112),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_74),
.Y(n_487)
);

BUFx8_ASAP7_75t_SL g488 ( 
.A(n_296),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_298),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_327),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_78),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_280),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_57),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_308),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_220),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_141),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_82),
.Y(n_497)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_371),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_183),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_367),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_17),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_351),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_201),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_243),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_256),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_11),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_230),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_130),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_281),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_167),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_107),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_340),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_189),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_379),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_129),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_121),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_283),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_382),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_244),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_194),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_234),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_114),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_68),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_390),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_360),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_99),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_301),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_9),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_258),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_15),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_241),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_144),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_16),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_36),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_261),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_64),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_245),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_52),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_118),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_259),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_174),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_309),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_365),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_150),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_83),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_247),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_307),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_164),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_249),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_9),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_8),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_144),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_206),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_339),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_300),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_209),
.Y(n_556)
);

BUFx8_ASAP7_75t_SL g557 ( 
.A(n_2),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_255),
.Y(n_558)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_289),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_358),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_389),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_313),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_264),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_205),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_33),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_342),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_278),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_173),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_82),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_60),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_139),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_67),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_34),
.Y(n_573)
);

BUFx2_ASAP7_75t_SL g574 ( 
.A(n_63),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_335),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_332),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_302),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_328),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_130),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_98),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_221),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_352),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_344),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g584 ( 
.A(n_329),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_84),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_303),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_13),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_292),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_293),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_288),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_187),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_290),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_181),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_376),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_357),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_355),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_18),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_228),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_69),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_88),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_372),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_354),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_19),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_108),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_229),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_13),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_37),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_373),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_95),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_297),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_138),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_92),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_88),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_24),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_121),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_240),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_4),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_173),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_167),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_237),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_319),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_65),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_317),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_137),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_90),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_178),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_345),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_8),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_174),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_50),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_114),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_40),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_147),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_381),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_191),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_216),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_268),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_370),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_324),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_75),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_58),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_199),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_22),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_246),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_383),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_219),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_63),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_248),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_106),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_77),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_267),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_175),
.Y(n_652)
);

CKINVDCx16_ASAP7_75t_R g653 ( 
.A(n_44),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_109),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_284),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_176),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_304),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_178),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_166),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_55),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_28),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_331),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_146),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_74),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_96),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_175),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_0),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_235),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_49),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_80),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_36),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_153),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_132),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_225),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_170),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_104),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_364),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_200),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_334),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_101),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_282),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_0),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_113),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_348),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_333),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_26),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_122),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_377),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_262),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_198),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_165),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_122),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_96),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_270),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_322),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_12),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_128),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_341),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_163),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_35),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_257),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_299),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_330),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_326),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_92),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_31),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_28),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_66),
.Y(n_708)
);

INVxp33_ASAP7_75t_SL g709 ( 
.A(n_172),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_7),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_55),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_343),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_369),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_86),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_78),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_62),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_39),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_29),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_45),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_176),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_168),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_137),
.Y(n_722)
);

BUFx8_ASAP7_75t_SL g723 ( 
.A(n_294),
.Y(n_723)
);

INVxp33_ASAP7_75t_L g724 ( 
.A(n_113),
.Y(n_724)
);

BUFx8_ASAP7_75t_SL g725 ( 
.A(n_196),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_242),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_56),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_87),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_312),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_287),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_163),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_279),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_207),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_316),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_73),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_93),
.Y(n_736)
);

BUFx8_ASAP7_75t_SL g737 ( 
.A(n_66),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_35),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_273),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_266),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_41),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_10),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_368),
.Y(n_743)
);

CKINVDCx16_ASAP7_75t_R g744 ( 
.A(n_253),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_251),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_321),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_353),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_129),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_104),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_391),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_391),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_557),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_442),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_569),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_569),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_442),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_737),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_572),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_572),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_579),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_579),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_666),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_622),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_442),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_455),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_622),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_480),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_671),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_642),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_664),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_671),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_442),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_442),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_528),
.Y(n_774)
);

CKINVDCx14_ASAP7_75t_R g775 ( 
.A(n_498),
.Y(n_775)
);

BUFx5_ASAP7_75t_L g776 ( 
.A(n_406),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_440),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_528),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_528),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_745),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_528),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_528),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_412),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_488),
.Y(n_784)
);

INVxp33_ASAP7_75t_L g785 ( 
.A(n_714),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_585),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_585),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_418),
.Y(n_788)
);

CKINVDCx14_ASAP7_75t_R g789 ( 
.A(n_559),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_451),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_585),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_585),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_585),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_735),
.Y(n_794)
);

CKINVDCx16_ASAP7_75t_R g795 ( 
.A(n_653),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_480),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_735),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_482),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_480),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_735),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_735),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_735),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_742),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_742),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_742),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_742),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_626),
.Y(n_807)
);

INVxp33_ASAP7_75t_L g808 ( 
.A(n_724),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_742),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_626),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_434),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_459),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_461),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_485),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_626),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_396),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_464),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_399),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_404),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_493),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_497),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_396),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_469),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_499),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_399),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_501),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_523),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_532),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_534),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_544),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_597),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_609),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_423),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_570),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_573),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_554),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_614),
.Y(n_837)
);

INVxp33_ASAP7_75t_L g838 ( 
.A(n_465),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_628),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_640),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_643),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_649),
.Y(n_842)
);

CKINVDCx14_ASAP7_75t_R g843 ( 
.A(n_584),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_440),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_654),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_723),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_665),
.Y(n_847)
);

INVxp33_ASAP7_75t_SL g848 ( 
.A(n_397),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_667),
.Y(n_849)
);

INVxp33_ASAP7_75t_SL g850 ( 
.A(n_397),
.Y(n_850)
);

INVxp33_ASAP7_75t_L g851 ( 
.A(n_465),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_473),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_669),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_680),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_682),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_725),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_683),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_687),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_398),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_692),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_693),
.Y(n_861)
);

CKINVDCx14_ASAP7_75t_R g862 ( 
.A(n_467),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_705),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_707),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_744),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_708),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_719),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_722),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_727),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_600),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_502),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_484),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_486),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_619),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_487),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_686),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_625),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_502),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_421),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_425),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_668),
.Y(n_882)
);

CKINVDCx16_ASAP7_75t_R g883 ( 
.A(n_686),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_436),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_446),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_473),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_398),
.Y(n_887)
);

INVxp33_ASAP7_75t_L g888 ( 
.A(n_496),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_400),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_496),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_491),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_450),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_452),
.Y(n_893)
);

INVxp33_ASAP7_75t_L g894 ( 
.A(n_548),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_548),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_457),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_458),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_474),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_467),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_476),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_633),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_552),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_494),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_506),
.Y(n_904)
);

INVxp33_ASAP7_75t_L g905 ( 
.A(n_552),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_503),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_512),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_514),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_519),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_466),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_525),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_537),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_540),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_618),
.Y(n_914)
);

INVxp33_ASAP7_75t_SL g915 ( 
.A(n_400),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_543),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_686),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_553),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_508),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_661),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_558),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_691),
.Y(n_922)
);

CKINVDCx16_ASAP7_75t_R g923 ( 
.A(n_413),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_563),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_577),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_578),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_590),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_594),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_595),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_411),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_574),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_467),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_510),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_407),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_407),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_618),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_637),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_638),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_645),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_511),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_651),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_679),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_410),
.Y(n_943)
);

INVxp33_ASAP7_75t_SL g944 ( 
.A(n_410),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_685),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_690),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_411),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_422),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_422),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_695),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_663),
.Y(n_951)
);

CKINVDCx14_ASAP7_75t_R g952 ( 
.A(n_621),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_701),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_712),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_729),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_515),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_431),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_427),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_663),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_431),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_507),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_621),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_639),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_507),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_621),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_509),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_509),
.Y(n_967)
);

CKINVDCx16_ASAP7_75t_R g968 ( 
.A(n_444),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_468),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_549),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_470),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_549),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_646),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_427),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_646),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_684),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_684),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_747),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_747),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_430),
.Y(n_980)
);

CKINVDCx14_ASAP7_75t_R g981 ( 
.A(n_704),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_430),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_445),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_704),
.Y(n_984)
);

INVxp67_ASAP7_75t_SL g985 ( 
.A(n_749),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_428),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_445),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_542),
.Y(n_988)
);

BUFx5_ASAP7_75t_L g989 ( 
.A(n_704),
.Y(n_989)
);

INVxp67_ASAP7_75t_SL g990 ( 
.A(n_612),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_542),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_428),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_576),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_639),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_748),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_576),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_583),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_583),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_702),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_702),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_734),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_734),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_603),
.B(n_1),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_603),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_639),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_516),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_522),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_526),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_432),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_530),
.Y(n_1010)
);

BUFx2_ASAP7_75t_SL g1011 ( 
.A(n_447),
.Y(n_1011)
);

CKINVDCx14_ASAP7_75t_R g1012 ( 
.A(n_392),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_533),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_432),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_536),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_435),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_435),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_538),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_539),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_639),
.Y(n_1020)
);

INVxp33_ASAP7_75t_SL g1021 ( 
.A(n_443),
.Y(n_1021)
);

CKINVDCx14_ASAP7_75t_R g1022 ( 
.A(n_392),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_541),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_545),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_550),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_551),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_565),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_394),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_568),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_393),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_571),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_639),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_580),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_587),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_591),
.Y(n_1035)
);

NOR2xp67_ASAP7_75t_L g1036 ( 
.A(n_593),
.B(n_1),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_472),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_599),
.Y(n_1038)
);

AND2x6_ASAP7_75t_L g1039 ( 
.A(n_963),
.B(n_402),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_997),
.B(n_709),
.Y(n_1040)
);

INVx5_ASAP7_75t_L g1041 ( 
.A(n_879),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_757),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1037),
.B(n_477),
.Y(n_1043)
);

BUFx8_ASAP7_75t_SL g1044 ( 
.A(n_752),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1028),
.B(n_456),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_753),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_808),
.B(n_475),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_808),
.B(n_564),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_1037),
.B(n_394),
.Y(n_1049)
);

AND2x6_ASAP7_75t_L g1050 ( 
.A(n_963),
.B(n_471),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_1028),
.B(n_395),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_775),
.B(n_395),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_910),
.B(n_478),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_757),
.Y(n_1054)
);

INVx5_ASAP7_75t_L g1055 ( 
.A(n_879),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_784),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_777),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_753),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_756),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_756),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_969),
.B(n_401),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_764),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_899),
.B(n_401),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_846),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_971),
.B(n_403),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_879),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_899),
.B(n_403),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_836),
.B(n_405),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_1012),
.B(n_405),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_764),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_989),
.B(n_479),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_930),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_772),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_772),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_800),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_800),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1030),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_930),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_777),
.Y(n_1079)
);

INVx6_ASAP7_75t_L g1080 ( 
.A(n_932),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_775),
.B(n_408),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_994),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_932),
.B(n_408),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1012),
.B(n_409),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_962),
.B(n_505),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_788),
.B(n_409),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_789),
.B(n_843),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_962),
.B(n_414),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_773),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_989),
.B(n_481),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_984),
.B(n_414),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_789),
.B(n_843),
.Y(n_1092)
);

BUFx12f_ASAP7_75t_L g1093 ( 
.A(n_856),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_783),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_984),
.B(n_415),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_930),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_989),
.B(n_844),
.Y(n_1097)
);

INVx5_ASAP7_75t_L g1098 ( 
.A(n_947),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_994),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1005),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_862),
.B(n_415),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_817),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_1032),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_SL g1104 ( 
.A(n_798),
.B(n_521),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1032),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_774),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_778),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_779),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1022),
.B(n_416),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_781),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_782),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1022),
.B(n_416),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_788),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_786),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_871),
.B(n_417),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1006),
.B(n_417),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1011),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_790),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_989),
.B(n_483),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1007),
.B(n_419),
.Y(n_1120)
);

INVx5_ASAP7_75t_L g1121 ( 
.A(n_947),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_947),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_989),
.B(n_489),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_989),
.B(n_490),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_989),
.B(n_1008),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_790),
.B(n_419),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_787),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_817),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1010),
.B(n_492),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_823),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_823),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_873),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_965),
.B(n_769),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_873),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_791),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_792),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_793),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_934),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_862),
.B(n_420),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1013),
.B(n_420),
.Y(n_1140)
);

AND2x6_ASAP7_75t_L g1141 ( 
.A(n_957),
.B(n_604),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_794),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_952),
.B(n_424),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_865),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_780),
.B(n_424),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_767),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_797),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1018),
.B(n_495),
.Y(n_1148)
);

INVx5_ASAP7_75t_L g1149 ( 
.A(n_807),
.Y(n_1149)
);

BUFx8_ASAP7_75t_L g1150 ( 
.A(n_859),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_874),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_801),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_882),
.B(n_426),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1019),
.B(n_500),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_802),
.Y(n_1155)
);

INVx5_ASAP7_75t_L g1156 ( 
.A(n_815),
.Y(n_1156)
);

CKINVDCx6p67_ASAP7_75t_R g1157 ( 
.A(n_752),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_934),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1023),
.B(n_504),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_931),
.B(n_426),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_803),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_804),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1024),
.B(n_513),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1025),
.B(n_429),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1027),
.B(n_1029),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1031),
.B(n_517),
.Y(n_1166)
);

BUFx8_ASAP7_75t_SL g1167 ( 
.A(n_819),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_874),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_876),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_876),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1033),
.B(n_1034),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_891),
.B(n_429),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_805),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_877),
.B(n_443),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_806),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_809),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1038),
.B(n_518),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_985),
.B(n_433),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_891),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_952),
.B(n_433),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_904),
.B(n_919),
.Y(n_1181)
);

INVx6_ASAP7_75t_L g1182 ( 
.A(n_883),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_818),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_818),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_990),
.B(n_437),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_825),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_884),
.B(n_520),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_904),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_935),
.B(n_986),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_995),
.B(n_1017),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_919),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_933),
.B(n_437),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_825),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_896),
.B(n_908),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_852),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_852),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_886),
.Y(n_1197)
);

AND2x6_ASAP7_75t_L g1198 ( 
.A(n_960),
.B(n_617),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_981),
.B(n_438),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_933),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_940),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_886),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_981),
.B(n_438),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_890),
.Y(n_1204)
);

BUFx8_ASAP7_75t_SL g1205 ( 
.A(n_819),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_890),
.Y(n_1206)
);

INVx5_ASAP7_75t_L g1207 ( 
.A(n_895),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_816),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_895),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_911),
.B(n_439),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_902),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_940),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_902),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_943),
.Y(n_1214)
);

INVx6_ASAP7_75t_L g1215 ( 
.A(n_917),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_928),
.B(n_524),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_914),
.Y(n_1217)
);

INVx5_ASAP7_75t_L g1218 ( 
.A(n_914),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_942),
.B(n_1020),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_776),
.B(n_527),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_770),
.B(n_750),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_956),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1079),
.B(n_936),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1079),
.B(n_1057),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1097),
.B(n_1125),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1106),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1077),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1082),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1059),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1059),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1082),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1041),
.B(n_936),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1047),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1220),
.A2(n_964),
.B(n_961),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1048),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1106),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1062),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1062),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_1117),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1106),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1082),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1049),
.B(n_1043),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1179),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1219),
.B(n_776),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1108),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1146),
.B(n_765),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1099),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1127),
.A2(n_967),
.B(n_966),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1108),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1108),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1146),
.B(n_956),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1075),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1114),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1041),
.B(n_1055),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1094),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1114),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1099),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1189),
.A2(n_1026),
.B1(n_1035),
.B2(n_1015),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1114),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1146),
.B(n_1015),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1099),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1135),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1041),
.B(n_951),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1135),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1135),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1040),
.A2(n_850),
.B1(n_915),
.B2(n_848),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1137),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1137),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1153),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1046),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1149),
.B(n_1026),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1075),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1149),
.B(n_1035),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1137),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1127),
.A2(n_972),
.B(n_970),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1155),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1149),
.B(n_785),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1055),
.B(n_951),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1076),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1055),
.B(n_959),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1066),
.B(n_776),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1155),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1046),
.Y(n_1283)
);

OA21x2_ASAP7_75t_L g1284 ( 
.A1(n_1136),
.A2(n_975),
.B(n_973),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1046),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1066),
.B(n_776),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1066),
.B(n_776),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1115),
.B(n_959),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1156),
.B(n_1101),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1187),
.B(n_776),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1076),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1216),
.B(n_776),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1184),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1115),
.B(n_980),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1155),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1129),
.B(n_1148),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1051),
.B(n_982),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1184),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1161),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1161),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1154),
.B(n_880),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1159),
.B(n_881),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1163),
.B(n_885),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1162),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1166),
.B(n_892),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1100),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1162),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1058),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1184),
.Y(n_1310)
);

BUFx8_ASAP7_75t_L g1311 ( 
.A(n_1138),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1195),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1177),
.B(n_1061),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1162),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1195),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1189),
.A2(n_848),
.B1(n_915),
.B2(n_850),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1195),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1058),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1145),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1196),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1136),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1196),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1100),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1156),
.B(n_785),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1142),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1142),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1051),
.B(n_983),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1190),
.A2(n_944),
.B1(n_1021),
.B2(n_795),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1196),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1065),
.B(n_893),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1173),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1190),
.A2(n_1021),
.B1(n_944),
.B2(n_556),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1167),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1173),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1116),
.B(n_987),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1165),
.B(n_887),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1206),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1160),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1176),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1176),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1089),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1206),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1107),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1110),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1156),
.B(n_949),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1058),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1222),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1111),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1206),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1103),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1147),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1152),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1209),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1060),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1175),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1209),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1209),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1063),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1071),
.A2(n_977),
.B(n_976),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1213),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1213),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1103),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1213),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1139),
.B(n_958),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1217),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1103),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1205),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1116),
.B(n_988),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1217),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1217),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1105),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1171),
.B(n_897),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1060),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1060),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1063),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1105),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1128),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1070),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1174),
.A2(n_992),
.B1(n_1009),
.B2(n_943),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1105),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1143),
.B(n_822),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1045),
.B(n_529),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1227),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1227),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1228),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1223),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1297),
.B(n_1045),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1233),
.B(n_1133),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1223),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1223),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1321),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1233),
.B(n_1178),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1325),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1229),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1229),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1230),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1230),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1326),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1331),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1334),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1248),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1228),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1235),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1339),
.Y(n_1404)
);

XNOR2xp5_ASAP7_75t_L g1405 ( 
.A(n_1333),
.B(n_833),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1358),
.B(n_1132),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1237),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1237),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1224),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1238),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1238),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1252),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1252),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1242),
.B(n_1130),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1340),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1225),
.A2(n_1039),
.B1(n_1050),
.B2(n_1120),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1338),
.B(n_1181),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1246),
.B(n_1178),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1336),
.B(n_1185),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1313),
.B(n_1090),
.Y(n_1420)
);

INVx5_ASAP7_75t_L g1421 ( 
.A(n_1228),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1288),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1272),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1239),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1244),
.B(n_1130),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1338),
.B(n_1119),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1288),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1288),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1224),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1272),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1279),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1279),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1228),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1269),
.B(n_1172),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1269),
.B(n_1290),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1291),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1231),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1292),
.B(n_1131),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1291),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1319),
.B(n_1131),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1336),
.B(n_1068),
.C(n_1192),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_SL g1442 ( 
.A(n_1330),
.B(n_547),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1248),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1248),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1302),
.B(n_1124),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1231),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1224),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1277),
.B(n_1185),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1275),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1341),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1294),
.B(n_1120),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1319),
.B(n_1169),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1239),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1231),
.Y(n_1454)
);

BUFx10_ASAP7_75t_L g1455 ( 
.A(n_1377),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1298),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1377),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1303),
.B(n_1169),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1275),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1343),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1344),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1284),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1348),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1367),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1284),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1284),
.Y(n_1466)
);

BUFx8_ASAP7_75t_SL g1467 ( 
.A(n_1243),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1304),
.B(n_1188),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1351),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1293),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1293),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1299),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1381),
.B(n_1084),
.C(n_1069),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1306),
.B(n_1123),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1352),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1355),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1372),
.B(n_1194),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1299),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1294),
.A2(n_1140),
.B1(n_1164),
.B2(n_1104),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1310),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1231),
.Y(n_1481)
);

NOR2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1251),
.B(n_1113),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1310),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1312),
.Y(n_1484)
);

INVxp33_ASAP7_75t_SL g1485 ( 
.A(n_1379),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1364),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1312),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1315),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1315),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1241),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1294),
.B(n_1210),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1317),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1317),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1359),
.A2(n_1382),
.B(n_1378),
.Y(n_1494)
);

NAND2xp33_ASAP7_75t_SL g1495 ( 
.A(n_1382),
.B(n_1375),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1266),
.B(n_1188),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_L g1497 ( 
.A(n_1320),
.B(n_1039),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1322),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1322),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1298),
.B(n_1102),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1329),
.B(n_1210),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1329),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1337),
.Y(n_1503)
);

BUFx10_ASAP7_75t_L g1504 ( 
.A(n_1298),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1327),
.B(n_1085),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1241),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1337),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1324),
.B(n_1180),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1342),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1342),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1349),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1327),
.B(n_1053),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1255),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1327),
.B(n_1144),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1255),
.Y(n_1515)
);

AOI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1281),
.A2(n_1287),
.B(n_1286),
.Y(n_1516)
);

NAND2xp33_ASAP7_75t_L g1517 ( 
.A(n_1349),
.B(n_1039),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1353),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1335),
.B(n_1144),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1353),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1356),
.B(n_1109),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1241),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1356),
.Y(n_1523)
);

BUFx10_ASAP7_75t_L g1524 ( 
.A(n_1335),
.Y(n_1524)
);

AND2x6_ASAP7_75t_L g1525 ( 
.A(n_1289),
.B(n_1087),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1380),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1369),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1369),
.B(n_1112),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1335),
.B(n_1144),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1311),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1234),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1258),
.B(n_1134),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1368),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1232),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1234),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1368),
.B(n_1140),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1386),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1389),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1390),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1467),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1420),
.A2(n_1234),
.B(n_1359),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1422),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1427),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1428),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1419),
.B(n_1345),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1513),
.B(n_875),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1394),
.Y(n_1547)
);

AND2x6_ASAP7_75t_L g1548 ( 
.A(n_1531),
.B(n_1368),
.Y(n_1548)
);

AOI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1435),
.A2(n_1373),
.B(n_1370),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1394),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1467),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1486),
.B(n_1347),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1395),
.Y(n_1553)
);

XOR2xp5_ASAP7_75t_L g1554 ( 
.A(n_1405),
.B(n_833),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1383),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1388),
.B(n_1260),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1395),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1396),
.Y(n_1558)
);

AOI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1435),
.A2(n_1360),
.B(n_1357),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1396),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1477),
.B(n_1316),
.Y(n_1561)
);

XOR2xp5_ASAP7_75t_L g1562 ( 
.A(n_1424),
.B(n_834),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1464),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1384),
.B(n_923),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1397),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1397),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_R g1567 ( 
.A(n_1403),
.B(n_1158),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1445),
.B(n_1039),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1407),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1407),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1408),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1531),
.A2(n_1208),
.B(n_1332),
.Y(n_1572)
);

XNOR2xp5_ASAP7_75t_L g1573 ( 
.A(n_1464),
.B(n_834),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1417),
.B(n_1271),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1408),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1410),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1410),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1434),
.B(n_968),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1411),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1473),
.B(n_1056),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_R g1581 ( 
.A(n_1532),
.B(n_1214),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1441),
.B(n_835),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1496),
.B(n_1151),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1456),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_R g1585 ( 
.A(n_1485),
.B(n_1067),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1411),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1412),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1412),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1413),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_SL g1590 ( 
.A(n_1524),
.B(n_1168),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1392),
.B(n_1418),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1387),
.B(n_835),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1413),
.Y(n_1593)
);

XNOR2xp5_ASAP7_75t_L g1594 ( 
.A(n_1424),
.B(n_870),
.Y(n_1594)
);

XOR2xp5_ASAP7_75t_L g1595 ( 
.A(n_1453),
.B(n_870),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1402),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1423),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1423),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1524),
.B(n_1170),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1432),
.Y(n_1600)
);

INVxp33_ASAP7_75t_L g1601 ( 
.A(n_1387),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1432),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1515),
.B(n_1273),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1426),
.B(n_878),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1448),
.B(n_1191),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1430),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1431),
.Y(n_1607)
);

AND2x2_ASAP7_75t_SL g1608 ( 
.A(n_1530),
.B(n_1328),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1491),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1436),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1439),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1456),
.Y(n_1612)
);

NOR2xp67_ASAP7_75t_L g1613 ( 
.A(n_1453),
.B(n_1064),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1406),
.B(n_1536),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1533),
.Y(n_1615)
);

XNOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1482),
.B(n_1174),
.Y(n_1616)
);

XNOR2xp5_ASAP7_75t_L g1617 ( 
.A(n_1479),
.B(n_878),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1451),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1414),
.B(n_901),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1455),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1508),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1414),
.B(n_1067),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1470),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1534),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1474),
.B(n_1050),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1391),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_SL g1627 ( 
.A(n_1524),
.B(n_1212),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1393),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1401),
.B(n_1444),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1398),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1409),
.B(n_1164),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1399),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1440),
.B(n_901),
.Y(n_1633)
);

INVxp33_ASAP7_75t_SL g1634 ( 
.A(n_1440),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1535),
.A2(n_1363),
.B(n_1361),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1400),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1404),
.Y(n_1637)
);

NAND2x1p5_ASAP7_75t_L g1638 ( 
.A(n_1533),
.B(n_1261),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1415),
.Y(n_1639)
);

BUFx8_ASAP7_75t_L g1640 ( 
.A(n_1536),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1452),
.B(n_920),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1401),
.B(n_1050),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1455),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1470),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1402),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1452),
.B(n_1200),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1471),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1471),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1472),
.Y(n_1649)
);

INVxp33_ASAP7_75t_L g1650 ( 
.A(n_1500),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1472),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1478),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1478),
.Y(n_1653)
);

CKINVDCx14_ASAP7_75t_R g1654 ( 
.A(n_1455),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1483),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1483),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1626),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1604),
.B(n_1458),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1557),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1574),
.B(n_1521),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1628),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1561),
.B(n_1578),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1634),
.B(n_1451),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1629),
.A2(n_1421),
.B(n_1385),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1556),
.B(n_1528),
.Y(n_1665)
);

OR2x6_ASAP7_75t_L g1666 ( 
.A(n_1614),
.B(n_1406),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1621),
.B(n_1451),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1555),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1609),
.B(n_1458),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1609),
.B(n_1468),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1621),
.B(n_1468),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1545),
.B(n_1512),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1591),
.B(n_1512),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1584),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1625),
.B(n_1568),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1601),
.B(n_1201),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1625),
.B(n_1416),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1552),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1630),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1568),
.B(n_1501),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1584),
.B(n_1536),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1560),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1650),
.B(n_1505),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1546),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1576),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1584),
.B(n_1504),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1632),
.B(n_1447),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1582),
.B(n_1485),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1636),
.B(n_1409),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1612),
.B(n_1615),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1637),
.B(n_1429),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1592),
.A2(n_1495),
.B1(n_1442),
.B2(n_1505),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1640),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1605),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1639),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1548),
.A2(n_1442),
.B1(n_1495),
.B2(n_1141),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1548),
.A2(n_1141),
.B1(n_1198),
.B2(n_1050),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1548),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1542),
.B(n_1429),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1619),
.A2(n_1500),
.B1(n_1525),
.B2(n_1425),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1612),
.B(n_1504),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1543),
.B(n_1425),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1544),
.B(n_1438),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1602),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1548),
.A2(n_1198),
.B1(n_1141),
.B2(n_1497),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1567),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1633),
.A2(n_1525),
.B1(n_1514),
.B2(n_1519),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1547),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1537),
.B(n_1438),
.Y(n_1709)
);

OR2x2_ASAP7_75t_SL g1710 ( 
.A(n_1646),
.B(n_1182),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1550),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1603),
.B(n_1221),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1538),
.B(n_1525),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1553),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1641),
.A2(n_1525),
.B1(n_1514),
.B2(n_1519),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1558),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1563),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1539),
.B(n_1525),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1572),
.A2(n_762),
.B1(n_948),
.B2(n_974),
.C(n_889),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1572),
.A2(n_1198),
.B1(n_1141),
.B2(n_1497),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1624),
.B(n_1450),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1631),
.A2(n_1529),
.B1(n_1517),
.B2(n_1460),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1565),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1612),
.B(n_1615),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1631),
.A2(n_1529),
.B1(n_1517),
.B2(n_1461),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1606),
.B(n_1463),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1564),
.B(n_1469),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1680),
.A2(n_1421),
.B(n_1675),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1660),
.B(n_1662),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1662),
.B(n_1617),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1702),
.A2(n_1421),
.B(n_1541),
.Y(n_1732)
);

A2O1A1Ixp33_ASAP7_75t_L g1733 ( 
.A1(n_1658),
.A2(n_1622),
.B(n_1583),
.C(n_1580),
.Y(n_1733)
);

BUFx4f_ASAP7_75t_L g1734 ( 
.A(n_1674),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1688),
.B(n_1583),
.Y(n_1735)
);

CKINVDCx6p67_ASAP7_75t_R g1736 ( 
.A(n_1693),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1703),
.A2(n_1421),
.B(n_1541),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1665),
.B(n_1615),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1688),
.B(n_920),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1658),
.B(n_1590),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1677),
.A2(n_1642),
.B(n_1635),
.Y(n_1741)
);

INVx8_ASAP7_75t_L g1742 ( 
.A(n_1674),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1671),
.B(n_1618),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1709),
.A2(n_1437),
.B(n_1385),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1674),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1672),
.A2(n_1437),
.B(n_1385),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1669),
.B(n_1613),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1676),
.B(n_1590),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1676),
.B(n_1678),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1670),
.A2(n_1642),
.B(n_1635),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1673),
.A2(n_1454),
.B(n_1437),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1706),
.B(n_1599),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1671),
.B(n_1607),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1664),
.A2(n_1490),
.B(n_1454),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1694),
.B(n_922),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1700),
.A2(n_1490),
.B(n_1454),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1692),
.B(n_1727),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1712),
.B(n_1610),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1663),
.B(n_922),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1707),
.A2(n_1596),
.B1(n_1645),
.B2(n_1611),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1657),
.B(n_1629),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1713),
.A2(n_1522),
.B(n_1490),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1661),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1683),
.A2(n_1126),
.B(n_1476),
.C(n_1475),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1679),
.B(n_1579),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1718),
.A2(n_1522),
.B(n_1596),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1668),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1695),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1667),
.B(n_1566),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1708),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1721),
.B(n_1597),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1726),
.B(n_1598),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1689),
.B(n_1569),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1708),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1715),
.B(n_1696),
.Y(n_1775)
);

OR2x6_ASAP7_75t_L g1776 ( 
.A(n_1757),
.B(n_1666),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1729),
.B(n_1599),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1770),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1738),
.B(n_1710),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1775),
.A2(n_1645),
.B(n_1720),
.Y(n_1780)
);

O2A1O1Ixp5_ASAP7_75t_L g1781 ( 
.A1(n_1735),
.A2(n_1686),
.B(n_1701),
.C(n_1690),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1775),
.A2(n_1756),
.B(n_1737),
.Y(n_1782)
);

OR2x6_ASAP7_75t_L g1783 ( 
.A(n_1740),
.B(n_1666),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1742),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1763),
.Y(n_1785)
);

BUFx12f_ASAP7_75t_L g1786 ( 
.A(n_1736),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1768),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1732),
.A2(n_1720),
.B(n_1705),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1731),
.B(n_1719),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_L g1790 ( 
.A(n_1733),
.B(n_1620),
.Y(n_1790)
);

OR2x6_ASAP7_75t_L g1791 ( 
.A(n_1748),
.B(n_1666),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1728),
.A2(n_1754),
.B(n_1750),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1753),
.B(n_1711),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1749),
.B(n_1714),
.Y(n_1794)
);

A2O1A1Ixp33_ASAP7_75t_L g1795 ( 
.A1(n_1735),
.A2(n_1696),
.B(n_1725),
.C(n_1722),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1774),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1731),
.A2(n_1697),
.B1(n_1705),
.B2(n_1691),
.Y(n_1797)
);

INVx11_ASAP7_75t_L g1798 ( 
.A(n_1734),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1747),
.B(n_1627),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1739),
.A2(n_1608),
.B1(n_1697),
.B2(n_1573),
.Y(n_1800)
);

BUFx4f_ASAP7_75t_L g1801 ( 
.A(n_1742),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1744),
.A2(n_1522),
.B(n_1535),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1746),
.A2(n_1681),
.B(n_1724),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1739),
.B(n_1627),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1743),
.B(n_1717),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1751),
.A2(n_1699),
.B(n_1481),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1761),
.B(n_1711),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1759),
.B(n_1643),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_SL g1809 ( 
.A(n_1759),
.B(n_1693),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1758),
.B(n_1687),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1771),
.B(n_1083),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1741),
.A2(n_1762),
.B(n_1766),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1772),
.B(n_1716),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1730),
.Y(n_1814)
);

AO32x1_ASAP7_75t_L g1815 ( 
.A1(n_1760),
.A2(n_1723),
.A3(n_1716),
.B1(n_1648),
.B2(n_1649),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1765),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1767),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1755),
.A2(n_1581),
.B1(n_1585),
.B2(n_1554),
.Y(n_1818)
);

AOI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1752),
.A2(n_1559),
.B(n_1549),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1769),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1773),
.B(n_1723),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1755),
.B(n_1221),
.Y(n_1822)
);

BUFx12f_ASAP7_75t_L g1823 ( 
.A(n_1786),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1816),
.B(n_1764),
.Y(n_1824)
);

OAI21x1_ASAP7_75t_SL g1825 ( 
.A1(n_1793),
.A2(n_1616),
.B(n_1659),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1789),
.A2(n_1086),
.B(n_762),
.Y(n_1826)
);

OAI21x1_ASAP7_75t_L g1827 ( 
.A1(n_1782),
.A2(n_1516),
.B(n_1698),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1812),
.A2(n_1494),
.B(n_1734),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1784),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1820),
.B(n_1745),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1795),
.A2(n_1614),
.B(n_1406),
.Y(n_1831)
);

NOR2xp67_ASAP7_75t_SL g1832 ( 
.A(n_1799),
.B(n_1093),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1814),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_L g1834 ( 
.A(n_1777),
.B(n_1745),
.Y(n_1834)
);

OAI21x1_ASAP7_75t_L g1835 ( 
.A1(n_1792),
.A2(n_1698),
.B(n_1571),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1785),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1810),
.B(n_1198),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1793),
.B(n_1594),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1796),
.Y(n_1839)
);

OAI21x1_ASAP7_75t_L g1840 ( 
.A1(n_1802),
.A2(n_1575),
.B(n_1570),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1805),
.B(n_1813),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1791),
.B(n_1674),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1781),
.A2(n_1811),
.B(n_1818),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1791),
.B(n_1494),
.Y(n_1844)
);

AOI21x1_ASAP7_75t_SL g1845 ( 
.A1(n_1821),
.A2(n_1088),
.B(n_1083),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1803),
.A2(n_1586),
.B(n_1577),
.Y(n_1846)
);

BUFx2_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1813),
.B(n_1659),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_L g1849 ( 
.A(n_1800),
.B(n_1311),
.C(n_1150),
.Y(n_1849)
);

OAI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1804),
.A2(n_1009),
.B(n_992),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1780),
.A2(n_1449),
.B(n_1443),
.Y(n_1851)
);

AO31x2_ASAP7_75t_L g1852 ( 
.A1(n_1788),
.A2(n_1449),
.A3(n_1459),
.B(n_1443),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1779),
.A2(n_1654),
.B1(n_1562),
.B2(n_1595),
.Y(n_1853)
);

OAI21x1_ASAP7_75t_L g1854 ( 
.A1(n_1806),
.A2(n_1819),
.B(n_1821),
.Y(n_1854)
);

AO22x2_ASAP7_75t_L g1855 ( 
.A1(n_1797),
.A2(n_1685),
.B1(n_1704),
.B2(n_1682),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1787),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1791),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1794),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1783),
.A2(n_1016),
.B1(n_1614),
.B2(n_1406),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1776),
.Y(n_1860)
);

OAI21x1_ASAP7_75t_L g1861 ( 
.A1(n_1807),
.A2(n_1588),
.B(n_1587),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1790),
.A2(n_1016),
.B(n_1036),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1783),
.A2(n_1215),
.B1(n_1182),
.B2(n_1157),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1807),
.A2(n_1593),
.B(n_1589),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1783),
.B(n_1776),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1778),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1815),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1815),
.A2(n_1465),
.B(n_1462),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1809),
.B(n_1682),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1776),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1822),
.B(n_1685),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1809),
.B(n_1704),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1797),
.A2(n_1808),
.B(n_799),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1801),
.B(n_1457),
.Y(n_1874)
);

A2O1A1Ixp33_ASAP7_75t_L g1875 ( 
.A1(n_1801),
.A2(n_1003),
.B(n_677),
.C(n_726),
.Y(n_1875)
);

NAND3x1_ASAP7_75t_L g1876 ( 
.A(n_1784),
.B(n_1004),
.C(n_754),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1798),
.A2(n_1600),
.B(n_1644),
.Y(n_1877)
);

AO31x2_ASAP7_75t_L g1878 ( 
.A1(n_1782),
.A2(n_1466),
.A3(n_1465),
.B(n_1655),
.Y(n_1878)
);

OAI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1782),
.A2(n_1651),
.B(n_1647),
.Y(n_1879)
);

AND3x4_ASAP7_75t_L g1880 ( 
.A(n_1814),
.B(n_1091),
.C(n_1088),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1816),
.B(n_1014),
.Y(n_1881)
);

AOI222xp33_ASAP7_75t_L g1882 ( 
.A1(n_1826),
.A2(n_810),
.B1(n_796),
.B2(n_449),
.C1(n_462),
.C2(n_656),
.Y(n_1882)
);

BUFx4f_ASAP7_75t_L g1883 ( 
.A(n_1823),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1856),
.Y(n_1884)
);

NAND2x1p5_ASAP7_75t_L g1885 ( 
.A(n_1834),
.B(n_1652),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1856),
.Y(n_1886)
);

A2O1A1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1862),
.A2(n_562),
.B(n_993),
.C(n_991),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1847),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1828),
.A2(n_1831),
.B(n_1843),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1870),
.B(n_1480),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1858),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1833),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1841),
.B(n_978),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1836),
.Y(n_1894)
);

A2O1A1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1873),
.A2(n_996),
.B(n_999),
.C(n_998),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1839),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1839),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1823),
.Y(n_1898)
);

NAND2x1p5_ASAP7_75t_L g1899 ( 
.A(n_1874),
.B(n_1653),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1860),
.Y(n_1900)
);

INVx5_ASAP7_75t_L g1901 ( 
.A(n_1829),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1829),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1860),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1880),
.A2(n_454),
.B1(n_462),
.B2(n_449),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1866),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1842),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1857),
.B(n_811),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1875),
.A2(n_1001),
.B(n_1000),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1870),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1865),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1832),
.B(n_1457),
.Y(n_1911)
);

NAND2x1_ASAP7_75t_L g1912 ( 
.A(n_1824),
.B(n_1523),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1855),
.Y(n_1913)
);

CKINVDCx20_ASAP7_75t_R g1914 ( 
.A(n_1838),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_1874),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1844),
.B(n_812),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1853),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1855),
.Y(n_1918)
);

A2O1A1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1875),
.A2(n_1849),
.B(n_1850),
.C(n_1859),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1828),
.A2(n_1742),
.B(n_1638),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_1871),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1869),
.B(n_813),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1855),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1872),
.B(n_814),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1825),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1830),
.B(n_820),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1848),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1854),
.B(n_821),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1881),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1877),
.B(n_1484),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1880),
.A2(n_652),
.B1(n_656),
.B2(n_454),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1861),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1835),
.B(n_1487),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1876),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1876),
.Y(n_1935)
);

AOI21xp33_ASAP7_75t_L g1936 ( 
.A1(n_1837),
.A2(n_1150),
.B(n_1311),
.Y(n_1936)
);

INVx1_ASAP7_75t_SL g1937 ( 
.A(n_1851),
.Y(n_1937)
);

INVx2_ASAP7_75t_SL g1938 ( 
.A(n_1863),
.Y(n_1938)
);

BUFx10_ASAP7_75t_L g1939 ( 
.A(n_1845),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1851),
.A2(n_1433),
.B(n_1402),
.Y(n_1940)
);

NOR2x1_ASAP7_75t_SL g1941 ( 
.A(n_1867),
.B(n_1845),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1864),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1827),
.B(n_1623),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1879),
.B(n_1044),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1878),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1878),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1878),
.Y(n_1947)
);

CKINVDCx11_ASAP7_75t_R g1948 ( 
.A(n_1867),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1852),
.B(n_1492),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1852),
.B(n_1846),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1840),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1868),
.Y(n_1952)
);

OR2x2_ASAP7_75t_SL g1953 ( 
.A(n_1849),
.B(n_1215),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1856),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1847),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1838),
.B(n_1540),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1911),
.B(n_1457),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1884),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1883),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1883),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1894),
.Y(n_1961)
);

BUFx12f_ASAP7_75t_L g1962 ( 
.A(n_1898),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1905),
.Y(n_1963)
);

CKINVDCx11_ASAP7_75t_R g1964 ( 
.A(n_1914),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_SL g1965 ( 
.A1(n_1889),
.A2(n_1118),
.B1(n_658),
.B2(n_659),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_1929),
.Y(n_1966)
);

BUFx8_ASAP7_75t_L g1967 ( 
.A(n_1916),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1888),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1954),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1910),
.B(n_824),
.Y(n_1970)
);

CKINVDCx16_ASAP7_75t_R g1971 ( 
.A(n_1915),
.Y(n_1971)
);

INVx6_ASAP7_75t_L g1972 ( 
.A(n_1901),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1902),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1891),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1902),
.Y(n_1975)
);

BUFx12f_ASAP7_75t_L g1976 ( 
.A(n_1953),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1906),
.B(n_826),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1900),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1886),
.Y(n_1979)
);

BUFx10_ASAP7_75t_L g1980 ( 
.A(n_1944),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1882),
.A2(n_851),
.B(n_838),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1955),
.Y(n_1982)
);

INVx6_ASAP7_75t_L g1983 ( 
.A(n_1901),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1882),
.A2(n_828),
.B1(n_829),
.B2(n_827),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1896),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1925),
.A2(n_831),
.B1(n_832),
.B2(n_830),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_SL g1987 ( 
.A1(n_1911),
.A2(n_658),
.B1(n_659),
.B2(n_652),
.Y(n_1987)
);

INVx6_ASAP7_75t_L g1988 ( 
.A(n_1901),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1909),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_SL g1990 ( 
.A1(n_1935),
.A2(n_670),
.B1(n_672),
.B2(n_660),
.Y(n_1990)
);

OAI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1887),
.A2(n_1002),
.B(n_979),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1892),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1927),
.B(n_606),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1903),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1938),
.A2(n_1931),
.B1(n_1904),
.B2(n_1936),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1904),
.A2(n_670),
.B1(n_672),
.B2(n_660),
.Y(n_1996)
);

NAND2x1p5_ASAP7_75t_L g1997 ( 
.A(n_1912),
.B(n_1942),
.Y(n_1997)
);

OAI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1931),
.A2(n_675),
.B1(n_676),
.B2(n_673),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1902),
.Y(n_1999)
);

BUFx10_ASAP7_75t_L g2000 ( 
.A(n_1890),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1919),
.A2(n_675),
.B1(n_676),
.B2(n_673),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1921),
.B(n_1897),
.Y(n_2002)
);

CKINVDCx20_ASAP7_75t_R g2003 ( 
.A(n_1917),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1934),
.A2(n_697),
.B1(n_699),
.B2(n_696),
.Y(n_2004)
);

CKINVDCx20_ASAP7_75t_R g2005 ( 
.A(n_1956),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1936),
.A2(n_839),
.B1(n_840),
.B2(n_837),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1913),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1934),
.A2(n_842),
.B1(n_845),
.B2(n_841),
.Y(n_2008)
);

CKINVDCx6p67_ASAP7_75t_R g2009 ( 
.A(n_1907),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1918),
.B(n_847),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1948),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_SL g2012 ( 
.A1(n_1957),
.A2(n_1920),
.B(n_1899),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1981),
.A2(n_1928),
.B(n_1893),
.Y(n_2013)
);

O2A1O1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1981),
.A2(n_1908),
.B(n_1895),
.C(n_1893),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1989),
.B(n_1923),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1989),
.B(n_1941),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1965),
.A2(n_1885),
.B1(n_1924),
.B2(n_1922),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1995),
.A2(n_1926),
.B1(n_1890),
.B2(n_1930),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2007),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1958),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1969),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_SL g2022 ( 
.A1(n_2001),
.A2(n_1930),
.B(n_1908),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1994),
.Y(n_2023)
);

AOI21xp5_ASAP7_75t_SL g2024 ( 
.A1(n_2001),
.A2(n_1950),
.B(n_1932),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1978),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1968),
.B(n_1950),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1982),
.B(n_2002),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1974),
.Y(n_2028)
);

O2A1O1Ixp33_ASAP7_75t_L g2029 ( 
.A1(n_1996),
.A2(n_1937),
.B(n_1943),
.C(n_1952),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1973),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_2010),
.B(n_1943),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1961),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_2010),
.B(n_1943),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1997),
.A2(n_1937),
.B(n_1940),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1964),
.Y(n_2035)
);

BUFx3_ASAP7_75t_L g2036 ( 
.A(n_1967),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_SL g2037 ( 
.A1(n_1997),
.A2(n_1951),
.B(n_1933),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1979),
.B(n_1951),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1972),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_SL g2040 ( 
.A1(n_2011),
.A2(n_1971),
.B1(n_2003),
.B2(n_1976),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1963),
.Y(n_2041)
);

OA21x2_ASAP7_75t_L g2042 ( 
.A1(n_1985),
.A2(n_1946),
.B(n_1945),
.Y(n_2042)
);

OR2x6_ASAP7_75t_L g2043 ( 
.A(n_2012),
.B(n_1972),
.Y(n_2043)
);

BUFx10_ASAP7_75t_L g2044 ( 
.A(n_2035),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2025),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2025),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_2036),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_2036),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2023),
.B(n_1970),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_2015),
.Y(n_2050)
);

AOI21xp33_ASAP7_75t_L g2051 ( 
.A1(n_2029),
.A2(n_1993),
.B(n_1996),
.Y(n_2051)
);

AND2x4_ASAP7_75t_SL g2052 ( 
.A(n_2027),
.B(n_2000),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_2030),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2039),
.B(n_1980),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_2039),
.B(n_1999),
.Y(n_2055)
);

NOR3xp33_ASAP7_75t_SL g2056 ( 
.A(n_2035),
.B(n_1960),
.C(n_1959),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_2018),
.A2(n_1939),
.B1(n_1967),
.B2(n_2009),
.Y(n_2057)
);

OAI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2022),
.A2(n_1993),
.B(n_1977),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_2039),
.B(n_1999),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_2040),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_2015),
.B(n_1947),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2019),
.Y(n_2062)
);

AOI21xp33_ASAP7_75t_L g2063 ( 
.A1(n_2014),
.A2(n_2004),
.B(n_2006),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2042),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_2030),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_2032),
.B(n_2041),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_2016),
.B(n_1999),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_2016),
.Y(n_2068)
);

OA21x2_ASAP7_75t_L g2069 ( 
.A1(n_2064),
.A2(n_2034),
.B(n_2013),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_L g2070 ( 
.A(n_2060),
.B(n_1980),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2061),
.B(n_2028),
.Y(n_2071)
);

INVxp67_ASAP7_75t_SL g2072 ( 
.A(n_2064),
.Y(n_2072)
);

AO21x2_ASAP7_75t_L g2073 ( 
.A1(n_2051),
.A2(n_2024),
.B(n_2012),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2061),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2066),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2045),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_2065),
.Y(n_2077)
);

AO21x2_ASAP7_75t_L g2078 ( 
.A1(n_2058),
.A2(n_2024),
.B(n_2037),
.Y(n_2078)
);

OA21x2_ASAP7_75t_L g2079 ( 
.A1(n_2046),
.A2(n_2021),
.B(n_2020),
.Y(n_2079)
);

OR2x6_ASAP7_75t_L g2080 ( 
.A(n_2043),
.B(n_2037),
.Y(n_2080)
);

NOR3xp33_ASAP7_75t_L g2081 ( 
.A(n_2063),
.B(n_1998),
.C(n_1990),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2066),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2068),
.B(n_2026),
.Y(n_2083)
);

BUFx12f_ASAP7_75t_L g2084 ( 
.A(n_2044),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_2050),
.Y(n_2085)
);

AO21x2_ASAP7_75t_L g2086 ( 
.A1(n_2062),
.A2(n_2004),
.B(n_2038),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2049),
.B(n_2027),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_2053),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2053),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2043),
.B(n_2026),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_2053),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2053),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2065),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_L g2094 ( 
.A(n_2047),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2043),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_2043),
.B(n_2038),
.Y(n_2096)
);

AOI221xp5_ASAP7_75t_L g2097 ( 
.A1(n_2060),
.A2(n_1990),
.B1(n_699),
.B2(n_700),
.C(n_697),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2054),
.B(n_2038),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_SL g2099 ( 
.A1(n_2048),
.A2(n_2017),
.B(n_1966),
.Y(n_2099)
);

NAND3xp33_ASAP7_75t_L g2100 ( 
.A(n_2047),
.B(n_1987),
.C(n_1984),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_2085),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2078),
.B(n_2054),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2085),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2081),
.A2(n_2047),
.B1(n_2048),
.B2(n_2057),
.Y(n_2104)
);

INVx3_ASAP7_75t_L g2105 ( 
.A(n_2084),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_2084),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2079),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2079),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2071),
.B(n_2067),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2071),
.B(n_2067),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_2081),
.A2(n_2047),
.B1(n_2033),
.B2(n_2031),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2078),
.B(n_2067),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_2070),
.B(n_2044),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2075),
.Y(n_2114)
);

OAI22xp33_ASAP7_75t_SL g2115 ( 
.A1(n_2077),
.A2(n_1992),
.B1(n_1983),
.B2(n_1988),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_2094),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2078),
.B(n_2055),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2093),
.B(n_2087),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_2094),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2079),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2079),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2078),
.B(n_2055),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2105),
.B(n_2094),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2113),
.A2(n_2073),
.B1(n_2069),
.B2(n_2084),
.Y(n_2124)
);

OAI211xp5_ASAP7_75t_L g2125 ( 
.A1(n_2104),
.A2(n_2097),
.B(n_2099),
.C(n_2069),
.Y(n_2125)
);

BUFx8_ASAP7_75t_SL g2126 ( 
.A(n_2106),
.Y(n_2126)
);

NAND2xp33_ASAP7_75t_R g2127 ( 
.A(n_2106),
.B(n_2105),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2115),
.A2(n_2097),
.B1(n_2073),
.B2(n_2100),
.C(n_2086),
.Y(n_2128)
);

AOI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_2115),
.A2(n_2073),
.B1(n_2100),
.B2(n_2086),
.C(n_2095),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2116),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2105),
.B(n_2083),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_2112),
.A2(n_2093),
.B(n_2072),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2105),
.B(n_2083),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_2118),
.B(n_2044),
.Y(n_2134)
);

OR2x6_ASAP7_75t_L g2135 ( 
.A(n_2116),
.B(n_2094),
.Y(n_2135)
);

OAI31xp33_ASAP7_75t_SL g2136 ( 
.A1(n_2112),
.A2(n_2122),
.A3(n_2117),
.B(n_2102),
.Y(n_2136)
);

OAI221xp5_ASAP7_75t_L g2137 ( 
.A1(n_2111),
.A2(n_2110),
.B1(n_2109),
.B2(n_2080),
.C(n_2095),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_SL g2138 ( 
.A1(n_2117),
.A2(n_2073),
.B1(n_2069),
.B2(n_2086),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2101),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2135),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2131),
.B(n_2094),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_2135),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2139),
.B(n_2103),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2133),
.B(n_2094),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2134),
.B(n_2094),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2123),
.B(n_2093),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2135),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2126),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2148),
.B(n_2123),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2146),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_2142),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2143),
.B(n_2136),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2141),
.Y(n_2153)
);

INVxp67_ASAP7_75t_L g2154 ( 
.A(n_2144),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2140),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2151),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2155),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2149),
.B(n_2147),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_2150),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2153),
.B(n_2145),
.Y(n_2160)
);

INVx1_ASAP7_75t_SL g2161 ( 
.A(n_2158),
.Y(n_2161)
);

NOR2x1p5_ASAP7_75t_L g2162 ( 
.A(n_2156),
.B(n_2143),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2159),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2161),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2163),
.B(n_2158),
.Y(n_2165)
);

OAI311xp33_ASAP7_75t_L g2166 ( 
.A1(n_2165),
.A2(n_2152),
.A3(n_2154),
.B1(n_2128),
.C1(n_2157),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2164),
.B(n_2160),
.Y(n_2167)
);

OAI221xp5_ASAP7_75t_L g2168 ( 
.A1(n_2165),
.A2(n_2125),
.B1(n_2136),
.B2(n_2152),
.C(n_2129),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2167),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_SL g2170 ( 
.A1(n_2168),
.A2(n_2162),
.B(n_2160),
.Y(n_2170)
);

NAND2xp33_ASAP7_75t_L g2171 ( 
.A(n_2169),
.B(n_2130),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2170),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2169),
.B(n_2103),
.Y(n_2173)
);

NAND4xp25_ASAP7_75t_L g2174 ( 
.A(n_2172),
.B(n_2173),
.C(n_2127),
.D(n_2166),
.Y(n_2174)
);

NAND3xp33_ASAP7_75t_L g2175 ( 
.A(n_2171),
.B(n_2138),
.C(n_2124),
.Y(n_2175)
);

OAI211xp5_ASAP7_75t_L g2176 ( 
.A1(n_2172),
.A2(n_1551),
.B(n_2137),
.C(n_2119),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2171),
.Y(n_2177)
);

AOI221x1_ASAP7_75t_L g2178 ( 
.A1(n_2174),
.A2(n_2114),
.B1(n_2122),
.B2(n_2102),
.C(n_2092),
.Y(n_2178)
);

INVxp33_ASAP7_75t_L g2179 ( 
.A(n_2177),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2176),
.B(n_2132),
.Y(n_2180)
);

NOR4xp25_ASAP7_75t_L g2181 ( 
.A(n_2175),
.B(n_2114),
.C(n_1054),
.D(n_1042),
.Y(n_2181)
);

NOR2x1_ASAP7_75t_L g2182 ( 
.A(n_2180),
.B(n_1092),
.Y(n_2182)
);

NOR3xp33_ASAP7_75t_L g2183 ( 
.A(n_2179),
.B(n_1203),
.C(n_1199),
.Y(n_2183)
);

NOR3xp33_ASAP7_75t_L g2184 ( 
.A(n_2181),
.B(n_2178),
.C(n_1095),
.Y(n_2184)
);

NOR2x1_ASAP7_75t_L g2185 ( 
.A(n_2180),
.B(n_849),
.Y(n_2185)
);

AOI221xp5_ASAP7_75t_L g2186 ( 
.A1(n_2181),
.A2(n_706),
.B1(n_710),
.B2(n_700),
.C(n_696),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_2179),
.B(n_2089),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2178),
.B(n_2089),
.Y(n_2188)
);

O2A1O1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_2179),
.A2(n_1991),
.B(n_851),
.C(n_888),
.Y(n_2189)
);

OAI211xp5_ASAP7_75t_L g2190 ( 
.A1(n_2181),
.A2(n_710),
.B(n_731),
.C(n_706),
.Y(n_2190)
);

AND2x2_ASAP7_75t_SL g2191 ( 
.A(n_2181),
.B(n_1986),
.Y(n_2191)
);

AOI211xp5_ASAP7_75t_L g2192 ( 
.A1(n_2181),
.A2(n_748),
.B(n_731),
.C(n_853),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2179),
.A2(n_1081),
.B(n_1052),
.Y(n_2193)
);

NOR3xp33_ASAP7_75t_L g2194 ( 
.A(n_2180),
.B(n_855),
.C(n_854),
.Y(n_2194)
);

NOR2x1_ASAP7_75t_L g2195 ( 
.A(n_2180),
.B(n_857),
.Y(n_2195)
);

NAND4xp25_ASAP7_75t_L g2196 ( 
.A(n_2178),
.B(n_2008),
.C(n_1991),
.D(n_860),
.Y(n_2196)
);

NOR3xp33_ASAP7_75t_SL g2197 ( 
.A(n_2190),
.B(n_611),
.C(n_607),
.Y(n_2197)
);

NAND3xp33_ASAP7_75t_L g2198 ( 
.A(n_2187),
.B(n_1640),
.C(n_615),
.Y(n_2198)
);

OAI211xp5_ASAP7_75t_SL g2199 ( 
.A1(n_2192),
.A2(n_861),
.B(n_863),
.C(n_858),
.Y(n_2199)
);

NAND4xp25_ASAP7_75t_L g2200 ( 
.A(n_2186),
.B(n_866),
.C(n_867),
.D(n_864),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2188),
.B(n_2089),
.Y(n_2201)
);

NAND3xp33_ASAP7_75t_L g2202 ( 
.A(n_2184),
.B(n_624),
.C(n_613),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2183),
.B(n_2191),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2189),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_SL g2205 ( 
.A(n_2193),
.B(n_2194),
.C(n_2182),
.Y(n_2205)
);

NOR3xp33_ASAP7_75t_L g2206 ( 
.A(n_2185),
.B(n_869),
.C(n_868),
.Y(n_2206)
);

AOI211x1_ASAP7_75t_SL g2207 ( 
.A1(n_2196),
.A2(n_2108),
.B(n_2120),
.C(n_2107),
.Y(n_2207)
);

NOR4xp25_ASAP7_75t_L g2208 ( 
.A(n_2195),
.B(n_872),
.C(n_2077),
.D(n_2092),
.Y(n_2208)
);

NAND3x1_ASAP7_75t_SL g2209 ( 
.A(n_2186),
.B(n_1080),
.C(n_630),
.Y(n_2209)
);

AOI21xp33_ASAP7_75t_SL g2210 ( 
.A1(n_2184),
.A2(n_631),
.B(n_629),
.Y(n_2210)
);

NAND3xp33_ASAP7_75t_L g2211 ( 
.A(n_2187),
.B(n_641),
.C(n_632),
.Y(n_2211)
);

NOR3xp33_ASAP7_75t_L g2212 ( 
.A(n_2190),
.B(n_755),
.C(n_751),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2187),
.B(n_2088),
.Y(n_2213)
);

AOI211xp5_ASAP7_75t_L g2214 ( 
.A1(n_2187),
.A2(n_650),
.B(n_711),
.C(n_647),
.Y(n_2214)
);

OAI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2188),
.A2(n_2056),
.B1(n_1080),
.B2(n_2072),
.C(n_2080),
.Y(n_2215)
);

AOI211xp5_ASAP7_75t_L g2216 ( 
.A1(n_2187),
.A2(n_716),
.B(n_717),
.C(n_715),
.Y(n_2216)
);

AND4x1_ASAP7_75t_L g2217 ( 
.A(n_2192),
.B(n_759),
.C(n_760),
.D(n_758),
.Y(n_2217)
);

AOI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2187),
.A2(n_2108),
.B1(n_2120),
.B2(n_2107),
.C(n_2091),
.Y(n_2218)
);

NAND4xp25_ASAP7_75t_L g2219 ( 
.A(n_2187),
.B(n_763),
.C(n_766),
.D(n_761),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_2187),
.B(n_1962),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2188),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2187),
.B(n_2109),
.Y(n_2222)
);

NAND3xp33_ASAP7_75t_L g2223 ( 
.A(n_2187),
.B(n_720),
.C(n_718),
.Y(n_2223)
);

NOR5xp2_ASAP7_75t_L g2224 ( 
.A(n_2190),
.B(n_771),
.C(n_768),
.D(n_2082),
.E(n_2075),
.Y(n_2224)
);

NOR3xp33_ASAP7_75t_L g2225 ( 
.A(n_2190),
.B(n_728),
.C(n_721),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2188),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_2187),
.B(n_2110),
.Y(n_2227)
);

AOI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_2193),
.A2(n_888),
.B(n_838),
.Y(n_2228)
);

AOI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_2187),
.A2(n_2086),
.B1(n_2121),
.B2(n_2108),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2187),
.B(n_2082),
.Y(n_2230)
);

OAI211xp5_ASAP7_75t_SL g2231 ( 
.A1(n_2192),
.A2(n_900),
.B(n_903),
.C(n_898),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2187),
.B(n_2069),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2188),
.Y(n_2233)
);

AND3x1_ASAP7_75t_L g2234 ( 
.A(n_2184),
.B(n_2121),
.C(n_2120),
.Y(n_2234)
);

NOR3xp33_ASAP7_75t_L g2235 ( 
.A(n_2190),
.B(n_738),
.C(n_736),
.Y(n_2235)
);

NAND4xp25_ASAP7_75t_L g2236 ( 
.A(n_2187),
.B(n_907),
.C(n_909),
.D(n_906),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2188),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_2187),
.B(n_2005),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_2187),
.B(n_2098),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2188),
.Y(n_2240)
);

NAND3xp33_ASAP7_75t_L g2241 ( 
.A(n_2187),
.B(n_905),
.C(n_894),
.Y(n_2241)
);

NOR3xp33_ASAP7_75t_L g2242 ( 
.A(n_2190),
.B(n_913),
.C(n_912),
.Y(n_2242)
);

CKINVDCx14_ASAP7_75t_R g2243 ( 
.A(n_2203),
.Y(n_2243)
);

AOI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2227),
.A2(n_2107),
.B1(n_2096),
.B2(n_2090),
.Y(n_2244)
);

OAI22xp33_ASAP7_75t_L g2245 ( 
.A1(n_2222),
.A2(n_2080),
.B1(n_2074),
.B2(n_2098),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2201),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2238),
.B(n_2069),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_R g2248 ( 
.A(n_2205),
.B(n_2),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2213),
.B(n_2074),
.Y(n_2249)
);

NOR2xp67_ASAP7_75t_L g2250 ( 
.A(n_2241),
.B(n_3),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2234),
.Y(n_2251)
);

NOR4xp75_ASAP7_75t_L g2252 ( 
.A(n_2215),
.B(n_2232),
.C(n_2230),
.D(n_2209),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2239),
.B(n_2076),
.Y(n_2253)
);

INVx1_ASAP7_75t_SL g2254 ( 
.A(n_2221),
.Y(n_2254)
);

O2A1O1Ixp33_ASAP7_75t_L g2255 ( 
.A1(n_2210),
.A2(n_905),
.B(n_894),
.C(n_2080),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2220),
.B(n_2076),
.Y(n_2256)
);

BUFx2_ASAP7_75t_L g2257 ( 
.A(n_2240),
.Y(n_2257)
);

AOI211xp5_ASAP7_75t_L g2258 ( 
.A1(n_2226),
.A2(n_918),
.B(n_921),
.C(n_916),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2233),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2237),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2207),
.Y(n_2261)
);

A2O1A1Ixp33_ASAP7_75t_L g2262 ( 
.A1(n_2228),
.A2(n_2074),
.B(n_2076),
.C(n_2090),
.Y(n_2262)
);

NAND3xp33_ASAP7_75t_L g2263 ( 
.A(n_2197),
.B(n_925),
.C(n_924),
.Y(n_2263)
);

NOR4xp25_ASAP7_75t_L g2264 ( 
.A(n_2198),
.B(n_927),
.C(n_929),
.D(n_926),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2208),
.B(n_2090),
.Y(n_2265)
);

AOI221xp5_ASAP7_75t_L g2266 ( 
.A1(n_2202),
.A2(n_939),
.B1(n_941),
.B2(n_938),
.C(n_937),
.Y(n_2266)
);

O2A1O1Ixp33_ASAP7_75t_L g2267 ( 
.A1(n_2225),
.A2(n_2080),
.B(n_946),
.C(n_950),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2217),
.B(n_2087),
.Y(n_2268)
);

XNOR2x1_ASAP7_75t_L g2269 ( 
.A(n_2204),
.B(n_3),
.Y(n_2269)
);

NAND3xp33_ASAP7_75t_L g2270 ( 
.A(n_2214),
.B(n_953),
.C(n_945),
.Y(n_2270)
);

AOI211xp5_ASAP7_75t_L g2271 ( 
.A1(n_2235),
.A2(n_955),
.B(n_954),
.C(n_441),
.Y(n_2271)
);

AOI211x1_ASAP7_75t_L g2272 ( 
.A1(n_2211),
.A2(n_2083),
.B(n_6),
.C(n_4),
.Y(n_2272)
);

NAND2xp33_ASAP7_75t_SL g2273 ( 
.A(n_2224),
.B(n_2096),
.Y(n_2273)
);

INVx2_ASAP7_75t_SL g2274 ( 
.A(n_2223),
.Y(n_2274)
);

AOI221xp5_ASAP7_75t_SL g2275 ( 
.A1(n_2216),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.C(n_10),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_R g2276 ( 
.A(n_2199),
.B(n_5),
.Y(n_2276)
);

AOI222xp33_ASAP7_75t_L g2277 ( 
.A1(n_2218),
.A2(n_2096),
.B1(n_2059),
.B2(n_2055),
.C1(n_453),
.C2(n_441),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2212),
.B(n_2096),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2229),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2231),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2242),
.B(n_2096),
.Y(n_2281)
);

INVxp67_ASAP7_75t_L g2282 ( 
.A(n_2219),
.Y(n_2282)
);

OAI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2206),
.A2(n_2080),
.B(n_2059),
.Y(n_2283)
);

OAI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2236),
.A2(n_2059),
.B(n_448),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2200),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_2201),
.Y(n_2286)
);

O2A1O1Ixp33_ASAP7_75t_L g2287 ( 
.A1(n_2210),
.A2(n_14),
.B(n_11),
.C(n_12),
.Y(n_2287)
);

INVx1_ASAP7_75t_SL g2288 ( 
.A(n_2201),
.Y(n_2288)
);

AND4x1_ASAP7_75t_L g2289 ( 
.A(n_2197),
.B(n_20),
.C(n_18),
.D(n_19),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_2222),
.B(n_20),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2227),
.A2(n_2079),
.B1(n_2052),
.B2(n_2030),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2222),
.Y(n_2292)
);

OA211x2_ASAP7_75t_L g2293 ( 
.A1(n_2203),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2227),
.B(n_23),
.Y(n_2294)
);

NOR2xp67_ASAP7_75t_L g2295 ( 
.A(n_2241),
.B(n_24),
.Y(n_2295)
);

NOR3xp33_ASAP7_75t_L g2296 ( 
.A(n_2209),
.B(n_448),
.C(n_439),
.Y(n_2296)
);

O2A1O1Ixp33_ASAP7_75t_L g2297 ( 
.A1(n_2210),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_2297)
);

AOI221xp5_ASAP7_75t_L g2298 ( 
.A1(n_2220),
.A2(n_463),
.B1(n_655),
.B2(n_460),
.C(n_453),
.Y(n_2298)
);

AOI332xp33_ASAP7_75t_L g2299 ( 
.A1(n_2221),
.A2(n_25),
.A3(n_27),
.B1(n_29),
.B2(n_30),
.B3(n_31),
.C1(n_32),
.C2(n_33),
.Y(n_2299)
);

OAI221xp5_ASAP7_75t_L g2300 ( 
.A1(n_2201),
.A2(n_655),
.B1(n_657),
.B2(n_463),
.C(n_460),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_R g2301 ( 
.A(n_2205),
.B(n_32),
.Y(n_2301)
);

NOR2x1_ASAP7_75t_L g2302 ( 
.A(n_2241),
.B(n_34),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_2230),
.B(n_2052),
.Y(n_2303)
);

NOR2x1p5_ASAP7_75t_L g2304 ( 
.A(n_2201),
.B(n_657),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2222),
.A2(n_2030),
.B1(n_1983),
.B2(n_1988),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2222),
.A2(n_1983),
.B1(n_1988),
.B2(n_1972),
.Y(n_2306)
);

O2A1O1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_2210),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2307)
);

INVxp67_ASAP7_75t_SL g2308 ( 
.A(n_2201),
.Y(n_2308)
);

NAND2xp33_ASAP7_75t_R g2309 ( 
.A(n_2197),
.B(n_38),
.Y(n_2309)
);

NAND2xp33_ASAP7_75t_SL g2310 ( 
.A(n_2197),
.B(n_662),
.Y(n_2310)
);

OAI31xp33_ASAP7_75t_L g2311 ( 
.A1(n_2215),
.A2(n_42),
.A3(n_40),
.B(n_41),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2201),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_2201),
.Y(n_2313)
);

INVx1_ASAP7_75t_SL g2314 ( 
.A(n_2201),
.Y(n_2314)
);

NAND3x1_ASAP7_75t_L g2315 ( 
.A(n_2217),
.B(n_42),
.C(n_43),
.Y(n_2315)
);

AOI211xp5_ASAP7_75t_L g2316 ( 
.A1(n_2201),
.A2(n_674),
.B(n_678),
.C(n_662),
.Y(n_2316)
);

CKINVDCx16_ASAP7_75t_R g2317 ( 
.A(n_2203),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2222),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_R g2319 ( 
.A(n_2205),
.B(n_43),
.Y(n_2319)
);

INVx1_ASAP7_75t_SL g2320 ( 
.A(n_2201),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2222),
.Y(n_2321)
);

INVx1_ASAP7_75t_SL g2322 ( 
.A(n_2201),
.Y(n_2322)
);

OAI32xp33_ASAP7_75t_L g2323 ( 
.A1(n_2201),
.A2(n_48),
.A3(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2222),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2228),
.A2(n_678),
.B(n_674),
.Y(n_2325)
);

AOI322xp5_ASAP7_75t_L g2326 ( 
.A1(n_2227),
.A2(n_2031),
.A3(n_2033),
.B1(n_51),
.B2(n_53),
.C1(n_54),
.C2(n_56),
.Y(n_2326)
);

NAND4xp25_ASAP7_75t_SL g2327 ( 
.A(n_2222),
.B(n_51),
.C(n_48),
.D(n_50),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2227),
.A2(n_688),
.B1(n_689),
.B2(n_681),
.Y(n_2328)
);

NOR2x1_ASAP7_75t_L g2329 ( 
.A(n_2327),
.B(n_53),
.Y(n_2329)
);

NOR2x1_ASAP7_75t_L g2330 ( 
.A(n_2269),
.B(n_57),
.Y(n_2330)
);

NAND2x1_ASAP7_75t_L g2331 ( 
.A(n_2272),
.B(n_1204),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2303),
.Y(n_2332)
);

XOR2x2_ASAP7_75t_L g2333 ( 
.A(n_2289),
.B(n_58),
.Y(n_2333)
);

OR2x2_ASAP7_75t_L g2334 ( 
.A(n_2265),
.B(n_59),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2294),
.B(n_60),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2293),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2281),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2249),
.Y(n_2338)
);

NAND4xp75_ASAP7_75t_L g2339 ( 
.A(n_2259),
.B(n_64),
.C(n_61),
.D(n_62),
.Y(n_2339)
);

NOR2x1_ASAP7_75t_L g2340 ( 
.A(n_2263),
.B(n_67),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2303),
.B(n_68),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2278),
.Y(n_2342)
);

INVx1_ASAP7_75t_SL g2343 ( 
.A(n_2248),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2290),
.B(n_69),
.Y(n_2344)
);

NAND4xp75_ASAP7_75t_L g2345 ( 
.A(n_2260),
.B(n_72),
.C(n_70),
.D(n_71),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2315),
.Y(n_2346)
);

NAND4xp75_ASAP7_75t_L g2347 ( 
.A(n_2292),
.B(n_72),
.C(n_70),
.D(n_71),
.Y(n_2347)
);

NOR2x1_ASAP7_75t_L g2348 ( 
.A(n_2257),
.B(n_73),
.Y(n_2348)
);

NOR2x1_ASAP7_75t_L g2349 ( 
.A(n_2302),
.B(n_75),
.Y(n_2349)
);

NOR2x1p5_ASAP7_75t_L g2350 ( 
.A(n_2308),
.B(n_681),
.Y(n_2350)
);

INVx1_ASAP7_75t_SL g2351 ( 
.A(n_2301),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2318),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2288),
.B(n_76),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2244),
.A2(n_689),
.B1(n_694),
.B2(n_688),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2251),
.Y(n_2355)
);

AND2x4_ASAP7_75t_L g2356 ( 
.A(n_2250),
.B(n_76),
.Y(n_2356)
);

NOR2x1_ASAP7_75t_L g2357 ( 
.A(n_2261),
.B(n_77),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2253),
.Y(n_2358)
);

NAND2x1p5_ASAP7_75t_SL g2359 ( 
.A(n_2274),
.B(n_79),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2286),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2321),
.B(n_2031),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2324),
.B(n_2033),
.Y(n_2362)
);

NAND4xp75_ASAP7_75t_L g2363 ( 
.A(n_2275),
.B(n_83),
.C(n_79),
.D(n_81),
.Y(n_2363)
);

AOI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2243),
.A2(n_698),
.B1(n_739),
.B2(n_694),
.Y(n_2364)
);

CKINVDCx20_ASAP7_75t_R g2365 ( 
.A(n_2317),
.Y(n_2365)
);

AOI22xp5_ASAP7_75t_L g2366 ( 
.A1(n_2273),
.A2(n_739),
.B1(n_740),
.B2(n_698),
.Y(n_2366)
);

NOR2x1_ASAP7_75t_L g2367 ( 
.A(n_2304),
.B(n_84),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2268),
.B(n_1973),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2254),
.B(n_85),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2309),
.A2(n_743),
.B1(n_746),
.B2(n_740),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2312),
.Y(n_2371)
);

INVx4_ASAP7_75t_L g2372 ( 
.A(n_2280),
.Y(n_2372)
);

OA22x2_ASAP7_75t_L g2373 ( 
.A1(n_2284),
.A2(n_746),
.B1(n_743),
.B2(n_87),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2246),
.Y(n_2374)
);

INVxp67_ASAP7_75t_SL g2375 ( 
.A(n_2295),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2287),
.Y(n_2376)
);

NOR2x1p5_ASAP7_75t_L g2377 ( 
.A(n_2285),
.B(n_531),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2313),
.A2(n_1504),
.B1(n_546),
.B2(n_555),
.Y(n_2378)
);

NAND3xp33_ASAP7_75t_L g2379 ( 
.A(n_2271),
.B(n_560),
.C(n_535),
.Y(n_2379)
);

XNOR2xp5_ASAP7_75t_L g2380 ( 
.A(n_2252),
.B(n_85),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2297),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2307),
.Y(n_2382)
);

AND2x2_ASAP7_75t_SL g2383 ( 
.A(n_2296),
.B(n_86),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_2319),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2256),
.Y(n_2385)
);

NOR2x1_ASAP7_75t_L g2386 ( 
.A(n_2270),
.B(n_89),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2314),
.B(n_89),
.Y(n_2387)
);

NAND3xp33_ASAP7_75t_L g2388 ( 
.A(n_2298),
.B(n_566),
.C(n_561),
.Y(n_2388)
);

OR2x2_ASAP7_75t_L g2389 ( 
.A(n_2320),
.B(n_90),
.Y(n_2389)
);

NOR2xp67_ASAP7_75t_L g2390 ( 
.A(n_2325),
.B(n_93),
.Y(n_2390)
);

BUFx3_ASAP7_75t_L g2391 ( 
.A(n_2322),
.Y(n_2391)
);

NOR2x1_ASAP7_75t_L g2392 ( 
.A(n_2279),
.B(n_94),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2283),
.B(n_94),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2277),
.B(n_95),
.Y(n_2394)
);

OAI211xp5_ASAP7_75t_SL g2395 ( 
.A1(n_2311),
.A2(n_100),
.B(n_97),
.C(n_98),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2323),
.Y(n_2396)
);

NOR2x1_ASAP7_75t_L g2397 ( 
.A(n_2300),
.B(n_100),
.Y(n_2397)
);

NOR3xp33_ASAP7_75t_L g2398 ( 
.A(n_2355),
.B(n_2371),
.C(n_2360),
.Y(n_2398)
);

NAND4xp75_ASAP7_75t_L g2399 ( 
.A(n_2357),
.B(n_2328),
.C(n_2266),
.D(n_2247),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2341),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2353),
.B(n_2326),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2361),
.B(n_2264),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2362),
.B(n_2282),
.Y(n_2403)
);

AND2x4_ASAP7_75t_L g2404 ( 
.A(n_2348),
.B(n_2262),
.Y(n_2404)
);

NOR4xp25_ASAP7_75t_L g2405 ( 
.A(n_2396),
.B(n_2267),
.C(n_2255),
.D(n_2276),
.Y(n_2405)
);

NOR3xp33_ASAP7_75t_L g2406 ( 
.A(n_2369),
.B(n_2310),
.C(n_2316),
.Y(n_2406)
);

NAND4xp75_ASAP7_75t_L g2407 ( 
.A(n_2392),
.B(n_2330),
.C(n_2349),
.D(n_2340),
.Y(n_2407)
);

NOR2x1_ASAP7_75t_L g2408 ( 
.A(n_2389),
.B(n_2299),
.Y(n_2408)
);

NOR5xp2_ASAP7_75t_L g2409 ( 
.A(n_2375),
.B(n_2382),
.C(n_2381),
.D(n_2376),
.E(n_2337),
.Y(n_2409)
);

NOR2x1_ASAP7_75t_L g2410 ( 
.A(n_2365),
.B(n_2245),
.Y(n_2410)
);

AND4x1_ASAP7_75t_L g2411 ( 
.A(n_2336),
.B(n_2258),
.C(n_2291),
.D(n_2305),
.Y(n_2411)
);

NAND4xp75_ASAP7_75t_L g2412 ( 
.A(n_2386),
.B(n_2306),
.C(n_103),
.D(n_101),
.Y(n_2412)
);

NAND4xp75_ASAP7_75t_L g2413 ( 
.A(n_2329),
.B(n_106),
.C(n_102),
.D(n_105),
.Y(n_2413)
);

NOR2x1p5_ASAP7_75t_L g2414 ( 
.A(n_2363),
.B(n_567),
.Y(n_2414)
);

AOI221xp5_ASAP7_75t_L g2415 ( 
.A1(n_2395),
.A2(n_582),
.B1(n_586),
.B2(n_581),
.C(n_575),
.Y(n_2415)
);

NAND4xp25_ASAP7_75t_L g2416 ( 
.A(n_2352),
.B(n_107),
.C(n_102),
.D(n_105),
.Y(n_2416)
);

NAND5xp2_ASAP7_75t_L g2417 ( 
.A(n_2342),
.B(n_112),
.C(n_110),
.D(n_111),
.E(n_115),
.Y(n_2417)
);

NOR3xp33_ASAP7_75t_L g2418 ( 
.A(n_2338),
.B(n_1204),
.C(n_1197),
.Y(n_2418)
);

NOR2x2_ASAP7_75t_L g2419 ( 
.A(n_2332),
.B(n_111),
.Y(n_2419)
);

NOR3xp33_ASAP7_75t_L g2420 ( 
.A(n_2372),
.B(n_1197),
.C(n_1183),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2334),
.Y(n_2421)
);

NOR4xp75_ASAP7_75t_SL g2422 ( 
.A(n_2394),
.B(n_2344),
.C(n_2354),
.D(n_2380),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2339),
.Y(n_2423)
);

NAND3x1_ASAP7_75t_L g2424 ( 
.A(n_2366),
.B(n_118),
.C(n_119),
.Y(n_2424)
);

NOR3xp33_ASAP7_75t_L g2425 ( 
.A(n_2374),
.B(n_1202),
.C(n_1183),
.Y(n_2425)
);

HB1xp67_ASAP7_75t_L g2426 ( 
.A(n_2345),
.Y(n_2426)
);

OAI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_2333),
.A2(n_589),
.B(n_588),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2387),
.B(n_2335),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2387),
.Y(n_2429)
);

NOR3xp33_ASAP7_75t_SL g2430 ( 
.A(n_2385),
.B(n_596),
.C(n_592),
.Y(n_2430)
);

NOR2x1_ASAP7_75t_L g2431 ( 
.A(n_2347),
.B(n_119),
.Y(n_2431)
);

NAND3xp33_ASAP7_75t_L g2432 ( 
.A(n_2370),
.B(n_601),
.C(n_598),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2359),
.Y(n_2433)
);

AND4x1_ASAP7_75t_L g2434 ( 
.A(n_2367),
.B(n_124),
.C(n_120),
.D(n_123),
.Y(n_2434)
);

AOI211xp5_ASAP7_75t_L g2435 ( 
.A1(n_2343),
.A2(n_2351),
.B(n_2393),
.C(n_2356),
.Y(n_2435)
);

NAND5xp2_ASAP7_75t_L g2436 ( 
.A(n_2368),
.B(n_124),
.C(n_120),
.D(n_123),
.E(n_125),
.Y(n_2436)
);

NOR3xp33_ASAP7_75t_SL g2437 ( 
.A(n_2358),
.B(n_605),
.C(n_602),
.Y(n_2437)
);

INVx2_ASAP7_75t_SL g2438 ( 
.A(n_2356),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2331),
.Y(n_2439)
);

NAND5xp2_ASAP7_75t_L g2440 ( 
.A(n_2384),
.B(n_127),
.C(n_125),
.D(n_126),
.E(n_128),
.Y(n_2440)
);

NAND3x2_ASAP7_75t_L g2441 ( 
.A(n_2393),
.B(n_126),
.C(n_127),
.Y(n_2441)
);

OA22x2_ASAP7_75t_L g2442 ( 
.A1(n_2346),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_2442)
);

NOR4xp25_ASAP7_75t_L g2443 ( 
.A(n_2379),
.B(n_134),
.C(n_131),
.D(n_133),
.Y(n_2443)
);

NOR2xp67_ASAP7_75t_L g2444 ( 
.A(n_2390),
.B(n_134),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2391),
.B(n_135),
.Y(n_2445)
);

NOR3xp33_ASAP7_75t_L g2446 ( 
.A(n_2388),
.B(n_1211),
.C(n_1202),
.Y(n_2446)
);

NOR3x2_ASAP7_75t_L g2447 ( 
.A(n_2350),
.B(n_2373),
.C(n_2377),
.Y(n_2447)
);

NAND4xp75_ASAP7_75t_L g2448 ( 
.A(n_2397),
.B(n_2383),
.C(n_2378),
.D(n_2364),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_2348),
.B(n_135),
.Y(n_2449)
);

NOR3xp33_ASAP7_75t_L g2450 ( 
.A(n_2355),
.B(n_1211),
.C(n_610),
.Y(n_2450)
);

AO211x2_ASAP7_75t_L g2451 ( 
.A1(n_2355),
.A2(n_139),
.B(n_136),
.C(n_138),
.Y(n_2451)
);

NOR5xp2_ASAP7_75t_L g2452 ( 
.A(n_2355),
.B(n_141),
.C(n_136),
.D(n_140),
.E(n_142),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2387),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2361),
.B(n_1973),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2445),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_2400),
.Y(n_2456)
);

NAND2xp33_ASAP7_75t_SL g2457 ( 
.A(n_2414),
.B(n_608),
.Y(n_2457)
);

BUFx2_ASAP7_75t_L g2458 ( 
.A(n_2449),
.Y(n_2458)
);

INVx1_ASAP7_75t_SL g2459 ( 
.A(n_2419),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2449),
.Y(n_2460)
);

HB1xp67_ASAP7_75t_L g2461 ( 
.A(n_2451),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2434),
.Y(n_2462)
);

BUFx2_ASAP7_75t_L g2463 ( 
.A(n_2442),
.Y(n_2463)
);

NOR2x1_ASAP7_75t_L g2464 ( 
.A(n_2407),
.B(n_140),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_2423),
.Y(n_2465)
);

INVx1_ASAP7_75t_SL g2466 ( 
.A(n_2445),
.Y(n_2466)
);

CKINVDCx20_ASAP7_75t_R g2467 ( 
.A(n_2426),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2438),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2413),
.Y(n_2469)
);

NAND3xp33_ASAP7_75t_L g2470 ( 
.A(n_2398),
.B(n_2435),
.C(n_2410),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2433),
.Y(n_2471)
);

INVx1_ASAP7_75t_SL g2472 ( 
.A(n_2431),
.Y(n_2472)
);

HB1xp67_ASAP7_75t_L g2473 ( 
.A(n_2444),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_2403),
.Y(n_2474)
);

CKINVDCx20_ASAP7_75t_R g2475 ( 
.A(n_2401),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_2429),
.Y(n_2476)
);

INVx3_ASAP7_75t_SL g2477 ( 
.A(n_2453),
.Y(n_2477)
);

HB1xp67_ASAP7_75t_L g2478 ( 
.A(n_2404),
.Y(n_2478)
);

INVx3_ASAP7_75t_SL g2479 ( 
.A(n_2404),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2454),
.Y(n_2480)
);

HB1xp67_ASAP7_75t_L g2481 ( 
.A(n_2412),
.Y(n_2481)
);

CKINVDCx16_ASAP7_75t_R g2482 ( 
.A(n_2408),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2424),
.Y(n_2483)
);

CKINVDCx20_ASAP7_75t_R g2484 ( 
.A(n_2428),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2421),
.Y(n_2485)
);

CKINVDCx20_ASAP7_75t_R g2486 ( 
.A(n_2402),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2409),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2439),
.Y(n_2488)
);

NAND3xp33_ASAP7_75t_L g2489 ( 
.A(n_2415),
.B(n_620),
.C(n_616),
.Y(n_2489)
);

CKINVDCx20_ASAP7_75t_R g2490 ( 
.A(n_2430),
.Y(n_2490)
);

NAND3xp33_ASAP7_75t_SL g2491 ( 
.A(n_2411),
.B(n_627),
.C(n_623),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2436),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_2441),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2440),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_R g2495 ( 
.A(n_2422),
.B(n_142),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2443),
.B(n_2000),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2437),
.Y(n_2497)
);

NAND4xp25_ASAP7_75t_L g2498 ( 
.A(n_2406),
.B(n_2417),
.C(n_2452),
.D(n_2450),
.Y(n_2498)
);

INVxp67_ASAP7_75t_L g2499 ( 
.A(n_2416),
.Y(n_2499)
);

INVx1_ASAP7_75t_SL g2500 ( 
.A(n_2447),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2427),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2448),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2399),
.Y(n_2503)
);

XNOR2x1_ASAP7_75t_L g2504 ( 
.A(n_2432),
.B(n_2405),
.Y(n_2504)
);

O2A1O1Ixp33_ASAP7_75t_L g2505 ( 
.A1(n_2420),
.A2(n_146),
.B(n_143),
.C(n_145),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2425),
.B(n_143),
.Y(n_2506)
);

NAND3xp33_ASAP7_75t_L g2507 ( 
.A(n_2446),
.B(n_635),
.C(n_634),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2418),
.Y(n_2508)
);

BUFx12f_ASAP7_75t_L g2509 ( 
.A(n_2438),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2449),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2449),
.Y(n_2511)
);

HB1xp67_ASAP7_75t_L g2512 ( 
.A(n_2451),
.Y(n_2512)
);

OR2x2_ASAP7_75t_L g2513 ( 
.A(n_2436),
.B(n_145),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2454),
.B(n_147),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2449),
.Y(n_2515)
);

CKINVDCx16_ASAP7_75t_R g2516 ( 
.A(n_2410),
.Y(n_2516)
);

INVx1_ASAP7_75t_SL g2517 ( 
.A(n_2495),
.Y(n_2517)
);

OAI221xp5_ASAP7_75t_L g2518 ( 
.A1(n_2470),
.A2(n_636),
.B1(n_644),
.B2(n_648),
.C(n_703),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2514),
.Y(n_2519)
);

OAI221xp5_ASAP7_75t_SL g2520 ( 
.A1(n_2500),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.C(n_151),
.Y(n_2520)
);

OAI322xp33_ASAP7_75t_SL g2521 ( 
.A1(n_2502),
.A2(n_151),
.A3(n_152),
.B1(n_153),
.B2(n_154),
.C1(n_155),
.C2(n_156),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2513),
.Y(n_2522)
);

OAI322xp33_ASAP7_75t_L g2523 ( 
.A1(n_2516),
.A2(n_152),
.A3(n_154),
.B1(n_155),
.B2(n_156),
.C1(n_157),
.C2(n_158),
.Y(n_2523)
);

AOI221xp5_ASAP7_75t_L g2524 ( 
.A1(n_2487),
.A2(n_713),
.B1(n_730),
.B2(n_732),
.C(n_733),
.Y(n_2524)
);

HB1xp67_ASAP7_75t_L g2525 ( 
.A(n_2464),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2461),
.Y(n_2526)
);

O2A1O1Ixp33_ASAP7_75t_L g2527 ( 
.A1(n_2478),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2527)
);

AOI322xp5_ASAP7_75t_L g2528 ( 
.A1(n_2472),
.A2(n_2496),
.A3(n_2482),
.B1(n_2512),
.B2(n_2459),
.C1(n_2466),
.C2(n_2469),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2458),
.Y(n_2529)
);

INVxp67_ASAP7_75t_L g2530 ( 
.A(n_2473),
.Y(n_2530)
);

A2O1A1Ixp33_ASAP7_75t_L g2531 ( 
.A1(n_2505),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2531)
);

OAI211xp5_ASAP7_75t_SL g2532 ( 
.A1(n_2499),
.A2(n_164),
.B(n_161),
.C(n_162),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2463),
.B(n_162),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2510),
.Y(n_2534)
);

AOI22xp33_ASAP7_75t_L g2535 ( 
.A1(n_2509),
.A2(n_1975),
.B1(n_168),
.B2(n_165),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2462),
.Y(n_2536)
);

NAND4xp25_ASAP7_75t_L g2537 ( 
.A(n_2498),
.B(n_170),
.C(n_166),
.D(n_169),
.Y(n_2537)
);

AOI322xp5_ASAP7_75t_L g2538 ( 
.A1(n_2503),
.A2(n_169),
.A3(n_171),
.B1(n_172),
.B2(n_177),
.C1(n_179),
.C2(n_180),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2468),
.Y(n_2539)
);

A2O1A1Ixp33_ASAP7_75t_L g2540 ( 
.A1(n_2494),
.A2(n_179),
.B(n_171),
.C(n_177),
.Y(n_2540)
);

INVxp33_ASAP7_75t_SL g2541 ( 
.A(n_2481),
.Y(n_2541)
);

OAI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2475),
.A2(n_1975),
.B1(n_182),
.B2(n_180),
.Y(n_2542)
);

AOI322xp5_ASAP7_75t_L g2543 ( 
.A1(n_2465),
.A2(n_2467),
.A3(n_2492),
.B1(n_2484),
.B2(n_2515),
.C1(n_2460),
.C2(n_2511),
.Y(n_2543)
);

OAI322xp33_ASAP7_75t_L g2544 ( 
.A1(n_2479),
.A2(n_181),
.A3(n_182),
.B1(n_183),
.B2(n_184),
.C1(n_186),
.C2(n_187),
.Y(n_2544)
);

AOI22xp33_ASAP7_75t_L g2545 ( 
.A1(n_2487),
.A2(n_1975),
.B1(n_184),
.B2(n_1263),
.Y(n_2545)
);

AOI322xp5_ASAP7_75t_L g2546 ( 
.A1(n_2480),
.A2(n_1933),
.A3(n_1949),
.B1(n_1527),
.B2(n_1498),
.C1(n_1502),
.C2(n_1510),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2476),
.A2(n_1263),
.B1(n_1278),
.B2(n_1232),
.Y(n_2547)
);

NOR2x1_ASAP7_75t_L g2548 ( 
.A(n_2455),
.B(n_1232),
.Y(n_2548)
);

OAI22x1_ASAP7_75t_L g2549 ( 
.A1(n_2477),
.A2(n_1278),
.B1(n_1280),
.B2(n_1263),
.Y(n_2549)
);

OAI22xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2490),
.A2(n_1078),
.B1(n_1096),
.B2(n_1072),
.Y(n_2550)
);

AOI322xp5_ASAP7_75t_L g2551 ( 
.A1(n_2486),
.A2(n_1949),
.A3(n_1507),
.B1(n_1656),
.B2(n_1520),
.C1(n_1518),
.C2(n_1511),
.Y(n_2551)
);

NOR3xp33_ASAP7_75t_L g2552 ( 
.A(n_2491),
.B(n_1254),
.C(n_1278),
.Y(n_2552)
);

AOI322xp5_ASAP7_75t_L g2553 ( 
.A1(n_2483),
.A2(n_1503),
.A3(n_1520),
.B1(n_1518),
.B2(n_1511),
.C1(n_1509),
.C2(n_1488),
.Y(n_2553)
);

OAI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_2456),
.A2(n_1365),
.B1(n_1072),
.B2(n_1122),
.Y(n_2554)
);

INVxp67_ASAP7_75t_L g2555 ( 
.A(n_2487),
.Y(n_2555)
);

NAND4xp25_ASAP7_75t_L g2556 ( 
.A(n_2493),
.B(n_1253),
.C(n_1226),
.D(n_1236),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2506),
.Y(n_2557)
);

INVx3_ASAP7_75t_L g2558 ( 
.A(n_2474),
.Y(n_2558)
);

AO22x2_ASAP7_75t_L g2559 ( 
.A1(n_2517),
.A2(n_2504),
.B1(n_2501),
.B2(n_2507),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2526),
.A2(n_2471),
.B1(n_2485),
.B2(n_2488),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2533),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2525),
.Y(n_2562)
);

AO22x2_ASAP7_75t_L g2563 ( 
.A1(n_2519),
.A2(n_2507),
.B1(n_2489),
.B2(n_2457),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2555),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2529),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2534),
.Y(n_2566)
);

OAI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2530),
.A2(n_2497),
.B1(n_2508),
.B2(n_1072),
.Y(n_2567)
);

OAI22x1_ASAP7_75t_L g2568 ( 
.A1(n_2539),
.A2(n_1280),
.B1(n_1096),
.B2(n_1098),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2548),
.Y(n_2569)
);

CKINVDCx20_ASAP7_75t_R g2570 ( 
.A(n_2558),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2541),
.A2(n_1280),
.B1(n_1276),
.B2(n_1250),
.Y(n_2571)
);

AO22x2_ASAP7_75t_L g2572 ( 
.A1(n_2522),
.A2(n_1301),
.B1(n_1265),
.B2(n_1267),
.Y(n_2572)
);

HB1xp67_ASAP7_75t_L g2573 ( 
.A(n_2542),
.Y(n_2573)
);

AOI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2536),
.A2(n_1282),
.B1(n_1295),
.B2(n_1240),
.Y(n_2574)
);

OAI22x1_ASAP7_75t_L g2575 ( 
.A1(n_2558),
.A2(n_1078),
.B1(n_1096),
.B2(n_1098),
.Y(n_2575)
);

OAI22xp5_ASAP7_75t_SL g2576 ( 
.A1(n_2545),
.A2(n_1078),
.B1(n_1098),
.B2(n_1121),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2531),
.Y(n_2577)
);

OAI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_2535),
.A2(n_1122),
.B1(n_1121),
.B2(n_1308),
.Y(n_2578)
);

OAI22x1_ASAP7_75t_L g2579 ( 
.A1(n_2557),
.A2(n_1121),
.B1(n_1122),
.B2(n_1186),
.Y(n_2579)
);

OAI22x1_ASAP7_75t_L g2580 ( 
.A1(n_2547),
.A2(n_1186),
.B1(n_1193),
.B2(n_1207),
.Y(n_2580)
);

AND4x1_ASAP7_75t_L g2581 ( 
.A(n_2527),
.B(n_1314),
.C(n_1305),
.D(n_1300),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2537),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2532),
.Y(n_2583)
);

OAI22xp5_ASAP7_75t_L g2584 ( 
.A1(n_2520),
.A2(n_1245),
.B1(n_1296),
.B2(n_1264),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2523),
.Y(n_2585)
);

AOI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2552),
.A2(n_1274),
.B1(n_1256),
.B2(n_1268),
.Y(n_2586)
);

OAI22xp33_ASAP7_75t_SL g2587 ( 
.A1(n_2518),
.A2(n_2554),
.B1(n_2528),
.B2(n_2543),
.Y(n_2587)
);

OAI311xp33_ASAP7_75t_L g2588 ( 
.A1(n_2565),
.A2(n_2556),
.A3(n_2540),
.B1(n_2524),
.C1(n_2538),
.Y(n_2588)
);

AOI321xp33_ASAP7_75t_L g2589 ( 
.A1(n_2560),
.A2(n_2550),
.A3(n_2521),
.B1(n_2549),
.B2(n_2544),
.C(n_2553),
.Y(n_2589)
);

AOI22xp5_ASAP7_75t_L g2590 ( 
.A1(n_2570),
.A2(n_2551),
.B1(n_2546),
.B2(n_1249),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2566),
.B(n_188),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2564),
.Y(n_2592)
);

NAND3xp33_ASAP7_75t_SL g2593 ( 
.A(n_2562),
.B(n_1262),
.C(n_1259),
.Y(n_2593)
);

XNOR2xp5_ASAP7_75t_L g2594 ( 
.A(n_2581),
.B(n_2561),
.Y(n_2594)
);

XNOR2xp5_ASAP7_75t_L g2595 ( 
.A(n_2582),
.B(n_190),
.Y(n_2595)
);

NOR4xp75_ASAP7_75t_L g2596 ( 
.A(n_2578),
.B(n_1074),
.C(n_1346),
.D(n_1318),
.Y(n_2596)
);

XNOR2x2_ASAP7_75t_L g2597 ( 
.A(n_2559),
.B(n_192),
.Y(n_2597)
);

NAND3xp33_ASAP7_75t_L g2598 ( 
.A(n_2585),
.B(n_1193),
.C(n_1186),
.Y(n_2598)
);

AOI211xp5_ASAP7_75t_L g2599 ( 
.A1(n_2587),
.A2(n_1073),
.B(n_1070),
.C(n_1433),
.Y(n_2599)
);

NAND4xp25_ASAP7_75t_L g2600 ( 
.A(n_2583),
.B(n_1074),
.C(n_1374),
.D(n_1346),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_2573),
.Y(n_2601)
);

NAND3xp33_ASAP7_75t_L g2602 ( 
.A(n_2577),
.B(n_1207),
.C(n_1193),
.Y(n_2602)
);

NAND5xp2_ASAP7_75t_L g2603 ( 
.A(n_2569),
.B(n_2571),
.C(n_2574),
.D(n_2586),
.E(n_2559),
.Y(n_2603)
);

OAI211xp5_ASAP7_75t_SL g2604 ( 
.A1(n_2567),
.A2(n_2563),
.B(n_2584),
.C(n_2576),
.Y(n_2604)
);

NAND4xp25_ASAP7_75t_L g2605 ( 
.A(n_2563),
.B(n_1374),
.C(n_1270),
.D(n_1318),
.Y(n_2605)
);

NAND3xp33_ASAP7_75t_L g2606 ( 
.A(n_2568),
.B(n_2575),
.C(n_2580),
.Y(n_2606)
);

NAND4xp25_ASAP7_75t_SL g2607 ( 
.A(n_2572),
.B(n_2579),
.C(n_195),
.D(n_197),
.Y(n_2607)
);

NAND3xp33_ASAP7_75t_L g2608 ( 
.A(n_2601),
.B(n_2572),
.C(n_1218),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2597),
.Y(n_2609)
);

AO22x2_ASAP7_75t_L g2610 ( 
.A1(n_2592),
.A2(n_2606),
.B1(n_2593),
.B2(n_2591),
.Y(n_2610)
);

AO22x2_ASAP7_75t_L g2611 ( 
.A1(n_2598),
.A2(n_2602),
.B1(n_2588),
.B2(n_2607),
.Y(n_2611)
);

INVxp67_ASAP7_75t_L g2612 ( 
.A(n_2603),
.Y(n_2612)
);

XNOR2xp5_ASAP7_75t_L g2613 ( 
.A(n_2594),
.B(n_193),
.Y(n_2613)
);

OAI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2590),
.A2(n_1218),
.B1(n_1207),
.B2(n_1506),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2604),
.A2(n_1218),
.B(n_1270),
.Y(n_2615)
);

AOI21x1_ASAP7_75t_L g2616 ( 
.A1(n_2595),
.A2(n_1489),
.B(n_1488),
.Y(n_2616)
);

OR2x6_ASAP7_75t_L g2617 ( 
.A(n_2589),
.B(n_1070),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2596),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2605),
.Y(n_2619)
);

OAI22xp33_ASAP7_75t_L g2620 ( 
.A1(n_2600),
.A2(n_1446),
.B1(n_1506),
.B2(n_1073),
.Y(n_2620)
);

AOI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2599),
.A2(n_1285),
.B(n_1283),
.Y(n_2621)
);

XNOR2xp5_ASAP7_75t_L g2622 ( 
.A(n_2601),
.B(n_204),
.Y(n_2622)
);

OAI21x1_ASAP7_75t_SL g2623 ( 
.A1(n_2615),
.A2(n_212),
.B(n_214),
.Y(n_2623)
);

AOI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2612),
.A2(n_1446),
.B1(n_1506),
.B2(n_1073),
.Y(n_2624)
);

OAI21xp5_ASAP7_75t_SL g2625 ( 
.A1(n_2609),
.A2(n_1285),
.B(n_1283),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2618),
.B(n_2622),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2610),
.Y(n_2627)
);

AOI21xp33_ASAP7_75t_L g2628 ( 
.A1(n_2617),
.A2(n_217),
.B(n_218),
.Y(n_2628)
);

OAI22xp5_ASAP7_75t_SL g2629 ( 
.A1(n_2619),
.A2(n_2608),
.B1(n_2613),
.B2(n_2614),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2611),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2616),
.B(n_222),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2620),
.B(n_223),
.Y(n_2632)
);

AOI21xp5_ASAP7_75t_L g2633 ( 
.A1(n_2621),
.A2(n_1261),
.B(n_1241),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2609),
.Y(n_2634)
);

AOI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2634),
.A2(n_2627),
.B1(n_2630),
.B2(n_2626),
.Y(n_2635)
);

OA22x2_ASAP7_75t_L g2636 ( 
.A1(n_2623),
.A2(n_2631),
.B1(n_2632),
.B2(n_2624),
.Y(n_2636)
);

AO21x2_ASAP7_75t_L g2637 ( 
.A1(n_2628),
.A2(n_1509),
.B(n_1503),
.Y(n_2637)
);

AO22x1_ASAP7_75t_L g2638 ( 
.A1(n_2629),
.A2(n_1261),
.B1(n_1247),
.B2(n_1257),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2625),
.A2(n_1309),
.B(n_1354),
.Y(n_2639)
);

AO21x2_ASAP7_75t_L g2640 ( 
.A1(n_2633),
.A2(n_1499),
.B(n_1493),
.Y(n_2640)
);

AOI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_2634),
.A2(n_1309),
.B(n_1354),
.Y(n_2641)
);

OAI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2634),
.A2(n_1506),
.B1(n_1446),
.B2(n_1493),
.Y(n_2642)
);

AOI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2634),
.A2(n_1499),
.B1(n_1489),
.B2(n_1526),
.Y(n_2643)
);

AOI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2635),
.A2(n_1309),
.B(n_1354),
.Y(n_2644)
);

AOI21xp5_ASAP7_75t_L g2645 ( 
.A1(n_2636),
.A2(n_1376),
.B(n_1371),
.Y(n_2645)
);

OA21x2_ASAP7_75t_L g2646 ( 
.A1(n_2641),
.A2(n_224),
.B(n_231),
.Y(n_2646)
);

AOI221xp5_ASAP7_75t_L g2647 ( 
.A1(n_2642),
.A2(n_1323),
.B1(n_1257),
.B2(n_1376),
.C(n_1371),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2639),
.A2(n_1376),
.B(n_1371),
.Y(n_2648)
);

A2O1A1Ixp33_ASAP7_75t_L g2649 ( 
.A1(n_2643),
.A2(n_1376),
.B(n_1371),
.C(n_1366),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2646),
.A2(n_2637),
.B1(n_2638),
.B2(n_2640),
.Y(n_2650)
);

AOI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2645),
.A2(n_1307),
.B1(n_1257),
.B2(n_1366),
.Y(n_2651)
);

AOI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2647),
.A2(n_2648),
.B1(n_2644),
.B2(n_2649),
.Y(n_2652)
);

OA21x2_ASAP7_75t_L g2653 ( 
.A1(n_2650),
.A2(n_232),
.B(n_233),
.Y(n_2653)
);

AOI21xp5_ASAP7_75t_L g2654 ( 
.A1(n_2652),
.A2(n_1366),
.B(n_1362),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2651),
.B(n_238),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2650),
.B(n_239),
.Y(n_2656)
);

OAI21xp5_ASAP7_75t_SL g2657 ( 
.A1(n_2654),
.A2(n_2656),
.B(n_2655),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2653),
.Y(n_2658)
);

AOI221xp5_ASAP7_75t_L g2659 ( 
.A1(n_2658),
.A2(n_1366),
.B1(n_1362),
.B2(n_1350),
.C(n_1323),
.Y(n_2659)
);

AOI221xp5_ASAP7_75t_L g2660 ( 
.A1(n_2657),
.A2(n_1362),
.B1(n_1350),
.B2(n_1323),
.C(n_1307),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2659),
.A2(n_1362),
.B(n_1350),
.Y(n_2661)
);

AOI211xp5_ASAP7_75t_L g2662 ( 
.A1(n_2661),
.A2(n_2660),
.B(n_1350),
.C(n_1323),
.Y(n_2662)
);


endmodule