module fake_jpeg_24090_n_308 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_27),
.Y(n_54)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_59),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_18),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_22),
.B1(n_31),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_72),
.B(n_75),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_24),
.B1(n_17),
.B2(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_17),
.B1(n_34),
.B2(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_31),
.B1(n_34),
.B2(n_26),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_78),
.B1(n_83),
.B2(n_28),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_19),
.B1(n_26),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_19),
.B1(n_32),
.B2(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_38),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_81),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_29),
.B1(n_37),
.B2(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_29),
.B1(n_35),
.B2(n_28),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_101),
.B(n_103),
.Y(n_132)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_89),
.B(n_108),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_1),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_102),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_110),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_28),
.B1(n_21),
.B2(n_27),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_98),
.A2(n_106),
.B1(n_60),
.B2(n_56),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_28),
.B(n_21),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_27),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_60),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_50),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_27),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

CKINVDCx6p67_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_27),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_5),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_28),
.B1(n_21),
.B2(n_36),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_74),
.B1(n_62),
.B2(n_56),
.Y(n_140)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_125),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_77),
.C(n_58),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_138),
.C(n_96),
.Y(n_156)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_55),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_136),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_6),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_21),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_134),
.Y(n_158)
);

AO21x1_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_112),
.B(n_50),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_21),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_137),
.B(n_141),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_7),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_120),
.B1(n_117),
.B2(n_100),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_151),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_82),
.B1(n_87),
.B2(n_119),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_154),
.B(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_166),
.B1(n_172),
.B2(n_180),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_86),
.B1(n_104),
.B2(n_101),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_171),
.B1(n_173),
.B2(n_36),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_167),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_89),
.C(n_118),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_183),
.C(n_143),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_86),
.B(n_115),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_175),
.B(n_182),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_118),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_91),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_174),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_102),
.B1(n_100),
.B2(n_82),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_126),
.A2(n_108),
.B1(n_107),
.B2(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

OAI22x1_ASAP7_75t_SL g180 ( 
.A1(n_132),
.A2(n_21),
.B1(n_28),
.B2(n_77),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_8),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_94),
.C(n_107),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_109),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_125),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_121),
.B(n_153),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_138),
.B(n_151),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_207),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_126),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_130),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_202),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_152),
.B(n_147),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_135),
.B(n_146),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_186),
.A2(n_141),
.B1(n_145),
.B2(n_109),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_216),
.B1(n_164),
.B2(n_156),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_182),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_149),
.C(n_142),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_142),
.C(n_144),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_92),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_92),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_166),
.A2(n_97),
.B1(n_36),
.B2(n_10),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_176),
.B1(n_171),
.B2(n_168),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_218),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_161),
.C(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_222),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_157),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_230),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_184),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_236),
.B(n_237),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_190),
.B1(n_210),
.B2(n_200),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_175),
.B1(n_182),
.B2(n_154),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_234),
.A2(n_195),
.B1(n_207),
.B2(n_192),
.Y(n_259)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_165),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_191),
.B(n_194),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_252),
.B(n_227),
.Y(n_274)
);

INVx3_ASAP7_75t_SL g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_230),
.B(n_204),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_254),
.C(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_213),
.B1(n_217),
.B2(n_200),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_258),
.B1(n_247),
.B2(n_255),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_194),
.B(n_203),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_201),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_209),
.B1(n_198),
.B2(n_212),
.Y(n_258)
);

AOI221xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_229),
.B1(n_220),
.B2(n_235),
.C(n_234),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_238),
.C(n_208),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_263),
.C(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_240),
.C(n_198),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_269),
.B1(n_274),
.B2(n_189),
.Y(n_285)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_224),
.Y(n_270)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_272),
.B(n_259),
.C(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_225),
.C(n_235),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_218),
.B1(n_253),
.B2(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_248),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_283),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_251),
.C(n_219),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_285),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_264),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_183),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_275),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_268),
.B(n_270),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_290),
.B(n_292),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_271),
.B(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_281),
.B1(n_278),
.B2(n_279),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_297),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_284),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_298),
.B1(n_9),
.B2(n_11),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_277),
.C(n_261),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_277),
.B1(n_178),
.B2(n_97),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_302),
.B(n_12),
.CI(n_13),
.CON(n_305),
.SN(n_305)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_9),
.B(n_11),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_301),
.C(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_305),
.B(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_305),
.Y(n_308)
);


endmodule