module fake_jpeg_15444_n_92 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_1),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_37),
.B1(n_41),
.B2(n_40),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_46),
.C(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_39),
.C(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_57),
.B1(n_59),
.B2(n_63),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_67),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_65),
.B(n_66),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_70),
.C(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_26),
.B(n_5),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_83),
.B1(n_79),
.B2(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_69),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_23),
.B1(n_9),
.B2(n_13),
.Y(n_85)
);

OAI31xp33_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_29),
.A3(n_14),
.B(n_15),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_30),
.C(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_32),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_33),
.C(n_18),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_21),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_22),
.CI(n_28),
.CON(n_92),
.SN(n_92)
);


endmodule