module fake_jpeg_20014_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_56),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_57),
.B1(n_52),
.B2(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_66),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_41),
.B1(n_46),
.B2(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_70),
.B1(n_47),
.B2(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_83),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_85),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_87),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_51),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_22),
.C(n_29),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_3),
.B(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_94),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_10),
.B1(n_12),
.B2(n_17),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_88),
.B1(n_81),
.B2(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_7),
.C(n_9),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_101),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_105),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_103),
.B(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_97),
.B1(n_106),
.B2(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_92),
.B1(n_95),
.B2(n_25),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_92),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_113),
.Y(n_114)
);


endmodule