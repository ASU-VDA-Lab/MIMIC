module real_jpeg_26141_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_292;
wire n_286;
wire n_221;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_98)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_65),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_45),
.B1(n_60),
.B2(n_61),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_45),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_52),
.Y(n_123)
);

INVx8_ASAP7_75t_SL g80 ( 
.A(n_7),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_30),
.B1(n_42),
.B2(n_43),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_9),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_70),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_70),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_70),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_11),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_11),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_11),
.B(n_82),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_11),
.B(n_43),
.C(n_57),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_11),
.B(n_154),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_182),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_29),
.C(n_48),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_11),
.A2(n_31),
.B(n_242),
.Y(n_270)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_13),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_13),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_87),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_87),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_15),
.A2(n_74),
.B1(n_86),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_15),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_135),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_135),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_135),
.Y(n_254)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_16),
.B(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_16),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_20),
.B(n_114),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_89),
.B2(n_113),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.C(n_67),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_25),
.A2(n_38),
.B1(n_39),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_25),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_26),
.A2(n_31),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_27),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_27),
.B(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_31),
.A2(n_33),
.B(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_31),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_31),
.A2(n_163),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_31),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_31),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_41),
.A2(n_50),
.B1(n_95),
.B2(n_127),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_43),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_43),
.B(n_249),
.Y(n_248)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_46),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_46),
.A2(n_53),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_50),
.A2(n_127),
.B(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_50),
.A2(n_178),
.B(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_50),
.B(n_182),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_53),
.B(n_179),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_54),
.B(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_66),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_56),
.B1(n_66),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_55),
.A2(n_151),
.B(n_153),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_55),
.A2(n_153),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_56),
.A2(n_64),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_56),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_56),
.A2(n_130),
.B(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_61),
.B1(n_78),
.B2(n_79),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_60),
.A2(n_74),
.A3(n_79),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_61),
.B(n_78),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_61),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_75),
.B(n_83),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_69),
.A2(n_76),
.B1(n_82),
.B2(n_134),
.Y(n_133)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_74),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_76),
.A2(n_84),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_81),
.A2(n_111),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_100),
.B2(n_101),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_99),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_94),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_95),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_95),
.A2(n_230),
.B(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_128),
.C(n_133),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_121),
.B(n_126),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_160)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_152),
.B1(n_154),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_167),
.B(n_293),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_165),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_140),
.B(n_165),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_147),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_147),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_155),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_150),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_160),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_161),
.A2(n_253),
.B1(n_255),
.B2(n_257),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_199),
.B(n_287),
.C(n_292),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_193),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.C(n_185),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_170),
.A2(n_171),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_182),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_184),
.B(n_185),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_281),
.B(n_286),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_231),
.B(n_280),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_220),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_204),
.B(n_220),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_213),
.C(n_217),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_205),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_208),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_227),
.C(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_274),
.B(n_279),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_250),
.B(n_273),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_244),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_244),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_248),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_260),
.B(n_272),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_258),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_266),
.B(n_271),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);


endmodule