module fake_jpeg_10115_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_1),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_16),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_31),
.C(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_57),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_22),
.B1(n_42),
.B2(n_31),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_67),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_40),
.B1(n_44),
.B2(n_28),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_78),
.B1(n_89),
.B2(n_90),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_75),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_30),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_30),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_84),
.C(n_65),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_44),
.B1(n_23),
.B2(n_29),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_23),
.B1(n_20),
.B2(n_24),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_88),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_22),
.Y(n_84)
);

AO22x1_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_61),
.B1(n_64),
.B2(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_32),
.B1(n_27),
.B2(n_31),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_32),
.B1(n_27),
.B2(n_37),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_107),
.B1(n_113),
.B2(n_106),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_105),
.Y(n_127)
);

NAND2x1_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_47),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_75),
.B1(n_87),
.B2(n_88),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_112),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_65),
.C(n_55),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_36),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_77),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_90),
.B(n_68),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_70),
.B1(n_66),
.B2(n_53),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_124),
.B1(n_108),
.B2(n_100),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_78),
.B1(n_87),
.B2(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_126),
.B1(n_129),
.B2(n_102),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_133),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_121),
.C(n_122),
.Y(n_136)
);

NOR4xp25_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_71),
.C(n_69),
.D(n_77),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_4),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_61),
.B1(n_76),
.B2(n_59),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_76),
.B1(n_34),
.B2(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_34),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_101),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_1),
.B(n_4),
.C(n_6),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_4),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_143),
.B1(n_128),
.B2(n_8),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_140),
.B1(n_135),
.B2(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_97),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_142),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_110),
.B1(n_114),
.B2(n_96),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_128),
.B(n_9),
.C(n_10),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_114),
.B1(n_96),
.B2(n_15),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_119),
.B(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_132),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_156),
.B1(n_161),
.B2(n_150),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_131),
.B(n_120),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_158),
.Y(n_169)
);

OAI321xp33_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_122),
.A3(n_121),
.B1(n_129),
.B2(n_133),
.C(n_125),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_164),
.B1(n_144),
.B2(n_146),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_12),
.B1(n_13),
.B2(n_10),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_141),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_136),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.C(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_147),
.C(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_147),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_12),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_7),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_162),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_160),
.C(n_161),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_165),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_184),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_182),
.B(n_181),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_166),
.B(n_176),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_187),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_9),
.B(n_11),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_176),
.B1(n_161),
.B2(n_175),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_183),
.C(n_11),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_9),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_189),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_195),
.C(n_189),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_196),
.Y(n_199)
);


endmodule