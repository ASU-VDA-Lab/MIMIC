module real_jpeg_22741_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_215;
wire n_221;
wire n_286;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_28),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_2),
.A2(n_21),
.B1(n_23),
.B2(n_56),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_56),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_56),
.B1(n_69),
.B2(n_70),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_6),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_21),
.B1(n_23),
.B2(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_32),
.B1(n_48),
.B2(n_50),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_6),
.A2(n_32),
.B1(n_69),
.B2(n_70),
.Y(n_133)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_9),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_21),
.B1(n_23),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_40),
.B1(n_48),
.B2(n_50),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_40),
.B1(n_69),
.B2(n_70),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_21),
.B1(n_23),
.B2(n_35),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_9),
.A2(n_35),
.B1(n_48),
.B2(n_50),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_35),
.B1(n_69),
.B2(n_70),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_20),
.C(n_23),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_9),
.B(n_19),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_9),
.B(n_45),
.C(n_48),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_9),
.B(n_66),
.C(n_69),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_11),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_9),
.B(n_115),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_9),
.B(n_59),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_11),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_88),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_87),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_72),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_16),
.B(n_72),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_16),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_38),
.CI(n_51),
.CON(n_16),
.SN(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B(n_33),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_18),
.A2(n_33),
.B(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_19),
.A2(n_34),
.B1(n_36),
.B2(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_19),
.B(n_36),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_24),
.B1(n_28),
.B2(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_21),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_21),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx6p67_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_23),
.B(n_221),
.Y(n_220)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_27),
.B(n_188),
.Y(n_187)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_42),
.A2(n_47),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_43),
.A2(n_59),
.B1(n_86),
.B2(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_47),
.A2(n_85),
.B(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_50),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_48),
.B(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.C(n_60),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_52),
.B(n_131),
.C(n_139),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_52),
.A2(n_78),
.B1(n_139),
.B2(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_52),
.A2(n_78),
.B1(n_117),
.B2(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_52),
.B(n_117),
.C(n_185),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_60),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_82),
.C(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_60),
.A2(n_76),
.B1(n_83),
.B2(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_71),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_62),
.B(n_105),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_64),
.A2(n_105),
.B1(n_115),
.B2(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_68),
.A2(n_104),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_69),
.B(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_71),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.C(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_73),
.A2(n_79),
.B1(n_82),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_82),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_79),
.B(n_158),
.C(n_167),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_79),
.A2(n_82),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_79),
.A2(n_82),
.B1(n_167),
.B2(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_80),
.A2(n_81),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_82),
.B(n_139),
.C(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_83),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_86),
.Y(n_168)
);

OAI211xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_141),
.B(n_148),
.C(n_287),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_125),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_125),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_110),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_112),
.C(n_120),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_101),
.B(n_106),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_92),
.A2(n_106),
.B1(n_107),
.B2(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_92),
.A2(n_102),
.B1(n_128),
.B2(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_94),
.B(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_100),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_95),
.B(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_102),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_120),
.B2(n_121),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_113),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_117),
.B(n_205),
.C(n_207),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_117),
.A2(n_195),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_130),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_129),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_278),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_132),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_136),
.A2(n_137),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_136),
.A2(n_137),
.B1(n_218),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_137),
.B(n_212),
.C(n_218),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_137),
.B(n_190),
.C(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_139),
.A2(n_140),
.B1(n_181),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_139),
.A2(n_140),
.B1(n_165),
.B2(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_140),
.B(n_165),
.C(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_149),
.C(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_143),
.B(n_144),
.Y(n_287)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_171),
.B(n_286),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_169),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_152),
.B(n_169),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_153),
.B(n_155),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_157),
.B(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_158),
.A2(n_159),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_165),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_192),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_165),
.A2(n_178),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_165),
.B(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_281),
.B(n_285),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_208),
.B(n_267),
.C(n_280),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_197),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_174),
.B(n_197),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_184),
.B2(n_196),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_177),
.B(n_183),
.C(n_196),
.Y(n_268)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_194),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_189),
.A2(n_190),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_241),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.C(n_204),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_199),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_204),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_207),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_266),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_227),
.B(n_265),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_224),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_211),
.B(n_224),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_212),
.A2(n_213),
.B1(n_261),
.B2(n_263),
.Y(n_260)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_258),
.B(n_264),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_252),
.B(n_257),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_244),
.B(n_251),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_236),
.B(n_243),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_233),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_240),
.B(n_242),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_269),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_279),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_276),
.B2(n_277),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_277),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);


endmodule