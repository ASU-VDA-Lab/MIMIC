module fake_jpeg_22071_n_144 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_144);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_35),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_34),
.B(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

OR2x4_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_18),
.B1(n_29),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_48),
.A2(n_63),
.B1(n_68),
.B2(n_71),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_18),
.B1(n_25),
.B2(n_21),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_42),
.B1(n_40),
.B2(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_66),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_31),
.B1(n_17),
.B2(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_46),
.B1(n_33),
.B2(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_75),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_27),
.B1(n_16),
.B2(n_23),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_22),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_92),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_55),
.C(n_70),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_90),
.C(n_88),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_109),
.C(n_74),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_69),
.C(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_81),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_60),
.B(n_21),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_76),
.B(n_75),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_65),
.B1(n_59),
.B2(n_51),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_105),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_51),
.B1(n_49),
.B2(n_72),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_72),
.B1(n_22),
.B2(n_5),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_22),
.C(n_4),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_11),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_12),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_81),
.B(n_98),
.C(n_105),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_124),
.B1(n_102),
.B2(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_73),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_74),
.C(n_77),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_10),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_111),
.B(n_113),
.C(n_107),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_110),
.C(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_108),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_114),
.B(n_110),
.C(n_109),
.D(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_130),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_103),
.C(n_13),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_115),
.B(n_123),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

BUFx4f_ASAP7_75t_SL g136 ( 
.A(n_133),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_136),
.B(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_134),
.B(n_131),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_137),
.C(n_136),
.Y(n_141)
);

AOI221xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_14),
.B1(n_6),
.B2(n_8),
.C(n_3),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_140),
.B1(n_3),
.B2(n_8),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_121),
.B(n_112),
.Y(n_144)
);


endmodule