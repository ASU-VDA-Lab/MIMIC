module fake_jpeg_3439_n_562 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_562);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_562;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_9),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_61),
.Y(n_193)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_20),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_74),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_66),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_67),
.B(n_68),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_71),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_72),
.B(n_84),
.Y(n_168)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_17),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_75),
.Y(n_209)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_79),
.Y(n_198)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_1),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_85),
.B(n_92),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_26),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_36),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_94),
.B(n_97),
.Y(n_208)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_36),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_36),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_108),
.B(n_110),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_2),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_55),
.A2(n_3),
.B(n_4),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_39),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_119),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_54),
.Y(n_114)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_52),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_117),
.B(n_118),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_52),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_42),
.B(n_3),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_123),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_43),
.B1(n_50),
.B2(n_47),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_127),
.B(n_61),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_57),
.B1(n_22),
.B2(n_45),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_130),
.A2(n_132),
.B1(n_140),
.B2(n_145),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_77),
.A2(n_57),
.B1(n_22),
.B2(n_45),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_70),
.A2(n_57),
.B1(n_22),
.B2(n_45),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_89),
.A2(n_27),
.B1(n_47),
.B2(n_43),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_50),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_147),
.B(n_150),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_27),
.B1(n_42),
.B2(n_38),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_149),
.A2(n_154),
.B1(n_155),
.B2(n_172),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_53),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_102),
.B1(n_81),
.B2(n_64),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_58),
.A2(n_53),
.B1(n_51),
.B2(n_19),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_76),
.B(n_37),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_162),
.Y(n_234)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_59),
.A2(n_51),
.B1(n_38),
.B2(n_37),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_80),
.A2(n_27),
.B1(n_25),
.B2(n_19),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_181),
.A2(n_183),
.B1(n_186),
.B2(n_195),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_95),
.A2(n_25),
.B1(n_46),
.B2(n_41),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_66),
.A2(n_99),
.B1(n_75),
.B2(n_109),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_90),
.B(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_188),
.B(n_202),
.Y(n_257)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_91),
.A2(n_41),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_101),
.A2(n_103),
.B1(n_105),
.B2(n_104),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_196),
.A2(n_201),
.B1(n_14),
.B2(n_15),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_63),
.A2(n_46),
.B1(n_41),
.B2(n_7),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_93),
.B(n_4),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_121),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_204),
.B1(n_61),
.B2(n_71),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_121),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_213),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_214),
.B(n_250),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_93),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_215),
.B(n_222),
.Y(n_316)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_216),
.Y(n_331)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_218),
.Y(n_335)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

OR2x4_ASAP7_75t_L g221 ( 
.A(n_160),
.B(n_125),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_221),
.A2(n_253),
.B(n_140),
.C(n_186),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_6),
.Y(n_222)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_230),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_128),
.B(n_9),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_231),
.B(n_232),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_10),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_133),
.B(n_10),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_241),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_235),
.A2(n_179),
.B1(n_132),
.B2(n_130),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_236),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_141),
.B(n_10),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_240),
.Y(n_299)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_239),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_168),
.B(n_137),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_10),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_152),
.B(n_11),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_255),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_243),
.B(n_244),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_162),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_178),
.B(n_11),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_127),
.Y(n_248)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_146),
.B(n_123),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_159),
.Y(n_252)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_127),
.A2(n_123),
.B(n_125),
.C(n_15),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_182),
.B(n_12),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_254),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_14),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_214),
.B1(n_259),
.B2(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_131),
.Y(n_262)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_176),
.Y(n_263)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_263),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_180),
.B(n_163),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_264),
.B(n_266),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_126),
.Y(n_265)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_142),
.Y(n_267)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_169),
.Y(n_268)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_138),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_269),
.A2(n_144),
.B1(n_205),
.B2(n_209),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_158),
.B(n_14),
.C(n_164),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_277),
.C(n_282),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_204),
.B(n_14),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_271),
.B(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_153),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_273),
.Y(n_302)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_175),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_170),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_279),
.Y(n_307)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_161),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_155),
.B(n_172),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_173),
.B(n_199),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_149),
.A2(n_181),
.B(n_183),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_278),
.A2(n_209),
.B(n_135),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_157),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_281),
.Y(n_328)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_145),
.A2(n_201),
.B(n_195),
.Y(n_282)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_161),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_283),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_286),
.A2(n_337),
.B1(n_215),
.B2(n_282),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_290),
.B(n_254),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

AO22x1_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_126),
.B1(n_211),
.B2(n_129),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_250),
.Y(n_338)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_221),
.B(n_135),
.CI(n_151),
.CON(n_301),
.SN(n_301)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_301),
.B(n_252),
.CI(n_219),
.CON(n_362),
.SN(n_362)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_309),
.A2(n_321),
.B(n_255),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_226),
.A2(n_144),
.B1(n_205),
.B2(n_151),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_318),
.A2(n_330),
.B1(n_216),
.B2(n_223),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_277),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_326),
.B(n_247),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_251),
.A2(n_131),
.B1(n_156),
.B2(n_191),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_240),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_237),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_222),
.B(n_156),
.C(n_191),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_279),
.C(n_220),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_246),
.A2(n_276),
.B1(n_234),
.B2(n_257),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_338),
.A2(n_349),
.B1(n_350),
.B2(n_365),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_363),
.C(n_367),
.Y(n_383)
);

AO22x1_ASAP7_75t_L g340 ( 
.A1(n_288),
.A2(n_235),
.B1(n_253),
.B2(n_278),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_323),
.Y(n_341)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_343),
.Y(n_389)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_345),
.A2(n_373),
.B1(n_301),
.B2(n_293),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_258),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_346),
.Y(n_412)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_296),
.Y(n_351)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_352),
.B(n_354),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_312),
.A2(n_249),
.B(n_218),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_328),
.B(n_307),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_299),
.B(n_270),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_224),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_356),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_217),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_254),
.Y(n_361)
);

XNOR2x1_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_370),
.Y(n_396)
);

AOI31xp67_ASAP7_75t_L g400 ( 
.A1(n_362),
.A2(n_294),
.A3(n_320),
.B(n_314),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_299),
.B(n_273),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_288),
.A2(n_262),
.B1(n_227),
.B2(n_220),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_364),
.A2(n_368),
.B1(n_371),
.B2(n_334),
.Y(n_390)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_369),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_284),
.B(n_274),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_290),
.A2(n_336),
.B1(n_321),
.B2(n_312),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_317),
.B(n_225),
.Y(n_369)
);

AOI22x1_ASAP7_75t_L g371 ( 
.A1(n_312),
.A2(n_212),
.B1(n_229),
.B2(n_239),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_374),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_336),
.A2(n_212),
.B1(n_228),
.B2(n_283),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_317),
.B(n_275),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_263),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_376),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_245),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_304),
.B(n_268),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_378),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_368),
.A2(n_286),
.B1(n_332),
.B2(n_293),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_382),
.A2(n_393),
.B1(n_409),
.B2(n_338),
.Y(n_413)
);

AOI32xp33_ASAP7_75t_L g384 ( 
.A1(n_357),
.A2(n_301),
.A3(n_287),
.B1(n_315),
.B2(n_291),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_384),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_387),
.A2(n_394),
.B(n_400),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_390),
.A2(n_411),
.B1(n_410),
.B2(n_406),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_340),
.A2(n_289),
.B1(n_298),
.B2(n_302),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_364),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_402),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_357),
.A2(n_319),
.B1(n_289),
.B2(n_298),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_397),
.A2(n_343),
.B1(n_344),
.B2(n_376),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_363),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_350),
.A2(n_294),
.B(n_320),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_403),
.A2(n_406),
.B(n_410),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_349),
.A2(n_353),
.B(n_345),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_374),
.A2(n_311),
.B1(n_297),
.B2(n_314),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_340),
.A2(n_327),
.B(n_308),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_413),
.A2(n_414),
.B1(n_442),
.B2(n_393),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_390),
.A2(n_378),
.B1(n_377),
.B2(n_373),
.Y(n_414)
);

AOI22x1_ASAP7_75t_L g415 ( 
.A1(n_385),
.A2(n_365),
.B1(n_362),
.B2(n_371),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_418),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_354),
.C(n_369),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_417),
.B(n_420),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_405),
.B(n_402),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_407),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_419),
.B(n_423),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_412),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_421),
.Y(n_453)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_398),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_431),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_370),
.Y(n_425)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_425),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_426),
.B(n_427),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_SL g427 ( 
.A(n_396),
.B(n_362),
.C(n_375),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_372),
.Y(n_428)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_428),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_310),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_429),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_361),
.C(n_371),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_403),
.C(n_394),
.Y(n_444)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_379),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_432),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_327),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_433),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_380),
.B(n_366),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_434),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_385),
.B(n_342),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_436),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_360),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_438),
.A2(n_380),
.B1(n_391),
.B2(n_401),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_439),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_447),
.C(n_456),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_386),
.C(n_382),
.Y(n_447)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_449),
.A2(n_454),
.B1(n_460),
.B2(n_465),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_413),
.A2(n_416),
.B1(n_414),
.B2(n_440),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_386),
.C(n_404),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_408),
.C(n_404),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_459),
.C(n_437),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_384),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_416),
.A2(n_395),
.B1(n_397),
.B2(n_400),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_440),
.A2(n_408),
.B1(n_401),
.B2(n_399),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_419),
.A2(n_399),
.B1(n_381),
.B2(n_379),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_466),
.A2(n_467),
.B1(n_438),
.B2(n_431),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_441),
.A2(n_381),
.B1(n_347),
.B2(n_341),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_427),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_470),
.B(n_472),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_437),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_483),
.Y(n_504)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_421),
.C(n_424),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_481),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_445),
.B(n_359),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_476),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_455),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_478),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_459),
.A2(n_415),
.B(n_435),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_479),
.A2(n_480),
.B1(n_482),
.B2(n_464),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_443),
.A2(n_415),
.B(n_434),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_422),
.C(n_428),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_450),
.A2(n_432),
.B(n_423),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_447),
.B(n_432),
.C(n_329),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_358),
.Y(n_484)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_484),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_450),
.B(n_347),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_486),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_351),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_444),
.B(n_329),
.C(n_348),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_492),
.Y(n_495)
);

OAI22x1_ASAP7_75t_L g489 ( 
.A1(n_452),
.A2(n_311),
.B1(n_331),
.B2(n_322),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_489),
.A2(n_451),
.B1(n_465),
.B2(n_467),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_335),
.Y(n_490)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_490),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_468),
.B(n_446),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_491),
.Y(n_506)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_493),
.A2(n_498),
.B1(n_502),
.B2(n_474),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_477),
.A2(n_463),
.B1(n_461),
.B2(n_464),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_500),
.A2(n_482),
.B(n_460),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_466),
.Y(n_501)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_488),
.A2(n_463),
.B1(n_461),
.B2(n_469),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_469),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_503),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_483),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_511),
.B(n_515),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_478),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_514),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_487),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_472),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_517),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_454),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_499),
.B(n_471),
.C(n_473),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_519),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_452),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_471),
.C(n_486),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_521),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_502),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_498),
.B1(n_496),
.B2(n_449),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_507),
.B(n_446),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_523),
.A2(n_495),
.B(n_505),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_534),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_528),
.B(n_530),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_501),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_531),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_513),
.B(n_509),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_508),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_510),
.B(n_496),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_532),
.B(n_522),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_516),
.B(n_508),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_520),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_536),
.B(n_542),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_525),
.A2(n_518),
.B(n_512),
.Y(n_537)
);

AOI21x1_ASAP7_75t_SL g550 ( 
.A1(n_537),
.A2(n_531),
.B(n_533),
.Y(n_550)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_540),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_514),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_541),
.B(n_485),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_494),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_527),
.B(n_494),
.C(n_470),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_544),
.B(n_527),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_546),
.B(n_548),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_543),
.B(n_534),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_538),
.A2(n_533),
.B(n_493),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_549),
.A2(n_544),
.B(n_453),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_550),
.A2(n_551),
.B(n_539),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_547),
.B(n_541),
.C(n_539),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_553),
.B(n_554),
.Y(n_557)
);

AOI321xp33_ASAP7_75t_L g556 ( 
.A1(n_555),
.A2(n_545),
.A3(n_453),
.B1(n_451),
.B2(n_455),
.C(n_489),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_556),
.A2(n_308),
.B1(n_331),
.B2(n_335),
.Y(n_559)
);

A2O1A1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_557),
.A2(n_552),
.B(n_545),
.C(n_458),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_558),
.B(n_559),
.C(n_305),
.Y(n_560)
);

AOI322xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_269),
.A3(n_305),
.B1(n_325),
.B2(n_322),
.C1(n_256),
.C2(n_230),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_325),
.Y(n_562)
);


endmodule