module fake_jpeg_15773_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_6),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_21),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_7),
.B(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_10),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_7),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_9),
.B(n_11),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.C(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_12),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_26),
.B1(n_28),
.B2(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.C(n_18),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_14),
.B(n_9),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_29),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_20),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_8),
.C(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_11),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_18),
.Y(n_46)
);

AOI322xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.A3(n_45),
.B1(n_11),
.B2(n_2),
.C1(n_5),
.C2(n_6),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_46),
.B(n_5),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_2),
.Y(n_50)
);


endmodule