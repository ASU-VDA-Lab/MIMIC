module fake_netlist_6_2045_n_1685 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_361, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1685);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1685;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_1664;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_527;
wire n_1207;
wire n_474;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_351),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_94),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_200),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_145),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_232),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_128),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_91),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_9),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_230),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_22),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_9),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_345),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_133),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_27),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_203),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_112),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_69),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_187),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_202),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_146),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_192),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_27),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_82),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_216),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_124),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_83),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_336),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_237),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_165),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_250),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_201),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_127),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_14),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_185),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_270),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_48),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_355),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_249),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_257),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_104),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_277),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_38),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_177),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_99),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_108),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_244),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_39),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_163),
.B(n_274),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_38),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_89),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_329),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_309),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_110),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_291),
.Y(n_421)
);

BUFx5_ASAP7_75t_L g422 ( 
.A(n_207),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_312),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_217),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_294),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_105),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_195),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_147),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_258),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_65),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_188),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_73),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_254),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_130),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_106),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_162),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_12),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_181),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_218),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_346),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_209),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_344),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_178),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_47),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_273),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_260),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_221),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_284),
.Y(n_448)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_20),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_33),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_213),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_90),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_161),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_48),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_136),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_348),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_324),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_63),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_44),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_358),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_45),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_263),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_304),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_164),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_142),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_226),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_349),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_68),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_60),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_321),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_340),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_88),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_220),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_137),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_148),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_158),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_211),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_272),
.B(n_305),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_129),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_55),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_228),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_97),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_134),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_15),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_240),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_229),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_319),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_208),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_153),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_333),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_316),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_343),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_40),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_212),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_126),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_117),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_172),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_215),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_169),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_111),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_17),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_17),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_361),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_184),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_198),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_248),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_292),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_323),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_120),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_16),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_7),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_118),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_261),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_199),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_363),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_266),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_58),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_53),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_239),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_101),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_57),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_66),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_10),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_114),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_233),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_342),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_241),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_26),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_77),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_0),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_243),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_42),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_338),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_23),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_22),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_14),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_320),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_341),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_356),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_71),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_326),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_186),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_75),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_194),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_42),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_50),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_285),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_26),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_150),
.Y(n_549)
);

BUFx5_ASAP7_75t_L g550 ( 
.A(n_311),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_317),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_0),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_337),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_39),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_251),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_157),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_113),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_189),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_268),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_282),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_13),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_271),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_359),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_330),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_152),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_196),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_55),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_279),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_7),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_50),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_52),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_286),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_132),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_131),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_160),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_331),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_252),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_60),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_167),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_302),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_328),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_287),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_298),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_155),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_235),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_144),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_52),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_191),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_109),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_8),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_327),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_154),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_19),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_86),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_98),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_179),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_204),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_238),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_590),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_428),
.B(n_1),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_449),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_399),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_449),
.Y(n_603)
);

NOR2x1_ASAP7_75t_L g604 ( 
.A(n_495),
.B(n_62),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_449),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_444),
.B(n_1),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_399),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_449),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_491),
.B(n_2),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_444),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_449),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_590),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_399),
.Y(n_613)
);

BUFx12f_ASAP7_75t_L g614 ( 
.A(n_420),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_511),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_399),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_379),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_420),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_379),
.Y(n_620)
);

CKINVDCx6p67_ASAP7_75t_R g621 ( 
.A(n_593),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_371),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_423),
.B(n_3),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_380),
.A2(n_67),
.B(n_64),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_374),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_379),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_491),
.B(n_4),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_373),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_381),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_432),
.B(n_5),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_381),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_449),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_422),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_501),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_422),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_515),
.B(n_5),
.Y(n_636)
);

BUFx12f_ASAP7_75t_L g637 ( 
.A(n_398),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_381),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_591),
.B(n_6),
.Y(n_639)
);

OA21x2_ASAP7_75t_L g640 ( 
.A1(n_369),
.A2(n_6),
.B(n_8),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_451),
.B(n_10),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_487),
.B(n_11),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_402),
.B(n_11),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_364),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_403),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_406),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_442),
.B(n_16),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_403),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_401),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_430),
.B(n_18),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_422),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_403),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_561),
.B(n_18),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_422),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_533),
.B(n_19),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_570),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_377),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_422),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_436),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_386),
.Y(n_660)
);

BUFx12f_ASAP7_75t_L g661 ( 
.A(n_407),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_436),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_437),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_436),
.Y(n_664)
);

BUFx8_ASAP7_75t_SL g665 ( 
.A(n_459),
.Y(n_665)
);

AOI22x1_ASAP7_75t_SL g666 ( 
.A1(n_461),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_422),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_414),
.B(n_24),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_450),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_454),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_412),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_480),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_482),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_482),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_469),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_550),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_493),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_521),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_592),
.B(n_25),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_494),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_487),
.B(n_28),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_494),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_534),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_567),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_382),
.B(n_28),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_484),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_569),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_502),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_494),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_537),
.Y(n_692)
);

BUFx12f_ASAP7_75t_L g693 ( 
.A(n_510),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_370),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_365),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_517),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_400),
.B(n_29),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_523),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_SL g699 ( 
.A1(n_552),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_528),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_438),
.B(n_30),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_532),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_368),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_453),
.B(n_31),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_535),
.Y(n_705)
);

BUFx12f_ASAP7_75t_L g706 ( 
.A(n_536),
.Y(n_706)
);

BUFx8_ASAP7_75t_L g707 ( 
.A(n_537),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_545),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_378),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_550),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_537),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_546),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_384),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_550),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_548),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_563),
.Y(n_716)
);

BUFx12f_ASAP7_75t_L g717 ( 
.A(n_554),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_571),
.B(n_32),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_578),
.B(n_32),
.Y(n_719)
);

BUFx8_ASAP7_75t_SL g720 ( 
.A(n_587),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_513),
.B(n_33),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_563),
.Y(n_722)
);

OA21x2_ASAP7_75t_L g723 ( 
.A1(n_387),
.A2(n_34),
.B(n_35),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_388),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_372),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_389),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_560),
.B(n_34),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_375),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_563),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_589),
.B(n_35),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_588),
.Y(n_731)
);

OAI21x1_ASAP7_75t_L g732 ( 
.A1(n_574),
.A2(n_72),
.B(n_70),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_589),
.B(n_36),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_588),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_392),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_376),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_367),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_588),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_395),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_396),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_366),
.B(n_36),
.Y(n_741)
);

INVxp33_ASAP7_75t_SL g742 ( 
.A(n_383),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_397),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_405),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_391),
.Y(n_745)
);

OAI22x1_ASAP7_75t_SL g746 ( 
.A1(n_394),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_550),
.Y(n_747)
);

BUFx8_ASAP7_75t_SL g748 ( 
.A(n_418),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_550),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_550),
.B(n_37),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_410),
.Y(n_751)
);

BUFx12f_ASAP7_75t_L g752 ( 
.A(n_385),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_417),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_390),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_419),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_408),
.B(n_41),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_424),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_748),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_703),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_617),
.Y(n_760)
);

CKINVDCx6p67_ASAP7_75t_R g761 ( 
.A(n_614),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_617),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_707),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_617),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_620),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_728),
.B(n_425),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_620),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_649),
.Y(n_768)
);

AND3x2_ASAP7_75t_L g769 ( 
.A(n_623),
.B(n_435),
.C(n_434),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_620),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_665),
.Y(n_771)
);

AOI21x1_ASAP7_75t_L g772 ( 
.A1(n_632),
.A2(n_446),
.B(n_445),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_725),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_752),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_599),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_720),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_626),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_737),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_676),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_626),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_R g781 ( 
.A(n_698),
.B(n_564),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_742),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_745),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_612),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_626),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_R g786 ( 
.A(n_698),
.B(n_582),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_644),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_R g788 ( 
.A(n_628),
.B(n_43),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_L g789 ( 
.A(n_702),
.B(n_447),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_700),
.B(n_708),
.Y(n_790)
);

BUFx10_ASAP7_75t_L g791 ( 
.A(n_618),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_638),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_R g793 ( 
.A(n_705),
.B(n_43),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_754),
.B(n_452),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_695),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_736),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_754),
.B(n_455),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_601),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_638),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_637),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_638),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_661),
.Y(n_802)
);

CKINVDCx16_ASAP7_75t_R g803 ( 
.A(n_671),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_693),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_712),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_621),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_603),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_605),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_645),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_645),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_706),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_645),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_717),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_630),
.B(n_741),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_608),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_636),
.B(n_470),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_648),
.Y(n_817)
);

XNOR2xp5_ASAP7_75t_L g818 ( 
.A(n_699),
.B(n_44),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_648),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_754),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_R g821 ( 
.A(n_715),
.B(n_393),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_715),
.B(n_507),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_611),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_622),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_619),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_707),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_669),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_688),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_690),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_648),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_659),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_696),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_739),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_659),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_740),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_659),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_664),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_610),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_609),
.B(n_45),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_629),
.B(n_456),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_625),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_664),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_751),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_744),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_R g845 ( 
.A(n_735),
.B(n_404),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_744),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_744),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_757),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_602),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_650),
.Y(n_850)
);

CKINVDCx16_ASAP7_75t_R g851 ( 
.A(n_636),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_R g852 ( 
.A(n_730),
.B(n_409),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_757),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_R g854 ( 
.A(n_694),
.B(n_411),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_664),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_675),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_724),
.B(n_549),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_694),
.B(n_415),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_757),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_629),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_652),
.Y(n_861)
);

AO221x1_ASAP7_75t_L g862 ( 
.A1(n_779),
.A2(n_646),
.B1(n_472),
.B2(n_475),
.C(n_466),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_SL g863 ( 
.A(n_850),
.B(n_655),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_849),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_841),
.B(n_718),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_838),
.B(n_639),
.Y(n_866)
);

NAND2xp33_ASAP7_75t_L g867 ( 
.A(n_852),
.B(n_627),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_849),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_857),
.B(n_822),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_827),
.B(n_639),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_798),
.B(n_633),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_814),
.B(n_631),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_839),
.A2(n_606),
.B1(n_647),
.B2(n_687),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_844),
.Y(n_874)
);

INVx4_ASAP7_75t_SL g875 ( 
.A(n_763),
.Y(n_875)
);

NOR3xp33_ASAP7_75t_L g876 ( 
.A(n_851),
.B(n_641),
.C(n_756),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_835),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_791),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_L g879 ( 
.A(n_852),
.B(n_643),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_790),
.B(n_833),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_798),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_843),
.A2(n_668),
.B1(n_682),
.B2(n_642),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_846),
.B(n_847),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_762),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_848),
.B(n_631),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_853),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_807),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_828),
.B(n_647),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_789),
.B(n_600),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_807),
.B(n_635),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_799),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_829),
.B(n_680),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_859),
.B(n_631),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_832),
.B(n_719),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_808),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_785),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_808),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_781),
.B(n_600),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_766),
.B(n_662),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_816),
.B(n_662),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_785),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_L g902 ( 
.A(n_821),
.B(n_653),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_837),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_759),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_837),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_781),
.B(n_687),
.Y(n_906)
);

OA21x2_ASAP7_75t_L g907 ( 
.A1(n_772),
.A2(n_732),
.B(n_624),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_815),
.B(n_662),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_773),
.B(n_733),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_815),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_840),
.B(n_750),
.C(n_701),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_L g912 ( 
.A(n_769),
.B(n_721),
.C(n_697),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_823),
.B(n_760),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_823),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_786),
.B(n_704),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_764),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_765),
.B(n_670),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_825),
.B(n_755),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_787),
.B(n_727),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_768),
.B(n_673),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_786),
.B(n_704),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_791),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_767),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_796),
.B(n_652),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_770),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_860),
.B(n_729),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_777),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_780),
.B(n_670),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_792),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_803),
.B(n_615),
.C(n_663),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_861),
.B(n_729),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_788),
.B(n_713),
.C(n_709),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_854),
.B(n_709),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_801),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_782),
.B(n_734),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_809),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_854),
.B(n_416),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_810),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_812),
.B(n_651),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_788),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_817),
.B(n_670),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_819),
.B(n_674),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_830),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_820),
.B(n_734),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_SL g945 ( 
.A(n_824),
.B(n_579),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_831),
.B(n_674),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_794),
.A2(n_723),
.B(n_640),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_834),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_836),
.B(n_674),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_842),
.B(n_713),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_855),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_858),
.B(n_726),
.Y(n_952)
);

AND2x2_ASAP7_75t_SL g953 ( 
.A(n_775),
.B(n_640),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_856),
.B(n_726),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_919),
.B(n_821),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_892),
.B(n_795),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_933),
.B(n_858),
.Y(n_957)
);

O2A1O1Ixp5_ASAP7_75t_L g958 ( 
.A1(n_947),
.A2(n_753),
.B(n_743),
.C(n_658),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_878),
.B(n_784),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_939),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_918),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_940),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_939),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_913),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_864),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_866),
.B(n_869),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_909),
.B(n_805),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_868),
.Y(n_968)
);

NAND2xp33_ASAP7_75t_L g969 ( 
.A(n_952),
.B(n_873),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_872),
.A2(n_613),
.B(n_413),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_884),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_889),
.B(n_657),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_903),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_910),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_889),
.B(n_845),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_916),
.B(n_679),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_877),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_891),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_881),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_925),
.B(n_660),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_887),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_902),
.B(n_911),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_903),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_870),
.B(n_845),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_947),
.A2(n_723),
.B(n_604),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_894),
.B(n_778),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_895),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_897),
.Y(n_988)
);

NOR2x2_ASAP7_75t_L g989 ( 
.A(n_945),
.B(n_746),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_874),
.B(n_826),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_888),
.B(n_783),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_922),
.Y(n_992)
);

NOR2x2_ASAP7_75t_L g993 ( 
.A(n_945),
.B(n_793),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_914),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_SL g995 ( 
.A1(n_923),
.A2(n_483),
.B(n_488),
.C(n_463),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_911),
.B(n_797),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_877),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_874),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_865),
.B(n_497),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_924),
.B(n_504),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_953),
.A2(n_509),
.B1(n_520),
.B2(n_519),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_886),
.B(n_763),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_927),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_871),
.B(n_654),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_901),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_905),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_912),
.A2(n_525),
.B1(n_531),
.B2(n_529),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_929),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_934),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_886),
.B(n_774),
.Y(n_1010)
);

AND3x1_ASAP7_75t_L g1011 ( 
.A(n_930),
.B(n_793),
.C(n_818),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_912),
.A2(n_862),
.B1(n_863),
.B2(n_867),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_926),
.B(n_931),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_906),
.B(n_539),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_923),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_943),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_938),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_903),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_915),
.B(n_776),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_936),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_908),
.B(n_743),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_921),
.B(n_541),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_SL g1023 ( 
.A(n_882),
.B(n_806),
.C(n_802),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_879),
.B(n_547),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_951),
.Y(n_1025)
);

AND3x2_ASAP7_75t_SL g1026 ( 
.A(n_876),
.B(n_666),
.C(n_771),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_880),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_920),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_932),
.A2(n_753),
.B1(n_478),
.B2(n_559),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_871),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_883),
.B(n_556),
.Y(n_1031)
);

O2A1O1Ixp5_ASAP7_75t_L g1032 ( 
.A1(n_898),
.A2(n_677),
.B(n_710),
.C(n_667),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_890),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_935),
.B(n_761),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_936),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_936),
.B(n_584),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_948),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_948),
.B(n_596),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_890),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_948),
.B(n_597),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_904),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_932),
.A2(n_747),
.B(n_714),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_950),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_885),
.B(n_421),
.Y(n_1044)
);

NOR2x2_ASAP7_75t_L g1045 ( 
.A(n_875),
.B(n_666),
.Y(n_1045)
);

BUFx4f_ASAP7_75t_L g1046 ( 
.A(n_907),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_907),
.A2(n_749),
.B1(n_672),
.B2(n_678),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_944),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_896),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_896),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_900),
.B(n_813),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_937),
.B(n_800),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_875),
.B(n_804),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_969),
.A2(n_893),
.B1(n_954),
.B2(n_427),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_998),
.B(n_875),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_974),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_982),
.A2(n_429),
.B1(n_431),
.B2(n_426),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_999),
.A2(n_917),
.B(n_941),
.C(n_928),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_981),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_998),
.B(n_896),
.Y(n_1060)
);

CKINVDCx16_ASAP7_75t_R g1061 ( 
.A(n_1053),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_960),
.B(n_433),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1046),
.A2(n_946),
.B(n_942),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1028),
.B(n_811),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_997),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_980),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1001),
.A2(n_440),
.B(n_441),
.C(n_439),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_979),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_L g1069 ( 
.A(n_998),
.B(n_1019),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_956),
.B(n_758),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_1030),
.A2(n_949),
.B(n_899),
.C(n_672),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1012),
.A2(n_448),
.B1(n_457),
.B2(n_443),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_972),
.B(n_961),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_985),
.A2(n_460),
.B(n_462),
.C(n_458),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_973),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1046),
.A2(n_613),
.B(n_692),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1033),
.A2(n_678),
.B(n_683),
.C(n_660),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_985),
.A2(n_613),
.B(n_692),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_963),
.B(n_964),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_987),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1039),
.A2(n_692),
.B(n_607),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1024),
.A2(n_955),
.B1(n_1013),
.B2(n_957),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_1042),
.A2(n_685),
.B(n_686),
.C(n_683),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1043),
.B(n_464),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_962),
.B(n_685),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1004),
.A2(n_607),
.B(n_602),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_1020),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1031),
.B(n_465),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1048),
.B(n_467),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_1018),
.B(n_686),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_1020),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_973),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1041),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_972),
.B(n_689),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_966),
.A2(n_471),
.B1(n_473),
.B2(n_468),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_973),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_980),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1000),
.B(n_474),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_983),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_967),
.B(n_476),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_SL g1101 ( 
.A(n_1020),
.B(n_477),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_988),
.B(n_479),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_977),
.Y(n_1103)
);

OAI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_1007),
.A2(n_689),
.B(n_656),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1047),
.A2(n_558),
.B1(n_485),
.B2(n_486),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_996),
.A2(n_656),
.B(n_634),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_986),
.B(n_1027),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1042),
.A2(n_634),
.B(n_481),
.C(n_557),
.Y(n_1108)
);

INVx8_ASAP7_75t_L g1109 ( 
.A(n_959),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_958),
.A2(n_565),
.B(n_490),
.C(n_492),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_SL g1111 ( 
.A1(n_995),
.A2(n_566),
.B(n_496),
.C(n_498),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1014),
.A2(n_572),
.B1(n_499),
.B2(n_500),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_977),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1034),
.B(n_489),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1003),
.B(n_74),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_994),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1004),
.A2(n_607),
.B(n_602),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_984),
.B(n_503),
.Y(n_1118)
);

CKINVDCx8_ASAP7_75t_R g1119 ( 
.A(n_959),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_983),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_976),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1022),
.A2(n_573),
.B(n_506),
.C(n_508),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_975),
.A2(n_576),
.B(n_512),
.C(n_514),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_SL g1124 ( 
.A(n_1023),
.B(n_991),
.C(n_1052),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1008),
.A2(n_577),
.B1(n_516),
.B2(n_522),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1015),
.A2(n_581),
.B1(n_524),
.B2(n_526),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_992),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_1011),
.B(n_1029),
.C(n_1016),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_992),
.B(n_505),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_L g1130 ( 
.A(n_1010),
.B(n_538),
.C(n_527),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1009),
.A2(n_586),
.B1(n_542),
.B2(n_543),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_993),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_976),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_965),
.B(n_968),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1044),
.A2(n_1037),
.B(n_1035),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1032),
.A2(n_616),
.B(n_675),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1025),
.A2(n_544),
.B(n_540),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_990),
.B(n_551),
.Y(n_1138)
);

CKINVDCx14_ASAP7_75t_R g1139 ( 
.A(n_1065),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1103),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1113),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_1109),
.B(n_959),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1093),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1128),
.A2(n_1029),
.B(n_1036),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1068),
.Y(n_1145)
);

AO21x2_ASAP7_75t_L g1146 ( 
.A1(n_1110),
.A2(n_1040),
.B(n_1038),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1132),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_1127),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1080),
.Y(n_1149)
);

AO21x1_ASAP7_75t_L g1150 ( 
.A1(n_1082),
.A2(n_970),
.B(n_971),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1074),
.A2(n_978),
.B(n_1021),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1135),
.A2(n_1006),
.B(n_1005),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_1109),
.B(n_1115),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1079),
.A2(n_1108),
.B(n_1078),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1116),
.Y(n_1155)
);

BUFx2_ASAP7_75t_SL g1156 ( 
.A(n_1087),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1073),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1073),
.Y(n_1158)
);

AOI22x1_ASAP7_75t_L g1159 ( 
.A1(n_1063),
.A2(n_1017),
.B1(n_1050),
.B2(n_1049),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1107),
.B(n_983),
.Y(n_1160)
);

BUFx4f_ASAP7_75t_L g1161 ( 
.A(n_1092),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1087),
.Y(n_1162)
);

BUFx12f_ASAP7_75t_L g1163 ( 
.A(n_1094),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1067),
.A2(n_1021),
.B(n_1011),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1087),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1134),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_1094),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1056),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1092),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1069),
.B(n_1002),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1092),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1059),
.Y(n_1172)
);

CKINVDCx6p67_ASAP7_75t_R g1173 ( 
.A(n_1061),
.Y(n_1173)
);

AO21x1_ASAP7_75t_L g1174 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1026),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_1091),
.B(n_616),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1072),
.A2(n_555),
.B(n_553),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1096),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1062),
.A2(n_568),
.B(n_562),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1091),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1054),
.A2(n_580),
.B(n_575),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1137),
.A2(n_585),
.B(n_583),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1066),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_1118),
.A2(n_46),
.B(n_47),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1097),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1121),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1096),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1085),
.Y(n_1187)
);

BUFx2_ASAP7_75t_SL g1188 ( 
.A(n_1096),
.Y(n_1188)
);

NAND2x1_ASAP7_75t_L g1189 ( 
.A(n_1099),
.B(n_1075),
.Y(n_1189)
);

AO21x2_ASAP7_75t_L g1190 ( 
.A1(n_1106),
.A2(n_595),
.B(n_594),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1099),
.B(n_616),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_1098),
.A2(n_598),
.B(n_78),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1133),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1120),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1136),
.A2(n_79),
.B(n_76),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1077),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_SL g1197 ( 
.A1(n_1058),
.A2(n_81),
.B(n_80),
.Y(n_1197)
);

AO21x2_ASAP7_75t_L g1198 ( 
.A1(n_1088),
.A2(n_85),
.B(n_84),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1099),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1083),
.Y(n_1200)
);

INVx3_ASAP7_75t_SL g1201 ( 
.A(n_1064),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1084),
.B(n_46),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1115),
.Y(n_1203)
);

CKINVDCx12_ASAP7_75t_R g1204 ( 
.A(n_1114),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1119),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1104),
.Y(n_1206)
);

OR3x4_ASAP7_75t_SL g1207 ( 
.A(n_1124),
.B(n_989),
.C(n_1045),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1086),
.A2(n_1117),
.B(n_1076),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1055),
.B(n_675),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1071),
.A2(n_245),
.B(n_362),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1090),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1089),
.B(n_87),
.Y(n_1212)
);

BUFx12f_ASAP7_75t_L g1213 ( 
.A(n_1060),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1102),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1123),
.A2(n_246),
.B(n_360),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1202),
.A2(n_1138),
.B1(n_1130),
.B2(n_1070),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1187),
.B(n_1095),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_SL g1218 ( 
.A1(n_1202),
.A2(n_1105),
.B1(n_1112),
.B2(n_1131),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1145),
.Y(n_1219)
);

INVx8_ASAP7_75t_L g1220 ( 
.A(n_1163),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1149),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1183),
.A2(n_1057),
.B1(n_1129),
.B2(n_1101),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1150),
.A2(n_1081),
.B(n_1126),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1155),
.Y(n_1224)
);

AO21x2_ASAP7_75t_L g1225 ( 
.A1(n_1154),
.A2(n_1122),
.B(n_1111),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1172),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1168),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1143),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1152),
.A2(n_1125),
.B(n_242),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1153),
.B(n_92),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1159),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1187),
.B(n_49),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1208),
.A2(n_247),
.B(n_357),
.Y(n_1233)
);

BUFx8_ASAP7_75t_SL g1234 ( 
.A(n_1148),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1140),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1154),
.A2(n_738),
.B(n_731),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1151),
.A2(n_236),
.B(n_353),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_SL g1238 ( 
.A1(n_1197),
.A2(n_234),
.B(n_352),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1166),
.A2(n_1203),
.B1(n_1214),
.B2(n_1160),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1147),
.B(n_49),
.Y(n_1240)
);

BUFx4f_ASAP7_75t_SL g1241 ( 
.A(n_1173),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1161),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1200),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1151),
.A2(n_231),
.B(n_350),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1179),
.B(n_681),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1174),
.A2(n_738),
.B1(n_731),
.B2(n_722),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1201),
.A2(n_738),
.B1(n_731),
.B2(n_722),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1182),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1184),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1167),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1162),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1201),
.A2(n_722),
.B1(n_716),
.B2(n_711),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1185),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1193),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1141),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1206),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1144),
.A2(n_716),
.B1(n_711),
.B2(n_691),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1162),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1161),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1139),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1153),
.B(n_93),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1177),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1160),
.A2(n_716),
.B1(n_711),
.B2(n_691),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1141),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1165),
.Y(n_1265)
);

AOI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1212),
.A2(n_691),
.B(n_684),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1179),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1177),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1194),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1144),
.A2(n_684),
.B1(n_681),
.B2(n_54),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1139),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1191),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1199),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1195),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1140),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1153),
.A2(n_684),
.B1(n_681),
.B2(n_54),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1191),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1186),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1196),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1186),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1210),
.A2(n_51),
.B(n_53),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1199),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1147),
.B(n_51),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1189),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1175),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1207),
.Y(n_1286)
);

AO21x1_ASAP7_75t_L g1287 ( 
.A1(n_1212),
.A2(n_56),
.B(n_57),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1175),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1164),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1157),
.Y(n_1290)
);

BUFx2_ASAP7_75t_SL g1291 ( 
.A(n_1165),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1158),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_SL g1293 ( 
.A(n_1242),
.B(n_1211),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1217),
.B(n_1204),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1242),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_R g1296 ( 
.A(n_1228),
.B(n_1213),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1234),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1219),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1231),
.A2(n_1192),
.A3(n_1190),
.B(n_1181),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1255),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1255),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1264),
.B(n_1164),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1242),
.Y(n_1303)
);

NOR2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1275),
.B(n_1205),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1264),
.B(n_1169),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1275),
.Y(n_1306)
);

OAI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1216),
.A2(n_1176),
.B(n_1178),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1217),
.A2(n_1181),
.B1(n_1176),
.B2(n_1180),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1273),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1243),
.B(n_1178),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1226),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1273),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1271),
.Y(n_1313)
);

AND2x4_ASAP7_75t_SL g1314 ( 
.A(n_1242),
.B(n_1142),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1231),
.A2(n_1192),
.A3(n_1190),
.B(n_1146),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1224),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1243),
.B(n_1146),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1256),
.B(n_1170),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1250),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1259),
.Y(n_1320)
);

OR2x6_ASAP7_75t_L g1321 ( 
.A(n_1230),
.B(n_1156),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1290),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1227),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1256),
.B(n_1170),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_R g1325 ( 
.A(n_1260),
.B(n_1205),
.Y(n_1325)
);

CKINVDCx16_ASAP7_75t_R g1326 ( 
.A(n_1271),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1274),
.A2(n_1287),
.A3(n_1279),
.B(n_1239),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1240),
.B(n_1171),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1221),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1230),
.A2(n_1180),
.B1(n_1207),
.B2(n_1198),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1216),
.A2(n_1142),
.B1(n_1198),
.B2(n_1188),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1248),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1259),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1292),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1259),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1283),
.B(n_1142),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1259),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_R g1338 ( 
.A(n_1261),
.B(n_1215),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_SL g1339 ( 
.A(n_1235),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1250),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1274),
.A2(n_1209),
.A3(n_61),
.B(n_59),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1241),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1220),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_SL g1344 ( 
.A(n_1218),
.B(n_1209),
.C(n_61),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1257),
.B(n_95),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1249),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1229),
.A2(n_1266),
.B(n_1223),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1241),
.Y(n_1348)
);

NAND2xp33_ASAP7_75t_R g1349 ( 
.A(n_1261),
.B(n_96),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1262),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1253),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1268),
.B(n_1282),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1220),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1232),
.B(n_100),
.Y(n_1354)
);

INVx4_ASAP7_75t_SL g1355 ( 
.A(n_1251),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1254),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1278),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1269),
.B(n_102),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1280),
.B(n_1267),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1251),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1258),
.B(n_103),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1220),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1272),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1258),
.B(n_107),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1277),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1289),
.B(n_115),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1298),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1302),
.B(n_1289),
.Y(n_1368)
);

INVx4_ASAP7_75t_SL g1369 ( 
.A(n_1341),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1305),
.B(n_1336),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1328),
.B(n_1222),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1316),
.Y(n_1372)
);

OAI33xp33_ASAP7_75t_L g1373 ( 
.A1(n_1307),
.A2(n_1276),
.A3(n_1252),
.B1(n_1247),
.B2(n_1263),
.B3(n_1284),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1311),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1301),
.B(n_1237),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1366),
.A2(n_1237),
.B1(n_1244),
.B2(n_1270),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1332),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1354),
.B(n_1222),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1307),
.A2(n_1270),
.B1(n_1276),
.B2(n_1246),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1300),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1308),
.A2(n_1246),
.B(n_1257),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1317),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1310),
.B(n_1318),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1310),
.B(n_1244),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1346),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1294),
.B(n_1285),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1318),
.B(n_1324),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1323),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1309),
.B(n_1225),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1352),
.B(n_1288),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1352),
.B(n_1265),
.Y(n_1391)
);

NOR2x1_ASAP7_75t_SL g1392 ( 
.A(n_1344),
.B(n_1225),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1350),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1312),
.B(n_1236),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1344),
.A2(n_1286),
.B1(n_1238),
.B2(n_1281),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1357),
.B(n_1265),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1306),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1329),
.B(n_1245),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1351),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1321),
.A2(n_1252),
.B1(n_1247),
.B2(n_1251),
.Y(n_1400)
);

OR2x2_ASAP7_75t_SL g1401 ( 
.A(n_1326),
.B(n_1281),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1356),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1321),
.B(n_1233),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1317),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1321),
.B(n_1245),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1324),
.B(n_1236),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1360),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1331),
.A2(n_1236),
.B(n_1281),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1322),
.B(n_1291),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1314),
.B(n_116),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1345),
.A2(n_1263),
.B(n_121),
.Y(n_1411)
);

INVxp67_ASAP7_75t_L g1412 ( 
.A(n_1334),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1327),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1359),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1363),
.B(n_1286),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1330),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1327),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1360),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1304),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1349),
.A2(n_125),
.B1(n_135),
.B2(n_138),
.Y(n_1420)
);

NAND2xp33_ASAP7_75t_R g1421 ( 
.A(n_1345),
.B(n_139),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1365),
.B(n_140),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1313),
.B(n_141),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1327),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1358),
.B(n_143),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1303),
.B(n_149),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1319),
.A2(n_151),
.B1(n_156),
.B2(n_159),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1293),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1331),
.B(n_166),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1303),
.B(n_1320),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1341),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1320),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1341),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1355),
.B(n_168),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1333),
.B(n_1335),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1299),
.B(n_170),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1315),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1315),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1333),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1343),
.B(n_171),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1315),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1335),
.B(n_1361),
.Y(n_1442)
);

AND2x2_ASAP7_75t_SL g1443 ( 
.A(n_1408),
.B(n_1379),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1382),
.B(n_1299),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1367),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1374),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1381),
.B(n_1361),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1388),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1414),
.B(n_1299),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1382),
.B(n_1404),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1370),
.B(n_1325),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1380),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1393),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1399),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1389),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1404),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1402),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1407),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1412),
.B(n_1364),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1377),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1403),
.B(n_1355),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1375),
.B(n_1347),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1412),
.Y(n_1463)
);

NAND2x1_ASAP7_75t_SL g1464 ( 
.A(n_1403),
.B(n_1378),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1409),
.Y(n_1465)
);

AND2x4_ASAP7_75t_SL g1466 ( 
.A(n_1396),
.B(n_1295),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1385),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1394),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1438),
.Y(n_1469)
);

AOI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1416),
.A2(n_1364),
.B1(n_1340),
.B2(n_1353),
.C(n_1362),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1431),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1441),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1433),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1372),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1383),
.B(n_1387),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1413),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1371),
.B(n_1347),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1417),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1384),
.B(n_1295),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1383),
.B(n_1295),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1384),
.B(n_1337),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1417),
.B(n_1337),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1424),
.B(n_1337),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1387),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1408),
.B(n_173),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1437),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1408),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1437),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1369),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1369),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1406),
.B(n_174),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1369),
.B(n_1338),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1406),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1401),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1436),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1386),
.B(n_1429),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1405),
.B(n_1342),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1390),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1432),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1368),
.B(n_1348),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1439),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1430),
.B(n_1435),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1461),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1461),
.B(n_1428),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1477),
.B(n_1392),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1450),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1477),
.B(n_1376),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1450),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1484),
.B(n_1376),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1494),
.B(n_1415),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1494),
.B(n_1391),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1468),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1479),
.B(n_1381),
.Y(n_1513)
);

NAND2x1p5_ASAP7_75t_L g1514 ( 
.A(n_1492),
.B(n_1407),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1479),
.B(n_1395),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1456),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1447),
.A2(n_1421),
.B1(n_1379),
.B2(n_1416),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1471),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1481),
.B(n_1395),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1475),
.B(n_1428),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1451),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1481),
.B(n_1443),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1473),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1443),
.B(n_1442),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1476),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1493),
.B(n_1398),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1447),
.A2(n_1427),
.B1(n_1420),
.B2(n_1373),
.Y(n_1527)
);

AND2x2_ASAP7_75t_SL g1528 ( 
.A(n_1492),
.B(n_1421),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1463),
.B(n_1411),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1444),
.B(n_1397),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1444),
.B(n_1397),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1455),
.B(n_1423),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1445),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1476),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1502),
.B(n_1411),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1446),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1502),
.B(n_1419),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1422),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1465),
.B(n_1426),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1485),
.B(n_1400),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1469),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1470),
.A2(n_1373),
.B1(n_1425),
.B2(n_1400),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1533),
.Y(n_1543)
);

NAND2x2_ASAP7_75t_L g1544 ( 
.A(n_1503),
.B(n_1500),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1533),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1536),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1536),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1512),
.B(n_1453),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1449),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1511),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1518),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1517),
.A2(n_1461),
.B1(n_1495),
.B2(n_1491),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1518),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1506),
.B(n_1462),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1523),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1452),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1530),
.B(n_1497),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1508),
.B(n_1495),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1516),
.B(n_1448),
.Y(n_1561)
);

NOR2xp67_ASAP7_75t_L g1562 ( 
.A(n_1529),
.B(n_1458),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1511),
.Y(n_1563)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1564 ( 
.A1(n_1509),
.A2(n_1498),
.B(n_1490),
.C(n_1488),
.D(n_1486),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1523),
.Y(n_1565)
);

INVxp33_ASAP7_75t_L g1566 ( 
.A(n_1538),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1517),
.A2(n_1496),
.B1(n_1459),
.B2(n_1480),
.Y(n_1567)
);

OAI32xp33_ASAP7_75t_L g1568 ( 
.A1(n_1527),
.A2(n_1485),
.A3(n_1489),
.B1(n_1487),
.B2(n_1457),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1528),
.A2(n_1491),
.B1(n_1497),
.B2(n_1440),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1520),
.A2(n_1489),
.B1(n_1458),
.B2(n_1440),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1541),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1507),
.B(n_1478),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1531),
.B(n_1497),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1568),
.A2(n_1528),
.B(n_1504),
.Y(n_1574)
);

AO22x1_ASAP7_75t_L g1575 ( 
.A1(n_1566),
.A2(n_1510),
.B1(n_1521),
.B2(n_1531),
.Y(n_1575)
);

AOI31xp33_ASAP7_75t_L g1576 ( 
.A1(n_1569),
.A2(n_1514),
.A3(n_1510),
.B(n_1542),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1571),
.Y(n_1577)
);

NAND4xp25_ASAP7_75t_SL g1578 ( 
.A(n_1553),
.B(n_1507),
.C(n_1540),
.D(n_1522),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1543),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1558),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1545),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1544),
.A2(n_1503),
.B1(n_1514),
.B2(n_1540),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1564),
.A2(n_1535),
.B(n_1513),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1573),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1567),
.A2(n_1535),
.B1(n_1515),
.B2(n_1519),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1547),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1557),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1572),
.B(n_1513),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1567),
.A2(n_1519),
.B1(n_1515),
.B2(n_1537),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1570),
.A2(n_1503),
.B1(n_1514),
.B2(n_1522),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1551),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_L g1593 ( 
.A(n_1552),
.B(n_1539),
.C(n_1532),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1554),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1555),
.B(n_1505),
.Y(n_1595)
);

OAI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1552),
.A2(n_1464),
.B(n_1505),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1560),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1576),
.A2(n_1562),
.B(n_1548),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1593),
.B(n_1537),
.Y(n_1599)
);

AOI211x1_ASAP7_75t_L g1600 ( 
.A1(n_1574),
.A2(n_1548),
.B(n_1549),
.C(n_1561),
.Y(n_1600)
);

OAI32xp33_ASAP7_75t_L g1601 ( 
.A1(n_1584),
.A2(n_1549),
.A3(n_1561),
.B1(n_1565),
.B2(n_1556),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1579),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1586),
.A2(n_1524),
.B1(n_1550),
.B2(n_1563),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1591),
.A2(n_1467),
.B(n_1499),
.C(n_1501),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1586),
.A2(n_1524),
.B(n_1538),
.C(n_1539),
.Y(n_1605)
);

OAI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1596),
.A2(n_1532),
.B1(n_1526),
.B2(n_1559),
.C(n_1474),
.Y(n_1606)
);

OAI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1590),
.A2(n_1559),
.B1(n_1487),
.B2(n_1541),
.Y(n_1607)
);

OAI211xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1590),
.A2(n_1454),
.B(n_1460),
.C(n_1541),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1297),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1581),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1597),
.B(n_1526),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1588),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1583),
.A2(n_1434),
.B1(n_1482),
.B2(n_1466),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1587),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1589),
.B(n_1575),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1592),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1594),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

NAND4xp25_ASAP7_75t_SL g1620 ( 
.A(n_1598),
.B(n_1595),
.C(n_1577),
.D(n_1296),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1600),
.B(n_1454),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1617),
.B(n_1483),
.Y(n_1622)
);

NOR3x1_ASAP7_75t_L g1623 ( 
.A(n_1612),
.B(n_1339),
.C(n_1466),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

NOR3x1_ASAP7_75t_L g1625 ( 
.A(n_1606),
.B(n_1434),
.C(n_1458),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_L g1626 ( 
.A(n_1609),
.B(n_1410),
.C(n_1460),
.Y(n_1626)
);

AOI221x1_ASAP7_75t_L g1627 ( 
.A1(n_1607),
.A2(n_1541),
.B1(n_1482),
.B2(n_1483),
.C(n_1525),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1601),
.B(n_1410),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1615),
.B(n_1525),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1610),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1599),
.B(n_1534),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1628),
.B(n_1605),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1624),
.Y(n_1633)
);

OA22x2_ASAP7_75t_SL g1634 ( 
.A1(n_1630),
.A2(n_1603),
.B1(n_1618),
.B2(n_1619),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1629),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1626),
.B(n_1613),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1622),
.Y(n_1637)
);

AOI211xp5_ASAP7_75t_L g1638 ( 
.A1(n_1620),
.A2(n_1604),
.B(n_1616),
.C(n_1621),
.Y(n_1638)
);

OAI222xp33_ASAP7_75t_L g1639 ( 
.A1(n_1625),
.A2(n_1599),
.B1(n_1611),
.B2(n_1614),
.C1(n_1608),
.C2(n_1534),
.Y(n_1639)
);

AOI211x1_ASAP7_75t_L g1640 ( 
.A1(n_1627),
.A2(n_1478),
.B(n_1534),
.C(n_180),
.Y(n_1640)
);

NAND2xp33_ASAP7_75t_SL g1641 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1639),
.A2(n_1631),
.B1(n_1472),
.B2(n_1469),
.C(n_1418),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1633),
.Y(n_1643)
);

OAI321xp33_ASAP7_75t_L g1644 ( 
.A1(n_1638),
.A2(n_1634),
.A3(n_1635),
.B1(n_1636),
.B2(n_1637),
.C(n_1640),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1636),
.A2(n_1472),
.B1(n_1418),
.B2(n_1407),
.C(n_183),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1638),
.B(n_1407),
.C(n_1418),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1633),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1632),
.A2(n_1418),
.B1(n_176),
.B2(n_182),
.C(n_190),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1641),
.A2(n_175),
.B1(n_193),
.B2(n_197),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1648),
.A2(n_205),
.B1(n_206),
.B2(n_210),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1643),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1647),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1646),
.Y(n_1653)
);

AO22x1_ASAP7_75t_L g1654 ( 
.A1(n_1644),
.A2(n_214),
.B1(n_219),
.B2(n_222),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_R g1655 ( 
.A(n_1653),
.B(n_1645),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1652),
.B(n_1642),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_223),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1649),
.B(n_224),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1656),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1655),
.Y(n_1660)
);

OA22x2_ASAP7_75t_L g1661 ( 
.A1(n_1658),
.A2(n_1654),
.B1(n_1650),
.B2(n_253),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1657),
.B(n_225),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1660),
.A2(n_227),
.B1(n_255),
.B2(n_256),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1659),
.A2(n_259),
.B1(n_262),
.B2(n_264),
.C(n_265),
.Y(n_1664)
);

XOR2xp5_ASAP7_75t_L g1665 ( 
.A(n_1661),
.B(n_267),
.Y(n_1665)
);

OAI22x1_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1662),
.B1(n_275),
.B2(n_276),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1663),
.Y(n_1667)
);

AO22x2_ASAP7_75t_L g1668 ( 
.A1(n_1664),
.A2(n_347),
.B1(n_278),
.B2(n_280),
.Y(n_1668)
);

INVx3_ASAP7_75t_SL g1669 ( 
.A(n_1665),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1669),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1667),
.A2(n_269),
.B1(n_281),
.B2(n_283),
.Y(n_1671)
);

OAI22x1_ASAP7_75t_L g1672 ( 
.A1(n_1666),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_1672)
);

INVx3_ASAP7_75t_SL g1673 ( 
.A(n_1668),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1670),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1672),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1671),
.A2(n_297),
.B(n_299),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1673),
.A2(n_300),
.B1(n_301),
.B2(n_303),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1674),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1677),
.B(n_1676),
.Y(n_1679)
);

AOI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1675),
.A2(n_306),
.B(n_307),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1678),
.A2(n_1679),
.B1(n_1680),
.B2(n_314),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1678),
.A2(n_308),
.B1(n_313),
.B2(n_315),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1679),
.A2(n_318),
.B1(n_325),
.B2(n_332),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1681),
.B(n_334),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1682),
.B1(n_1683),
.B2(n_335),
.Y(n_1685)
);


endmodule