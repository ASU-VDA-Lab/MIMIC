module real_aes_8795_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g238 ( .A1(n_0), .A2(n_239), .B(n_242), .C(n_246), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_1), .B(n_230), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g113 ( .A1(n_2), .A2(n_7), .B1(n_114), .B2(n_118), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_3), .A2(n_30), .B1(n_103), .B2(n_108), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_4), .B(n_240), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_5), .A2(n_200), .B(n_270), .Y(n_269) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_6), .A2(n_232), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g187 ( .A(n_8), .Y(n_187) );
AND2x6_ASAP7_75t_L g205 ( .A(n_8), .B(n_185), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_8), .B(n_514), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_9), .A2(n_205), .B(n_207), .C(n_296), .Y(n_295) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_10), .A2(n_22), .B1(n_92), .B2(n_93), .Y(n_91) );
INVx1_ASAP7_75t_L g225 ( .A(n_11), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_12), .B(n_240), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_13), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_170) );
INVx1_ASAP7_75t_L g173 ( .A(n_13), .Y(n_173) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_14), .A2(n_24), .B1(n_92), .B2(n_96), .Y(n_95) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_15), .A2(n_72), .B1(n_123), .B2(n_130), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_16), .A2(n_207), .B(n_210), .C(n_218), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_17), .A2(n_207), .B(n_218), .C(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_18), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_19), .A2(n_200), .B(n_235), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_20), .A2(n_38), .B1(n_136), .B2(n_140), .Y(n_135) );
INVx2_ASAP7_75t_L g203 ( .A(n_21), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_23), .A2(n_258), .B(n_259), .C(n_263), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g178 ( .A1(n_24), .A2(n_41), .B1(n_53), .B2(n_179), .C(n_180), .Y(n_178) );
INVxp67_ASAP7_75t_L g181 ( .A(n_24), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_25), .A2(n_58), .B1(n_160), .B2(n_161), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_26), .B(n_312), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_27), .A2(n_56), .B1(n_145), .B2(n_148), .Y(n_144) );
AOI22xp33_ASAP7_75t_SL g152 ( .A1(n_28), .A2(n_42), .B1(n_153), .B2(n_156), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_29), .B(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_31), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_32), .B(n_240), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_33), .B(n_200), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_34), .A2(n_258), .B(n_263), .C(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g243 ( .A(n_35), .Y(n_243) );
INVx1_ASAP7_75t_L g286 ( .A(n_36), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_37), .B(n_200), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_39), .Y(n_227) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_40), .Y(n_172) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_41), .A2(n_63), .B1(n_92), .B2(n_96), .Y(n_99) );
INVxp67_ASAP7_75t_L g182 ( .A(n_41), .Y(n_182) );
INVx1_ASAP7_75t_L g185 ( .A(n_43), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_44), .B(n_200), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_45), .B(n_230), .Y(n_277) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_46), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_46), .A2(n_217), .B(n_273), .C(n_275), .Y(n_272) );
OAI22xp5_ASAP7_75t_SL g165 ( .A1(n_47), .A2(n_166), .B1(n_167), .B2(n_168), .Y(n_165) );
INVx1_ASAP7_75t_L g168 ( .A(n_47), .Y(n_168) );
INVx1_ASAP7_75t_L g224 ( .A(n_48), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_49), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_50), .B(n_240), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_51), .B(n_241), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_52), .A2(n_82), .B1(n_83), .B2(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_52), .Y(n_522) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_53), .A2(n_68), .B1(n_92), .B2(n_93), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_54), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_55), .B(n_212), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_57), .A2(n_207), .B(n_263), .C(n_326), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_59), .Y(n_271) );
INVx1_ASAP7_75t_L g81 ( .A(n_60), .Y(n_81) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_61), .B(n_215), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_62), .Y(n_265) );
INVx2_ASAP7_75t_L g222 ( .A(n_64), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_65), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_66), .B(n_245), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_66), .A2(n_82), .B1(n_83), .B2(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_66), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_67), .B(n_200), .Y(n_256) );
INVx1_ASAP7_75t_L g260 ( .A(n_69), .Y(n_260) );
INVxp67_ASAP7_75t_L g276 ( .A(n_70), .Y(n_276) );
INVx1_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
INVx1_ASAP7_75t_L g94 ( .A(n_71), .Y(n_94) );
INVx1_ASAP7_75t_L g293 ( .A(n_73), .Y(n_293) );
INVx1_ASAP7_75t_L g327 ( .A(n_74), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_75), .Y(n_87) );
AND2x2_ASAP7_75t_L g288 ( .A(n_76), .B(n_221), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_175), .B1(n_188), .B2(n_503), .C(n_508), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_164), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_82), .B1(n_83), .B2(n_163), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_80), .Y(n_163) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND2xp5_ASAP7_75t_SL g84 ( .A(n_85), .B(n_133), .Y(n_84) );
NOR2xp33_ASAP7_75t_L g85 ( .A(n_86), .B(n_112), .Y(n_85) );
OAI21xp5_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_88), .B(n_102), .Y(n_86) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x6_ASAP7_75t_L g89 ( .A(n_90), .B(n_97), .Y(n_89) );
AND2x4_ASAP7_75t_L g109 ( .A(n_90), .B(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_95), .Y(n_90) );
AND2x2_ASAP7_75t_L g107 ( .A(n_91), .B(n_99), .Y(n_107) );
INVx2_ASAP7_75t_L g129 ( .A(n_91), .Y(n_129) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_94), .Y(n_96) );
INVx2_ASAP7_75t_L g117 ( .A(n_95), .Y(n_117) );
INVx1_ASAP7_75t_L g121 ( .A(n_95), .Y(n_121) );
OR2x2_ASAP7_75t_L g128 ( .A(n_95), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g132 ( .A(n_95), .B(n_129), .Y(n_132) );
AND2x2_ASAP7_75t_L g147 ( .A(n_97), .B(n_139), .Y(n_147) );
AND2x6_ASAP7_75t_L g150 ( .A(n_97), .B(n_127), .Y(n_150) );
AND2x4_ASAP7_75t_L g155 ( .A(n_97), .B(n_132), .Y(n_155) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
AND2x2_ASAP7_75t_L g126 ( .A(n_98), .B(n_101), .Y(n_126) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g138 ( .A(n_99), .B(n_111), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_99), .B(n_101), .Y(n_143) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g106 ( .A(n_101), .Y(n_106) );
INVx1_ASAP7_75t_L g111 ( .A(n_101), .Y(n_111) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g116 ( .A(n_106), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g115 ( .A(n_107), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g119 ( .A(n_107), .B(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_122), .Y(n_112) );
BUFx4f_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g139 ( .A(n_117), .B(n_129), .Y(n_139) );
BUFx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x6_ASAP7_75t_L g162 ( .A(n_121), .B(n_143), .Y(n_162) );
INVx5_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x6_ASAP7_75t_L g131 ( .A(n_126), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g160 ( .A(n_126), .B(n_139), .Y(n_160) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx4f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g158 ( .A(n_132), .B(n_138), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_151), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_144), .Y(n_134) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x4_ASAP7_75t_L g141 ( .A(n_139), .B(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx5_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
INVx11_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_159), .Y(n_151) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx8_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx6_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_169), .B1(n_170), .B2(n_174), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_165), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_166), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
AND3x1_ASAP7_75t_SL g177 ( .A(n_178), .B(n_183), .C(n_186), .Y(n_177) );
INVxp67_ASAP7_75t_L g514 ( .A(n_178), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g515 ( .A(n_183), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_183), .A2(n_518), .B(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_184), .B(n_187), .Y(n_520) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_186), .B(n_515), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_192), .B(n_439), .Y(n_191) );
NOR5xp2_ASAP7_75t_L g192 ( .A(n_193), .B(n_370), .C(n_399), .D(n_419), .E(n_426), .Y(n_192) );
OAI211xp5_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_250), .B(n_314), .C(n_357), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_195), .A2(n_442), .B1(n_444), .B2(n_445), .Y(n_441) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_229), .Y(n_195) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_196), .Y(n_317) );
AND2x4_ASAP7_75t_L g350 ( .A(n_196), .B(n_351), .Y(n_350) );
INVx5_ASAP7_75t_L g368 ( .A(n_196), .Y(n_368) );
AND2x2_ASAP7_75t_L g377 ( .A(n_196), .B(n_369), .Y(n_377) );
AND2x2_ASAP7_75t_L g389 ( .A(n_196), .B(n_254), .Y(n_389) );
AND2x2_ASAP7_75t_L g485 ( .A(n_196), .B(n_353), .Y(n_485) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_226), .Y(n_196) );
AOI21xp5_ASAP7_75t_SL g197 ( .A1(n_198), .A2(n_206), .B(n_219), .Y(n_197) );
BUFx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_205), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_201), .B(n_205), .Y(n_294) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
INVx1_ASAP7_75t_L g217 ( .A(n_202), .Y(n_217) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g208 ( .A(n_203), .Y(n_208) );
INVx1_ASAP7_75t_L g301 ( .A(n_203), .Y(n_301) );
INVx1_ASAP7_75t_L g209 ( .A(n_204), .Y(n_209) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_204), .Y(n_213) );
INVx3_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_204), .Y(n_245) );
INVx1_ASAP7_75t_L g312 ( .A(n_204), .Y(n_312) );
BUFx3_ASAP7_75t_L g218 ( .A(n_205), .Y(n_218) );
INVx4_ASAP7_75t_SL g248 ( .A(n_205), .Y(n_248) );
INVx5_ASAP7_75t_L g237 ( .A(n_207), .Y(n_237) );
AND2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
BUFx3_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_208), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_216), .Y(n_210) );
INVx2_ASAP7_75t_L g215 ( .A(n_212), .Y(n_215) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx4_ASAP7_75t_L g274 ( .A(n_213), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_215), .A2(n_260), .B(n_261), .C(n_262), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_215), .A2(n_262), .B(n_286), .C(n_287), .Y(n_285) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_215), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_216), .B(n_248), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_216), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g228 ( .A(n_221), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_221), .A2(n_256), .B(n_257), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_221), .A2(n_283), .B(n_284), .Y(n_282) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_222), .B(n_223), .Y(n_221) );
AND2x2_ASAP7_75t_L g233 ( .A(n_222), .B(n_223), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g351 ( .A(n_229), .Y(n_351) );
AND2x2_ASAP7_75t_L g369 ( .A(n_229), .B(n_323), .Y(n_369) );
AND2x2_ASAP7_75t_L g388 ( .A(n_229), .B(n_322), .Y(n_388) );
AND2x2_ASAP7_75t_L g428 ( .A(n_229), .B(n_368), .Y(n_428) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_234), .B(n_249), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_231), .B(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_231), .A2(n_292), .B(n_302), .Y(n_291) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_231), .A2(n_324), .B(n_332), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_231), .B(n_333), .Y(n_332) );
INVx4_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_232), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_232), .A2(n_308), .B(n_309), .Y(n_307) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g304 ( .A(n_233), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_236), .A2(n_237), .B(n_238), .C(n_248), .Y(n_235) );
INVx2_ASAP7_75t_L g258 ( .A(n_237), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_237), .A2(n_248), .B(n_271), .C(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_240), .B(n_276), .Y(n_275) );
INVx5_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx4_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_247), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_248), .Y(n_263) );
INVxp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_278), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI322xp5_ASAP7_75t_L g487 ( .A1(n_253), .A2(n_289), .A3(n_342), .B1(n_350), .B2(n_404), .C1(n_488), .C2(n_491), .Y(n_487) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_266), .Y(n_253) );
INVx5_ASAP7_75t_L g319 ( .A(n_254), .Y(n_319) );
AND2x2_ASAP7_75t_L g336 ( .A(n_254), .B(n_321), .Y(n_336) );
BUFx2_ASAP7_75t_L g414 ( .A(n_254), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_254), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g491 ( .A(n_254), .B(n_398), .Y(n_491) );
OR2x6_ASAP7_75t_L g254 ( .A(n_255), .B(n_264), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_266), .B(n_280), .Y(n_345) );
INVx1_ASAP7_75t_L g372 ( .A(n_266), .Y(n_372) );
AND2x2_ASAP7_75t_L g385 ( .A(n_266), .B(n_305), .Y(n_385) );
AND2x2_ASAP7_75t_L g486 ( .A(n_266), .B(n_404), .Y(n_486) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g340 ( .A(n_267), .B(n_280), .Y(n_340) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_267), .Y(n_348) );
OR2x2_ASAP7_75t_L g355 ( .A(n_267), .B(n_305), .Y(n_355) );
AND2x2_ASAP7_75t_L g365 ( .A(n_267), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_267), .B(n_291), .Y(n_394) );
INVxp67_ASAP7_75t_L g418 ( .A(n_267), .Y(n_418) );
AND2x2_ASAP7_75t_L g425 ( .A(n_267), .B(n_289), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_267), .B(n_305), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_267), .B(n_290), .Y(n_451) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_277), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_273), .A2(n_327), .B(n_328), .C(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_289), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_280), .B(n_306), .Y(n_395) );
OR2x2_ASAP7_75t_L g417 ( .A(n_280), .B(n_290), .Y(n_417) );
AND2x2_ASAP7_75t_L g430 ( .A(n_280), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_280), .B(n_385), .Y(n_436) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_280), .A2(n_441), .B(n_446), .C(n_455), .Y(n_440) );
AND2x2_ASAP7_75t_L g501 ( .A(n_280), .B(n_305), .Y(n_501) );
INVx5_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g354 ( .A(n_281), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_281), .B(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_281), .B(n_349), .Y(n_361) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_281), .Y(n_363) );
OR2x2_ASAP7_75t_L g374 ( .A(n_281), .B(n_290), .Y(n_374) );
AND2x2_ASAP7_75t_SL g379 ( .A(n_281), .B(n_365), .Y(n_379) );
AND2x2_ASAP7_75t_L g404 ( .A(n_281), .B(n_290), .Y(n_404) );
AND2x2_ASAP7_75t_L g424 ( .A(n_281), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g462 ( .A(n_281), .B(n_289), .Y(n_462) );
OR2x2_ASAP7_75t_L g465 ( .A(n_281), .B(n_451), .Y(n_465) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_288), .Y(n_281) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_305), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_290), .A2(n_409), .B(n_412), .C(n_418), .Y(n_408) );
INVx5_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_291), .B(n_305), .Y(n_339) );
AND2x2_ASAP7_75t_L g343 ( .A(n_291), .B(n_306), .Y(n_343) );
OR2x2_ASAP7_75t_L g349 ( .A(n_291), .B(n_305), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_295), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_299), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_299), .A2(n_311), .B(n_313), .Y(n_310) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_SL g366 ( .A(n_305), .Y(n_366) );
OR2x2_ASAP7_75t_L g494 ( .A(n_305), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_334), .B(n_337), .C(n_346), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI31xp33_ASAP7_75t_L g419 ( .A1(n_316), .A2(n_420), .A3(n_422), .B(n_423), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_317), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_318), .B(n_350), .Y(n_356) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_319), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g376 ( .A(n_319), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g381 ( .A(n_319), .B(n_351), .Y(n_381) );
AND2x2_ASAP7_75t_L g391 ( .A(n_319), .B(n_350), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_319), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g411 ( .A(n_319), .B(n_368), .Y(n_411) );
AND2x2_ASAP7_75t_L g416 ( .A(n_319), .B(n_388), .Y(n_416) );
OR2x2_ASAP7_75t_L g435 ( .A(n_319), .B(n_321), .Y(n_435) );
OR2x2_ASAP7_75t_L g437 ( .A(n_319), .B(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_319), .Y(n_484) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g384 ( .A(n_321), .B(n_351), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_321), .B(n_368), .Y(n_407) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g353 ( .A(n_323), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_331), .Y(n_324) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g444 ( .A(n_336), .B(n_368), .Y(n_444) );
AOI322xp5_ASAP7_75t_L g446 ( .A1(n_336), .A2(n_350), .A3(n_388), .B1(n_447), .B2(n_448), .C1(n_449), .C2(n_452), .Y(n_446) );
INVx1_ASAP7_75t_L g454 ( .A(n_336), .Y(n_454) );
NAND2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
INVx1_ASAP7_75t_SL g448 ( .A(n_338), .Y(n_448) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g400 ( .A(n_339), .B(n_345), .Y(n_400) );
INVx1_ASAP7_75t_L g431 ( .A(n_339), .Y(n_431) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI32xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .A3(n_352), .B1(n_354), .B2(n_356), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AOI21xp33_ASAP7_75t_SL g386 ( .A1(n_349), .A2(n_364), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g401 ( .A(n_350), .Y(n_401) );
AND2x4_ASAP7_75t_L g398 ( .A(n_351), .B(n_368), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_351), .B(n_434), .Y(n_433) );
AOI322xp5_ASAP7_75t_L g463 ( .A1(n_352), .A2(n_379), .A3(n_398), .B1(n_431), .B2(n_464), .C1(n_466), .C2(n_467), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_352), .A2(n_429), .B1(n_493), .B2(n_494), .C(n_496), .Y(n_492) );
AND2x2_ASAP7_75t_L g380 ( .A(n_353), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g360 ( .A(n_355), .Y(n_360) );
OR2x2_ASAP7_75t_L g432 ( .A(n_355), .B(n_417), .Y(n_432) );
OAI31xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .A3(n_362), .B(n_367), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_358), .A2(n_391), .B1(n_392), .B2(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g403 ( .A(n_360), .B(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_362), .A2(n_403), .B1(n_456), .B2(n_459), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g445 ( .A(n_365), .B(n_414), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_365), .B(n_404), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_366), .B(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g479 ( .A(n_366), .B(n_417), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_367), .A2(n_462), .B1(n_475), .B2(n_478), .Y(n_474) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
AND2x2_ASAP7_75t_L g466 ( .A(n_368), .B(n_388), .Y(n_466) );
OR2x2_ASAP7_75t_L g468 ( .A(n_368), .B(n_435), .Y(n_468) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_368), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_369), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_369), .B(n_414), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B(n_378), .C(n_390), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_382), .B2(n_385), .C(n_386), .Y(n_378) );
INVxp67_ASAP7_75t_L g490 ( .A(n_381), .Y(n_490) );
INVx1_ASAP7_75t_L g457 ( .A(n_382), .Y(n_457) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g421 ( .A(n_383), .B(n_388), .Y(n_421) );
INVx1_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_384), .B(n_411), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g453 ( .A(n_388), .Y(n_453) );
AND2x2_ASAP7_75t_L g459 ( .A(n_388), .B(n_414), .Y(n_459) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_SL g447 ( .A(n_395), .Y(n_447) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_398), .B(n_434), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_402), .B2(n_405), .C(n_408), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g495 ( .A(n_404), .Y(n_495) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g413 ( .A(n_407), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_411), .B(n_470), .Y(n_469) );
AOI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B(n_417), .Y(n_412) );
OAI211xp5_ASAP7_75t_SL g460 ( .A1(n_415), .A2(n_461), .B(n_463), .C(n_469), .Y(n_460) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g472 ( .A(n_417), .Y(n_472) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI222xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_432), .B2(n_433), .C1(n_436), .C2(n_437), .Y(n_426) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g502 ( .A(n_433), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_434), .B(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_434), .A2(n_481), .B1(n_483), .B2(n_486), .Y(n_480) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
NOR4xp25_ASAP7_75t_L g439 ( .A(n_440), .B(n_460), .C(n_473), .D(n_492), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_442), .B(n_472), .Y(n_482) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g449 ( .A(n_447), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_450), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_480), .C(n_487), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g489 ( .A(n_485), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_499), .B(n_502), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g519 ( .A(n_506), .Y(n_519) );
OAI322xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .A3(n_511), .B1(n_515), .B2(n_516), .C1(n_521), .C2(n_523), .Y(n_508) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
endmodule