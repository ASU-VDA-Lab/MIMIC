module fake_aes_3061_n_990 (n_117, n_219, n_44, n_133, n_149, n_81, n_69, n_214, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_990);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_990;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_844;
wire n_818;
wire n_230;
wire n_274;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_490;
wire n_247;
wire n_393;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_224;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_150), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_181), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_82), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_203), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_161), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_4), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_215), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_128), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_15), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_153), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_135), .Y(n_234) );
INVxp33_ASAP7_75t_SL g235 ( .A(n_70), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_218), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_149), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_213), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_141), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_205), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_219), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_147), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_120), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_112), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_40), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_187), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_42), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_162), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_35), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_36), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_49), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_85), .Y(n_252) );
NOR2xp67_ASAP7_75t_L g253 ( .A(n_197), .B(n_216), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_25), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_22), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_29), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_100), .B(n_66), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_173), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_127), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_62), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_186), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_118), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_121), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_140), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_182), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_52), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_172), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_204), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_139), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_137), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_94), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_69), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_0), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_68), .Y(n_274) );
NOR2xp67_ASAP7_75t_L g275 ( .A(n_180), .B(n_102), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_77), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_154), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_176), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_89), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_70), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_169), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_114), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_129), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_111), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_191), .Y(n_287) );
INVxp33_ASAP7_75t_L g288 ( .A(n_51), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_69), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_47), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_62), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_152), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_138), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_41), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_202), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_189), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_208), .Y(n_297) );
CKINVDCx14_ASAP7_75t_R g298 ( .A(n_131), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_123), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_211), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_77), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_90), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_86), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_17), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_179), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_217), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_84), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_97), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_6), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_142), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_83), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_108), .Y(n_312) );
BUFx2_ASAP7_75t_SL g313 ( .A(n_157), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_6), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_198), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_117), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_87), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_93), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_79), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_29), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_53), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_50), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_201), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_130), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_165), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_78), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_53), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_88), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_54), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_113), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_185), .Y(n_331) );
CKINVDCx16_ASAP7_75t_R g332 ( .A(n_34), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_107), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_170), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_24), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_109), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_75), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_171), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_124), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_68), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_15), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_214), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_200), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_274), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_324), .B(n_0), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_220), .B(n_248), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_322), .B(n_1), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_274), .B(n_1), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_228), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_269), .Y(n_351) );
NAND2xp33_ASAP7_75t_L g352 ( .A(n_279), .B(n_101), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_304), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_230), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_264), .B(n_2), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_228), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_245), .A2(n_5), .B1(n_2), .B2(n_3), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_258), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_251), .B(n_3), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_269), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_288), .B(n_5), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_258), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_264), .B(n_7), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_262), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_262), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_305), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_251), .B(n_7), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_305), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_310), .B(n_8), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_221), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_326), .B(n_8), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_222), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_315), .A2(n_104), .B(n_103), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_224), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_315), .Y(n_375) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_226), .A2(n_9), .B(n_10), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_323), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_323), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_333), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_227), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_354), .A2(n_332), .B1(n_235), .B2(n_306), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_344), .B(n_298), .Y(n_383) );
AND2x6_ASAP7_75t_L g384 ( .A(n_347), .B(n_233), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_351), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_346), .B(n_330), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_346), .B(n_231), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_347), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_344), .B(n_229), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_347), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_344), .B(n_229), .Y(n_395) );
NAND2xp33_ASAP7_75t_L g396 ( .A(n_370), .B(n_261), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_361), .A2(n_225), .B1(n_250), .B2(n_247), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_356), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
AND2x6_ASAP7_75t_L g402 ( .A(n_355), .B(n_234), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
AND2x6_ASAP7_75t_L g404 ( .A(n_355), .B(n_236), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_358), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_370), .B(n_232), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_361), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
INVx4_ASAP7_75t_L g410 ( .A(n_363), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_357), .B(n_329), .C(n_289), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g412 ( .A(n_371), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_363), .Y(n_413) );
OR2x6_ASAP7_75t_L g414 ( .A(n_357), .B(n_313), .Y(n_414) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_352), .B(n_237), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_363), .A2(n_256), .B1(n_271), .B2(n_254), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_351), .Y(n_417) );
XNOR2xp5_ASAP7_75t_L g418 ( .A(n_371), .B(n_249), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_372), .B(n_255), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_371), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_351), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_358), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_351), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_358), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_383), .B(n_345), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_410), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_407), .A2(n_352), .B1(n_345), .B2(n_369), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_410), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_388), .A2(n_393), .B(n_391), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_383), .B(n_372), .Y(n_433) );
BUFx6f_ASAP7_75t_SL g434 ( .A(n_414), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_392), .B(n_374), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_392), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_415), .A2(n_369), .B1(n_235), .B2(n_306), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_406), .B(n_374), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_390), .B(n_380), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_415), .A2(n_223), .B1(n_266), .B2(n_260), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_416), .B(n_240), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_419), .B(n_359), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_414), .B(n_367), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_397), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_395), .B(n_367), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_399), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_421), .B(n_266), .Y(n_448) );
NOR2xp33_ASAP7_75t_SL g449 ( .A(n_412), .B(n_249), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_421), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_389), .B(n_377), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_398), .A2(n_302), .B1(n_303), .B2(n_278), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_412), .B(n_278), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_388), .A2(n_303), .B1(n_307), .B2(n_302), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_418), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_381), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_384), .A2(n_308), .B1(n_320), .B2(n_314), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_399), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_408), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_387), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_400), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_384), .B(n_377), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_384), .B(n_402), .Y(n_464) );
CKINVDCx11_ASAP7_75t_R g465 ( .A(n_414), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_384), .B(n_348), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_393), .B(n_387), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_403), .Y(n_468) );
AND2x6_ASAP7_75t_SL g469 ( .A(n_414), .B(n_272), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_394), .B(n_238), .Y(n_470) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_414), .A2(n_311), .B1(n_341), .B2(n_337), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_394), .B(n_239), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_394), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_413), .A2(n_311), .B1(n_341), .B2(n_337), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_402), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_402), .B(n_243), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_408), .B(n_241), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_408), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_396), .B(n_353), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_402), .A2(n_376), .B1(n_375), .B2(n_368), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_402), .Y(n_481) );
INVx5_ASAP7_75t_L g482 ( .A(n_404), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_404), .A2(n_376), .B1(n_375), .B2(n_368), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_404), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_404), .A2(n_340), .B1(n_409), .B2(n_405), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_425), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_425), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_420), .B(n_242), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_404), .B(n_244), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_405), .B(n_340), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_404), .B(n_246), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_409), .B(n_246), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_423), .Y(n_493) );
INVx5_ASAP7_75t_L g494 ( .A(n_420), .Y(n_494) );
AND2x6_ASAP7_75t_SL g495 ( .A(n_423), .B(n_273), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_385), .B(n_259), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_385), .B(n_263), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_385), .A2(n_376), .B1(n_375), .B2(n_368), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_386), .A2(n_349), .B1(n_376), .B2(n_319), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_386), .B(n_263), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_386), .A2(n_376), .B1(n_375), .B2(n_368), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_488), .A2(n_373), .B(n_401), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_482), .B(n_265), .Y(n_503) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_429), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_493), .Y(n_505) );
BUFx12f_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_439), .A2(n_373), .B(n_362), .C(n_364), .Y(n_507) );
OAI22xp5_ASAP7_75t_SL g508 ( .A1(n_471), .A2(n_252), .B1(n_283), .B2(n_265), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_444), .A2(n_362), .B1(n_364), .B2(n_350), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_439), .A2(n_365), .B(n_366), .C(n_350), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_429), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_426), .B(n_446), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_490), .B(n_284), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_444), .A2(n_366), .B1(n_365), .B2(n_376), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_493), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_443), .B(n_286), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_468), .B(n_281), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_482), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_450), .B(n_282), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_469), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_482), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_450), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_433), .B(n_286), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_428), .A2(n_291), .B(n_294), .C(n_290), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_430), .B(n_448), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_482), .B(n_292), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_453), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_458), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_461), .Y(n_529) );
BUFx4f_ASAP7_75t_SL g530 ( .A(n_442), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_438), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_475), .B(n_301), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_467), .A2(n_422), .B(n_417), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_461), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_437), .B(n_309), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_467), .A2(n_422), .B(n_417), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_427), .Y(n_537) );
O2A1O1Ixp5_ASAP7_75t_L g538 ( .A1(n_451), .A2(n_422), .B(n_424), .C(n_257), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_434), .A2(n_318), .B1(n_321), .B2(n_317), .Y(n_539) );
INVx5_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_498), .A2(n_424), .B(n_366), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_431), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_452), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_480), .A2(n_365), .B1(n_328), .B2(n_335), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_481), .B(n_478), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_449), .B(n_327), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_441), .A2(n_343), .B1(n_342), .B2(n_267), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_454), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_432), .A2(n_270), .B(n_268), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_457), .B(n_312), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_456), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_470), .A2(n_277), .B(n_276), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_458), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_480), .A2(n_483), .B1(n_485), .B2(n_499), .Y(n_555) );
AOI21xp5_ASAP7_75t_SL g556 ( .A1(n_464), .A2(n_285), .B(n_280), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_473), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_487), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_472), .A2(n_293), .B(n_287), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_483), .A2(n_296), .B1(n_297), .B2(n_295), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_476), .B(n_299), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_460), .B(n_300), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_440), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_445), .B(n_9), .Y(n_564) );
INVx4_ASAP7_75t_L g565 ( .A(n_494), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_479), .B(n_316), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_479), .A2(n_477), .B1(n_459), .B2(n_462), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_447), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_492), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_489), .B(n_325), .Y(n_570) );
BUFx2_ASAP7_75t_L g571 ( .A(n_491), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_466), .A2(n_334), .B1(n_336), .B2(n_331), .Y(n_572) );
AOI21xp33_ASAP7_75t_L g573 ( .A1(n_463), .A2(n_339), .B(n_338), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_496), .B(n_10), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_498), .A2(n_501), .B1(n_500), .B2(n_497), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_494), .A2(n_378), .B(n_360), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_458), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_435), .B(n_253), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_486), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_486), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_486), .Y(n_581) );
NAND2x1p5_ASAP7_75t_L g582 ( .A(n_482), .B(n_275), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_488), .A2(n_378), .B(n_360), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_450), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_439), .A2(n_378), .B(n_13), .C(n_11), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_482), .B(n_378), .Y(n_586) );
NOR2xp33_ASAP7_75t_SL g587 ( .A(n_429), .B(n_105), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_488), .A2(n_110), .B(n_106), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_429), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_455), .B(n_12), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_435), .B(n_14), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_450), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_482), .B(n_14), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_436), .B(n_16), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_435), .B(n_16), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_444), .A2(n_19), .B1(n_17), .B2(n_18), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_493), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_493), .Y(n_598) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_449), .B(n_18), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_488), .A2(n_116), .B(n_115), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_488), .A2(n_122), .B(n_119), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_435), .B(n_19), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_493), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_436), .B(n_20), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_486), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_436), .B(n_20), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_444), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_592), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_584), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_512), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_522), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_543), .A2(n_23), .B(n_24), .C(n_25), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_531), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_525), .B(n_26), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_505), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_527), .B(n_27), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_549), .B(n_28), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_515), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_535), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_524), .A2(n_33), .B(n_34), .C(n_35), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_605), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_552), .B(n_33), .Y(n_622) );
INVx4_ASAP7_75t_L g623 ( .A(n_506), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_502), .A2(n_126), .B(n_125), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_563), .Y(n_625) );
BUFx12f_ASAP7_75t_L g626 ( .A(n_545), .Y(n_626) );
CKINVDCx8_ASAP7_75t_R g627 ( .A(n_520), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_569), .B(n_37), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_SL g629 ( .A1(n_507), .A2(n_510), .B(n_585), .C(n_514), .Y(n_629) );
INVx3_ASAP7_75t_SL g630 ( .A(n_599), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_597), .B(n_38), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_598), .A2(n_39), .B1(n_42), .B2(n_43), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_564), .Y(n_633) );
AO31x2_ASAP7_75t_L g634 ( .A1(n_555), .A2(n_44), .A3(n_45), .B(n_46), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_603), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_530), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_528), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_568), .Y(n_638) );
INVxp67_ASAP7_75t_L g639 ( .A(n_606), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_538), .A2(n_133), .B(n_132), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_596), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_519), .B(n_55), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_558), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_528), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_516), .B(n_55), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_548), .B(n_56), .Y(n_646) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_541), .A2(n_136), .B(n_134), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_540), .B(n_56), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_607), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_575), .A2(n_536), .B(n_533), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_591), .Y(n_651) );
NOR4xp25_ASAP7_75t_L g652 ( .A(n_544), .B(n_60), .C(n_61), .D(n_63), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_590), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_SL g654 ( .A1(n_514), .A2(n_167), .B(n_212), .C(n_210), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_547), .B(n_517), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_595), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_523), .B(n_63), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_528), .A2(n_166), .B(n_209), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_593), .A2(n_164), .B(n_207), .C(n_206), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_540), .B(n_64), .Y(n_660) );
BUFx10_ASAP7_75t_L g661 ( .A(n_594), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_513), .B(n_65), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_565), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_602), .A2(n_66), .B(n_67), .C(n_71), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_578), .B(n_72), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_540), .B(n_73), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_604), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_561), .A2(n_74), .B(n_75), .C(n_76), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g669 ( .A1(n_570), .A2(n_80), .B(n_81), .C(n_83), .Y(n_669) );
INVx5_ASAP7_75t_L g670 ( .A(n_521), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_539), .B(n_88), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_574), .B(n_91), .C(n_92), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_560), .A2(n_93), .B(n_94), .C(n_95), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_566), .B(n_95), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_504), .Y(n_675) );
AND2x6_ASAP7_75t_SL g676 ( .A(n_551), .B(n_96), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_567), .B(n_96), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_587), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_546), .Y(n_679) );
INVx4_ASAP7_75t_SL g680 ( .A(n_504), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_550), .A2(n_143), .B(n_144), .C(n_145), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_554), .A2(n_146), .B(n_148), .Y(n_682) );
AOI221x1_ASAP7_75t_L g683 ( .A1(n_509), .A2(n_576), .B1(n_573), .B2(n_583), .C(n_556), .Y(n_683) );
BUFx12f_ASAP7_75t_L g684 ( .A(n_582), .Y(n_684) );
AOI221x1_ASAP7_75t_L g685 ( .A1(n_588), .A2(n_156), .B1(n_158), .B2(n_159), .C(n_160), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_537), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_577), .A2(n_163), .B(n_168), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_546), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_518), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_579), .Y(n_690) );
AO32x2_ASAP7_75t_L g691 ( .A1(n_518), .A2(n_174), .A3(n_175), .B1(n_177), .B2(n_178), .Y(n_691) );
BUFx4_ASAP7_75t_R g692 ( .A(n_580), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_562), .Y(n_693) );
INVx3_ASAP7_75t_L g694 ( .A(n_521), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_581), .Y(n_695) );
INVx4_ASAP7_75t_L g696 ( .A(n_521), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_542), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_571), .A2(n_190), .B1(n_192), .B2(n_193), .Y(n_698) );
BUFx3_ASAP7_75t_L g699 ( .A(n_511), .Y(n_699) );
AO31x2_ASAP7_75t_L g700 ( .A1(n_600), .A2(n_194), .A3(n_195), .B(n_196), .Y(n_700) );
CKINVDCx11_ASAP7_75t_R g701 ( .A(n_511), .Y(n_701) );
CKINVDCx6p67_ASAP7_75t_R g702 ( .A(n_532), .Y(n_702) );
OAI21x1_ASAP7_75t_L g703 ( .A1(n_601), .A2(n_586), .B(n_553), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_557), .Y(n_704) );
AO31x2_ASAP7_75t_L g705 ( .A1(n_559), .A2(n_529), .A3(n_534), .B(n_572), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_503), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_589), .B(n_526), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_543), .A2(n_524), .B(n_525), .C(n_585), .Y(n_708) );
CKINVDCx8_ASAP7_75t_R g709 ( .A(n_545), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_549), .B(n_412), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_527), .A2(n_471), .B1(n_434), .B2(n_414), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_543), .A2(n_524), .B(n_525), .C(n_585), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_527), .A2(n_471), .B1(n_434), .B2(n_414), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_592), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_641), .A2(n_649), .B1(n_610), .B2(n_648), .Y(n_715) );
AO31x2_ASAP7_75t_L g716 ( .A1(n_683), .A2(n_685), .A3(n_624), .B(n_681), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_611), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_638), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_630), .A2(n_710), .B1(n_655), .B2(n_711), .Y(n_719) );
BUFx2_ASAP7_75t_L g720 ( .A(n_609), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_649), .A2(n_648), .B1(n_619), .B2(n_702), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_651), .B(n_656), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_665), .A2(n_633), .B1(n_713), .B2(n_652), .C(n_622), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_642), .B(n_616), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_608), .B(n_714), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_625), .Y(n_726) );
INVx3_ASAP7_75t_L g727 ( .A(n_670), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_613), .B(n_671), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_667), .A2(n_639), .B1(n_653), .B2(n_628), .C(n_646), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_645), .A2(n_654), .B(n_703), .Y(n_730) );
INVx2_ASAP7_75t_SL g731 ( .A(n_684), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_619), .A2(n_666), .B1(n_660), .B2(n_617), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_679), .B(n_662), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_674), .A2(n_657), .B(n_614), .Y(n_734) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_612), .A2(n_673), .B(n_677), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_660), .A2(n_666), .B1(n_678), .B2(n_672), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g737 ( .A1(n_672), .A2(n_664), .B(n_620), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_686), .Y(n_738) );
NOR2x1_ASAP7_75t_SL g739 ( .A(n_670), .B(n_663), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_631), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_688), .B(n_680), .Y(n_741) );
OAI21x1_ASAP7_75t_L g742 ( .A1(n_658), .A2(n_687), .B(n_682), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_692), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_621), .Y(n_744) );
OR2x6_ASAP7_75t_L g745 ( .A(n_688), .B(n_696), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_652), .A2(n_669), .B(n_668), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_704), .B(n_697), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_637), .A2(n_644), .B(n_659), .Y(n_748) );
AOI322xp5_ASAP7_75t_L g749 ( .A1(n_632), .A2(n_636), .A3(n_676), .B1(n_698), .B2(n_709), .C1(n_706), .C2(n_643), .Y(n_749) );
INVx3_ASAP7_75t_L g750 ( .A(n_696), .Y(n_750) );
BUFx2_ASAP7_75t_L g751 ( .A(n_699), .Y(n_751) );
AO31x2_ASAP7_75t_L g752 ( .A1(n_615), .A2(n_618), .A3(n_635), .B(n_634), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_690), .B(n_695), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_690), .A2(n_695), .B1(n_689), .B2(n_644), .Y(n_754) );
AO21x2_ASAP7_75t_L g755 ( .A1(n_707), .A2(n_634), .B(n_691), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_705), .B(n_689), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_705), .B(n_694), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_661), .B(n_680), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_701), .B(n_627), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_700), .Y(n_760) );
OAI21x1_ASAP7_75t_L g761 ( .A1(n_691), .A2(n_650), .B(n_647), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_641), .A2(n_649), .B1(n_610), .B2(n_648), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_610), .B(n_455), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_641), .A2(n_649), .B1(n_610), .B2(n_648), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_610), .B(n_455), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_625), .Y(n_766) );
INVx3_ASAP7_75t_L g767 ( .A(n_670), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_641), .A2(n_649), .B1(n_610), .B2(n_648), .Y(n_768) );
OA21x2_ASAP7_75t_L g769 ( .A1(n_640), .A2(n_507), .B(n_650), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_641), .A2(n_471), .B1(n_630), .B2(n_599), .Y(n_770) );
CKINVDCx11_ASAP7_75t_R g771 ( .A(n_623), .Y(n_771) );
INVx4_ASAP7_75t_L g772 ( .A(n_692), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_625), .Y(n_773) );
OA21x2_ASAP7_75t_L g774 ( .A1(n_640), .A2(n_507), .B(n_650), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_610), .B(n_531), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_675), .Y(n_776) );
NAND2x1p5_ASAP7_75t_L g777 ( .A(n_670), .B(n_663), .Y(n_777) );
INVx3_ASAP7_75t_L g778 ( .A(n_670), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_610), .B(n_512), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_610), .B(n_531), .Y(n_780) );
AO21x2_ASAP7_75t_L g781 ( .A1(n_640), .A2(n_629), .B(n_507), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_610), .B(n_693), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_625), .Y(n_783) );
CKINVDCx11_ASAP7_75t_R g784 ( .A(n_623), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_708), .A2(n_555), .B(n_712), .Y(n_785) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_610), .A2(n_411), .B1(n_535), .B2(n_524), .C(n_710), .Y(n_786) );
BUFx2_ASAP7_75t_L g787 ( .A(n_610), .Y(n_787) );
AO21x2_ASAP7_75t_L g788 ( .A1(n_640), .A2(n_629), .B(n_507), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_610), .B(n_693), .Y(n_789) );
BUFx2_ASAP7_75t_L g790 ( .A(n_610), .Y(n_790) );
BUFx8_ASAP7_75t_L g791 ( .A(n_626), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_610), .B(n_455), .Y(n_792) );
AOI222xp33_ASAP7_75t_L g793 ( .A1(n_610), .A2(n_471), .B1(n_474), .B2(n_508), .C1(n_357), .C2(n_599), .Y(n_793) );
AO31x2_ASAP7_75t_L g794 ( .A1(n_650), .A2(n_507), .A3(n_683), .B(n_514), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_610), .B(n_455), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_610), .B(n_512), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_610), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_641), .A2(n_649), .B1(n_610), .B2(n_648), .Y(n_798) );
OR2x6_ASAP7_75t_L g799 ( .A(n_684), .B(n_506), .Y(n_799) );
BUFx3_ASAP7_75t_L g800 ( .A(n_777), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_766), .B(n_773), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_783), .B(n_738), .Y(n_802) );
AOI21xp5_ASAP7_75t_SL g803 ( .A1(n_715), .A2(n_764), .B(n_762), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_756), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_757), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_726), .B(n_747), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_794), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_794), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_794), .Y(n_809) );
OA21x2_ASAP7_75t_L g810 ( .A1(n_785), .A2(n_760), .B(n_730), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_718), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_747), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_793), .A2(n_721), .B1(n_770), .B2(n_764), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_728), .B(n_717), .Y(n_814) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_787), .Y(n_815) );
AND2x4_ASAP7_75t_L g816 ( .A(n_750), .B(n_745), .Y(n_816) );
INVx5_ASAP7_75t_L g817 ( .A(n_772), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_793), .A2(n_721), .B1(n_715), .B2(n_762), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_790), .Y(n_819) );
INVx3_ASAP7_75t_L g820 ( .A(n_727), .Y(n_820) );
BUFx3_ASAP7_75t_L g821 ( .A(n_777), .Y(n_821) );
OR2x6_ASAP7_75t_L g822 ( .A(n_768), .B(n_798), .Y(n_822) );
INVx4_ASAP7_75t_L g823 ( .A(n_745), .Y(n_823) );
AO21x2_ASAP7_75t_L g824 ( .A1(n_746), .A2(n_781), .B(n_788), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_753), .Y(n_825) );
BUFx3_ASAP7_75t_L g826 ( .A(n_727), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_779), .B(n_796), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_763), .B(n_765), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_782), .B(n_789), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_753), .Y(n_830) );
OA21x2_ASAP7_75t_L g831 ( .A1(n_734), .A2(n_737), .B(n_735), .Y(n_831) );
OR2x2_ASAP7_75t_L g832 ( .A(n_782), .B(n_789), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_768), .A2(n_786), .B1(n_732), .B2(n_723), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_755), .Y(n_834) );
OR2x6_ASAP7_75t_L g835 ( .A(n_732), .B(n_736), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_755), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_769), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_774), .Y(n_838) );
INVx4_ASAP7_75t_L g839 ( .A(n_767), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g840 ( .A(n_749), .B(n_729), .C(n_719), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_722), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_775), .B(n_780), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_741), .B(n_767), .Y(n_843) );
BUFx2_ASAP7_75t_L g844 ( .A(n_754), .Y(n_844) );
NOR2x1_ASAP7_75t_R g845 ( .A(n_771), .B(n_784), .Y(n_845) );
AO21x2_ASAP7_75t_L g846 ( .A1(n_748), .A2(n_754), .B(n_742), .Y(n_846) );
BUFx2_ASAP7_75t_L g847 ( .A(n_720), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_740), .B(n_724), .Y(n_848) );
OAI31xp33_ASAP7_75t_L g849 ( .A1(n_780), .A2(n_792), .A3(n_795), .B(n_743), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_752), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_725), .B(n_778), .Y(n_851) );
OR2x2_ASAP7_75t_L g852 ( .A(n_752), .B(n_744), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_778), .B(n_752), .Y(n_853) );
AND2x4_ASAP7_75t_L g854 ( .A(n_741), .B(n_739), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_797), .B(n_733), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_751), .B(n_776), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_716), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g858 ( .A1(n_758), .A2(n_731), .B(n_759), .Y(n_858) );
OA21x2_ASAP7_75t_L g859 ( .A1(n_799), .A2(n_791), .B(n_761), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_799), .Y(n_860) );
OR2x6_ASAP7_75t_L g861 ( .A(n_803), .B(n_822), .Y(n_861) );
INVx4_ASAP7_75t_L g862 ( .A(n_823), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_835), .B(n_853), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_835), .B(n_853), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_835), .B(n_822), .Y(n_865) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_815), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_804), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_835), .B(n_822), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_819), .Y(n_869) );
AND2x4_ASAP7_75t_L g870 ( .A(n_822), .B(n_805), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_850), .B(n_814), .Y(n_871) );
BUFx2_ASAP7_75t_L g872 ( .A(n_844), .Y(n_872) );
OR2x2_ASAP7_75t_L g873 ( .A(n_832), .B(n_852), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_806), .B(n_829), .Y(n_874) );
NAND2x1_ASAP7_75t_L g875 ( .A(n_803), .B(n_823), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_827), .B(n_828), .Y(n_876) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_840), .A2(n_813), .B1(n_818), .B2(n_833), .C(n_829), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_847), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_806), .B(n_825), .Y(n_879) );
NAND3xp33_ASAP7_75t_L g880 ( .A(n_833), .B(n_849), .C(n_831), .Y(n_880) );
BUFx2_ASAP7_75t_L g881 ( .A(n_859), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_825), .B(n_830), .Y(n_882) );
HB1xp67_ASAP7_75t_L g883 ( .A(n_851), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_811), .B(n_848), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_852), .Y(n_885) );
CKINVDCx6p67_ASAP7_75t_R g886 ( .A(n_817), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_811), .B(n_801), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_801), .B(n_802), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_834), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_802), .B(n_841), .Y(n_890) );
INVx2_ASAP7_75t_SL g891 ( .A(n_854), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_812), .B(n_831), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_873), .B(n_807), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_882), .B(n_831), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_871), .B(n_808), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_889), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_892), .B(n_809), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_863), .B(n_857), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_886), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_876), .B(n_860), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_863), .B(n_857), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_864), .B(n_836), .Y(n_902) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_877), .A2(n_858), .B1(n_860), .B2(n_842), .C(n_855), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_874), .B(n_824), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_874), .B(n_810), .Y(n_905) );
AND2x4_ASAP7_75t_L g906 ( .A(n_861), .B(n_846), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_888), .B(n_810), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_888), .B(n_810), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_884), .B(n_810), .Y(n_909) );
NOR2x1_ASAP7_75t_L g910 ( .A(n_862), .B(n_839), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_884), .B(n_837), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_870), .B(n_838), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_878), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_867), .Y(n_914) );
INVxp67_ASAP7_75t_L g915 ( .A(n_900), .Y(n_915) );
INVx2_ASAP7_75t_SL g916 ( .A(n_910), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_914), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_904), .B(n_887), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_896), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_904), .B(n_887), .Y(n_920) );
NAND2x1_ASAP7_75t_L g921 ( .A(n_899), .B(n_881), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_914), .Y(n_922) );
OR2x2_ASAP7_75t_L g923 ( .A(n_894), .B(n_872), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_905), .B(n_865), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_905), .B(n_865), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_907), .B(n_868), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_913), .B(n_879), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_907), .B(n_868), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_908), .B(n_885), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_909), .B(n_890), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_908), .B(n_885), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_909), .B(n_890), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_911), .B(n_866), .Y(n_933) );
INVx1_ASAP7_75t_SL g934 ( .A(n_911), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_895), .B(n_869), .Y(n_935) );
NOR3xp33_ASAP7_75t_L g936 ( .A(n_903), .B(n_880), .C(n_845), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_919), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_929), .B(n_902), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_936), .A2(n_891), .B1(n_875), .B2(n_883), .Y(n_939) );
INVx4_ASAP7_75t_L g940 ( .A(n_916), .Y(n_940) );
AND2x4_ASAP7_75t_L g941 ( .A(n_916), .B(n_906), .Y(n_941) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_934), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_924), .B(n_902), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_924), .B(n_898), .Y(n_944) );
INVx2_ASAP7_75t_SL g945 ( .A(n_921), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_929), .B(n_898), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_931), .B(n_901), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_931), .B(n_901), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_917), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_927), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_933), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_918), .B(n_897), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_935), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_923), .B(n_893), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_922), .Y(n_955) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_915), .B(n_845), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_920), .B(n_897), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_925), .B(n_912), .Y(n_958) );
AOI21xp33_ASAP7_75t_SL g959 ( .A1(n_945), .A2(n_939), .B(n_956), .Y(n_959) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_942), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_940), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_944), .B(n_925), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_950), .B(n_926), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_937), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_954), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_951), .B(n_926), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_953), .B(n_928), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_960), .Y(n_968) );
AOI221xp5_ASAP7_75t_L g969 ( .A1(n_959), .A2(n_955), .B1(n_947), .B2(n_946), .C(n_948), .Y(n_969) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_961), .A2(n_938), .B1(n_930), .B2(n_932), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g971 ( .A1(n_965), .A2(n_941), .B1(n_943), .B2(n_949), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_962), .B(n_958), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_965), .A2(n_958), .B1(n_957), .B2(n_952), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_968), .B(n_962), .Y(n_974) );
O2A1O1Ixp33_ASAP7_75t_SL g975 ( .A1(n_969), .A2(n_967), .B(n_966), .C(n_963), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_970), .B(n_973), .Y(n_976) );
NAND2x1p5_ASAP7_75t_L g977 ( .A(n_972), .B(n_817), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_976), .B(n_971), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_974), .B(n_964), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_975), .B(n_964), .Y(n_980) );
AND2x4_ASAP7_75t_L g981 ( .A(n_978), .B(n_856), .Y(n_981) );
NAND3x1_ASAP7_75t_L g982 ( .A(n_980), .B(n_977), .C(n_820), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_981), .B(n_979), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_982), .Y(n_984) );
INVx2_ASAP7_75t_SL g985 ( .A(n_984), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_985), .B(n_983), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_986), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g988 ( .A(n_987), .B(n_800), .C(n_821), .Y(n_988) );
OAI22x1_ASAP7_75t_L g989 ( .A1(n_988), .A2(n_843), .B1(n_839), .B2(n_816), .Y(n_989) );
AOI21xp33_ASAP7_75t_L g990 ( .A1(n_989), .A2(n_826), .B(n_820), .Y(n_990) );
endmodule