module fake_jpeg_13665_n_571 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_571);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_571;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_18),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_63),
.Y(n_118)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_56),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_58),
.B(n_84),
.Y(n_155)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_59),
.Y(n_144)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx2_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_69),
.Y(n_135)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_23),
.B(n_18),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_36),
.A2(n_41),
.B1(n_28),
.B2(n_46),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_41),
.B1(n_49),
.B2(n_39),
.Y(n_122)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_25),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

CKINVDCx9p33_ASAP7_75t_R g158 ( 
.A(n_101),
.Y(n_158)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_47),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_109),
.B(n_130),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_25),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_111),
.B(n_117),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_120),
.B(n_127),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_122),
.A2(n_157),
.B1(n_29),
.B2(n_47),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_49),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_51),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_51),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_72),
.B(n_40),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_57),
.B(n_40),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_26),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_87),
.B(n_42),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_47),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_73),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_159),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_78),
.A2(n_28),
.B1(n_46),
.B2(n_33),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_42),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_160),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_54),
.A2(n_33),
.B1(n_46),
.B2(n_28),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_61),
.B1(n_95),
.B2(n_81),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_172),
.B(n_183),
.Y(n_264)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_182),
.A2(n_187),
.B1(n_213),
.B2(n_223),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_105),
.B1(n_103),
.B2(n_76),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_184),
.B(n_211),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_121),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_185),
.B(n_203),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_186),
.B(n_221),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_122),
.A2(n_101),
.B1(n_93),
.B2(n_82),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_202),
.B1(n_219),
.B2(n_160),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_197),
.Y(n_284)
);

CKINVDCx12_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_198),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_45),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_201),
.B(n_208),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_122),
.A2(n_77),
.B1(n_62),
.B2(n_71),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

CKINVDCx12_ASAP7_75t_R g205 ( 
.A(n_162),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_206),
.Y(n_282)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_108),
.B(n_44),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_138),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_209),
.B(n_212),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_27),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_210),
.B(n_181),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_118),
.A2(n_83),
.B1(n_79),
.B2(n_33),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_164),
.A2(n_29),
.B1(n_47),
.B2(n_69),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_220),
.B1(n_139),
.B2(n_170),
.Y(n_237)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_233),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_166),
.A2(n_29),
.B1(n_69),
.B2(n_47),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_1),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_229),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_142),
.A2(n_88),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_142),
.A2(n_144),
.B1(n_135),
.B2(n_125),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_224),
.A2(n_227),
.B1(n_228),
.B2(n_234),
.Y(n_254)
);

AO22x1_ASAP7_75t_SL g225 ( 
.A1(n_167),
.A2(n_88),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_226),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_118),
.B(n_2),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_144),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_171),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_113),
.B(n_4),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_5),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_161),
.Y(n_233)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_237),
.A2(n_239),
.B1(n_266),
.B2(n_273),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_139),
.B1(n_170),
.B2(n_165),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_238),
.A2(n_247),
.B1(n_285),
.B2(n_215),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_263),
.Y(n_292)
);

OAI22x1_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_112),
.B1(n_125),
.B2(n_165),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_189),
.A2(n_129),
.B(n_156),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_250),
.A2(n_185),
.B(n_195),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_262),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_186),
.Y(n_263)
);

OR2x4_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_119),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_222),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_220),
.A2(n_143),
.B1(n_147),
.B2(n_129),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_200),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_287),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_177),
.B(n_123),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_206),
.C(n_173),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_177),
.B(n_123),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_271),
.B(n_281),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_189),
.A2(n_147),
.B1(n_136),
.B2(n_124),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_183),
.A2(n_221),
.B1(n_232),
.B2(n_233),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_286),
.B1(n_199),
.B2(n_227),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_124),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_191),
.B(n_169),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_176),
.A2(n_169),
.B1(n_135),
.B2(n_112),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_203),
.A2(n_126),
.B1(n_156),
.B2(n_8),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_231),
.B(n_140),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_179),
.B(n_126),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_180),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_226),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_296),
.C(n_316),
.Y(n_348)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_291),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_175),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_212),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_299),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_209),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_301),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_229),
.Y(n_301)
);

OAI21x1_ASAP7_75t_SL g354 ( 
.A1(n_302),
.A2(n_318),
.B(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_304),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_257),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_306),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_307),
.A2(n_332),
.B1(n_335),
.B2(n_284),
.Y(n_353)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx4_ASAP7_75t_SL g343 ( 
.A(n_308),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_309),
.B(n_331),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_230),
.B(n_218),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_311),
.A2(n_262),
.B(n_261),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_312),
.A2(n_333),
.B1(n_247),
.B2(n_251),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_188),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_313),
.B(n_324),
.Y(n_380)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_317),
.Y(n_370)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_240),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_320),
.B(n_321),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_322),
.B(n_323),
.Y(n_359)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_280),
.B(n_275),
.Y(n_324)
);

INVx13_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_325),
.Y(n_339)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_235),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_326),
.B(n_327),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_204),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_275),
.A2(n_174),
.B1(n_192),
.B2(n_194),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_328),
.A2(n_244),
.B1(n_258),
.B2(n_252),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_279),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_338),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_214),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_242),
.B(n_190),
.Y(n_331)
);

BUFx4f_ASAP7_75t_L g332 ( 
.A(n_255),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_237),
.A2(n_178),
.B1(n_197),
.B2(n_196),
.Y(n_333)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_248),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_334),
.Y(n_356)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_244),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_264),
.B(n_207),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g374 ( 
.A1(n_336),
.A2(n_301),
.B(n_290),
.C(n_292),
.D(n_291),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_276),
.A2(n_217),
.B1(n_234),
.B2(n_8),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_255),
.B1(n_262),
.B2(n_241),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_240),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_349),
.B1(n_362),
.B2(n_381),
.Y(n_384)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_333),
.A2(n_239),
.B1(n_265),
.B2(n_276),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_344),
.Y(n_387)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_300),
.B(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_346),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_318),
.A2(n_266),
.B1(n_245),
.B2(n_254),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_347),
.A2(n_350),
.B1(n_351),
.B2(n_355),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_295),
.A2(n_253),
.B1(n_236),
.B2(n_269),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_318),
.A2(n_286),
.B1(n_253),
.B2(n_251),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_259),
.B1(n_236),
.B2(n_269),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_295),
.A2(n_259),
.B1(n_256),
.B2(n_284),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_302),
.A2(n_256),
.B(n_258),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_363),
.A2(n_330),
.B(n_338),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_252),
.C(n_162),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_365),
.C(n_378),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_289),
.B(n_6),
.C(n_7),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_324),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_377),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_374),
.B(n_346),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_306),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_296),
.B(n_10),
.C(n_11),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_297),
.A2(n_328),
.B1(n_290),
.B2(n_336),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_299),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_312),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_357),
.B(n_298),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_382),
.B(n_415),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_299),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_386),
.A2(n_394),
.B(n_395),
.Y(n_423)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_389),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_397),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_368),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_403),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_340),
.A2(n_349),
.B1(n_362),
.B2(n_369),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_393),
.A2(n_347),
.B1(n_345),
.B2(n_379),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_293),
.Y(n_394)
);

AO22x1_ASAP7_75t_L g395 ( 
.A1(n_354),
.A2(n_311),
.B1(n_321),
.B2(n_305),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_297),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_348),
.C(n_364),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_325),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_376),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_398),
.Y(n_420)
);

O2A1O1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_345),
.A2(n_330),
.B(n_322),
.C(n_314),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_408),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_400),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_315),
.Y(n_401)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_334),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_329),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_404),
.B(n_405),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_357),
.B(n_303),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_407),
.A2(n_339),
.B(n_356),
.Y(n_440)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_409),
.B(n_410),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_339),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_373),
.A2(n_294),
.B(n_323),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_412),
.A2(n_363),
.B(n_359),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_359),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_413),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_346),
.B(n_320),
.Y(n_415)
);

INVx13_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_416),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_305),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_417),
.B(n_370),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_424),
.A2(n_425),
.B1(n_433),
.B2(n_445),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_387),
.A2(n_393),
.B1(n_384),
.B2(n_345),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_434),
.C(n_448),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_387),
.A2(n_350),
.B1(n_377),
.B2(n_372),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_396),
.B(n_352),
.C(n_371),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_435),
.A2(n_440),
.B(n_407),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_409),
.B(n_365),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_437),
.B(n_400),
.Y(n_461)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_390),
.B(n_378),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_415),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_411),
.A2(n_356),
.B(n_375),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_10),
.B(n_12),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_412),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_451),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_384),
.A2(n_351),
.B1(n_355),
.B2(n_370),
.Y(n_445)
);

XOR2x2_ASAP7_75t_L g447 ( 
.A(n_386),
.B(n_367),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_395),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_391),
.B(n_310),
.C(n_361),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_402),
.A2(n_385),
.B1(n_382),
.B2(n_413),
.Y(n_449)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_411),
.A2(n_361),
.B1(n_360),
.B2(n_310),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_450),
.A2(n_402),
.B1(n_408),
.B2(n_388),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_391),
.B(n_307),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_452),
.A2(n_476),
.B1(n_436),
.B2(n_446),
.Y(n_488)
);

XNOR2x1_ASAP7_75t_L g503 ( 
.A(n_454),
.B(n_14),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_389),
.C(n_386),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_464),
.C(n_420),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_443),
.B1(n_425),
.B2(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_457),
.A2(n_479),
.B(n_435),
.Y(n_484)
);

OAI22x1_ASAP7_75t_L g459 ( 
.A1(n_433),
.A2(n_395),
.B1(n_394),
.B2(n_397),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_459),
.A2(n_446),
.B1(n_423),
.B2(n_419),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_461),
.B(n_446),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_426),
.A2(n_418),
.B1(n_417),
.B2(n_401),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_471),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_426),
.A2(n_418),
.B1(n_414),
.B2(n_383),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_398),
.C(n_406),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_474),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_429),
.A2(n_403),
.B1(n_375),
.B2(n_385),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_419),
.A2(n_381),
.B1(n_399),
.B2(n_416),
.Y(n_467)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_467),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_326),
.Y(n_469)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_469),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_304),
.Y(n_470)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_470),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_429),
.A2(n_335),
.B1(n_343),
.B2(n_332),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_438),
.Y(n_473)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_308),
.C(n_319),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_437),
.B(n_319),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_477),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_L g476 ( 
.A1(n_421),
.A2(n_343),
.B1(n_332),
.B2(n_14),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_332),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_432),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_432),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_496),
.C(n_501),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_495),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_442),
.C(n_423),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_491),
.Y(n_508)
);

OAI21xp33_ASAP7_75t_SL g521 ( 
.A1(n_484),
.A2(n_486),
.B(n_503),
.Y(n_521)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_457),
.A2(n_440),
.B(n_431),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_462),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_493),
.B(n_499),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g494 ( 
.A(n_455),
.B(n_431),
.CI(n_430),
.CON(n_494),
.SN(n_494)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_458),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_461),
.B(n_430),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_447),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_453),
.B(n_450),
.C(n_439),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_439),
.C(n_420),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_477),
.B(n_445),
.C(n_436),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_463),
.C(n_474),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_485),
.A2(n_472),
.B1(n_468),
.B2(n_460),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_506),
.A2(n_513),
.B1(n_515),
.B2(n_519),
.Y(n_528)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_492),
.Y(n_507)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_507),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_500),
.Y(n_509)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_512),
.A2(n_494),
.B(n_482),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_489),
.A2(n_472),
.B1(n_459),
.B2(n_466),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_480),
.A2(n_476),
.B1(n_465),
.B2(n_454),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_487),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_471),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_517),
.B(n_488),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_480),
.A2(n_479),
.B1(n_16),
.B2(n_17),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_518),
.A2(n_17),
.B1(n_503),
.B2(n_515),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_483),
.A2(n_15),
.B1(n_17),
.B2(n_502),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_501),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_494),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_491),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_522),
.A2(n_516),
.B(n_518),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_499),
.C(n_514),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_524),
.B(n_529),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_525),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_526),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_498),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_535),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_487),
.C(n_497),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_531),
.B(n_533),
.Y(n_548)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_532),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_497),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_496),
.C(n_495),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_534),
.B(n_511),
.C(n_521),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_484),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_536),
.B(n_533),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_511),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_535),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_538),
.A2(n_506),
.B1(n_513),
.B2(n_522),
.Y(n_540)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_542),
.B(n_550),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_544),
.B(n_546),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_524),
.B(n_531),
.C(n_530),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_545),
.C(n_546),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_541),
.A2(n_534),
.B(n_528),
.Y(n_551)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_551),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_548),
.A2(n_527),
.B(n_523),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_553),
.B(n_557),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_541),
.A2(n_537),
.B1(n_543),
.B2(n_539),
.Y(n_555)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_555),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_549),
.C(n_545),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_558),
.B(n_556),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_562),
.A2(n_563),
.B(n_564),
.Y(n_565)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_561),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_559),
.B(n_554),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_563),
.A2(n_560),
.B(n_556),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_566),
.A2(n_551),
.B(n_552),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_567),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_568),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_565),
.C(n_555),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_570),
.B(n_547),
.Y(n_571)
);


endmodule