module fake_jpeg_25007_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_23),
.B1(n_25),
.B2(n_19),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_46),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_47),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_21),
.B1(n_25),
.B2(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_15),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx10_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_27),
.B1(n_31),
.B2(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

OA21x2_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_44),
.B(n_27),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_73),
.B(n_76),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_55),
.B(n_56),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_34),
.B1(n_41),
.B2(n_32),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_49),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_80),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_52),
.B(n_27),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_85),
.B(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_87),
.B1(n_72),
.B2(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_67),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_31),
.B1(n_39),
.B2(n_41),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_32),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_72),
.B1(n_57),
.B2(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_88),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_54),
.B1(n_32),
.B2(n_30),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_95),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_63),
.B(n_67),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_93),
.B(n_2),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_66),
.A3(n_71),
.B1(n_69),
.B2(n_74),
.C1(n_7),
.C2(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_63),
.B(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_88),
.C(n_79),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_105),
.C(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_28),
.C(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_107),
.B(n_66),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_83),
.B1(n_28),
.B2(n_4),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_95),
.B1(n_93),
.B2(n_98),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_100),
.B(n_102),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_105),
.B1(n_108),
.B2(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_8),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_95),
.C(n_28),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2x1p5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_8),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_119),
.C(n_109),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_113),
.B(n_11),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_118),
.B1(n_3),
.B2(n_2),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_124),
.C(n_2),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_6),
.B(n_7),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_123),
.A2(n_3),
.B(n_14),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_10),
.C(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_14),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_128),
.Y(n_130)
);


endmodule