module fake_jpeg_4591_n_230 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_40),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_44),
.B1(n_28),
.B2(n_23),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_0),
.Y(n_74)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_6),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_15),
.Y(n_66)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_15),
.C(n_30),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_7),
.C(n_11),
.Y(n_117)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_56),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_16),
.B1(n_22),
.B2(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_64),
.B1(n_85),
.B2(n_20),
.Y(n_101)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_16),
.B1(n_22),
.B2(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NAND2x1_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_26),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_2),
.B(n_4),
.C(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_34),
.B(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

AO21x1_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_82),
.B(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_39),
.B(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_32),
.A2(n_26),
.B1(n_1),
.B2(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_33),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_33),
.B(n_18),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_20),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_26),
.B1(n_1),
.B2(n_0),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_102),
.B1(n_50),
.B2(n_75),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_26),
.B(n_3),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_101),
.B(n_64),
.C(n_52),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_86),
.B(n_48),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_80),
.Y(n_126)
);

AOI22x1_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_58),
.A2(n_19),
.B1(n_8),
.B2(n_10),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_113),
.B1(n_72),
.B2(n_11),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_61),
.B1(n_54),
.B2(n_68),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_79),
.B1(n_60),
.B2(n_7),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_108),
.Y(n_143)
);

HAxp5_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_136),
.CON(n_161),
.SN(n_161)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_143),
.Y(n_157)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_123),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_51),
.B1(n_55),
.B2(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_57),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_72),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_126),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_59),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_117),
.B1(n_112),
.B2(n_116),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_145),
.B(n_146),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_142),
.B(n_94),
.C(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_135),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_86),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_49),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_76),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_53),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_91),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_56),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_99),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_106),
.B(n_92),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_97),
.A2(n_94),
.B(n_107),
.Y(n_146)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_168),
.B1(n_162),
.B2(n_160),
.C(n_156),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_170),
.C(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_115),
.B1(n_112),
.B2(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_105),
.B1(n_115),
.B2(n_145),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_130),
.B1(n_123),
.B2(n_118),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_132),
.B(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_168),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_121),
.B(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_137),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_142),
.B1(n_122),
.B2(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_143),
.C(n_146),
.Y(n_172)
);

OA21x2_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_183),
.B(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_177),
.C(n_181),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_139),
.B1(n_131),
.B2(n_120),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_150),
.B(n_159),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_124),
.C(n_132),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_154),
.B(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_157),
.B(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_190),
.C(n_177),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_200),
.Y(n_202)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_148),
.B1(n_168),
.B2(n_161),
.C(n_158),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_194),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

AOI221xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_168),
.B1(n_157),
.B2(n_147),
.C(n_153),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_147),
.B1(n_153),
.B2(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_195),
.A2(n_175),
.B1(n_182),
.B2(n_187),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_178),
.B(n_179),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_176),
.Y(n_201)
);

INVxp33_ASAP7_75t_SL g204 ( 
.A(n_201),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_190),
.B(n_196),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_207),
.B(n_208),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_180),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_186),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_195),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_186),
.B1(n_174),
.B2(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_200),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_206),
.B(n_215),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_193),
.B1(n_204),
.B2(n_201),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_205),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_219),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_211),
.B1(n_198),
.B2(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_207),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_226),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_225),
.Y(n_230)
);


endmodule