module fake_jpeg_31654_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_45),
.B1(n_48),
.B2(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_3),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_60),
.B(n_61),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_44),
.C(n_42),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_68),
.C(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_49),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_40),
.B(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_39),
.B1(n_47),
.B2(n_40),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_5),
.C(n_6),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_4),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_54),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_67),
.C(n_58),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_17),
.B1(n_34),
.B2(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_4),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_5),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_78),
.C(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_6),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_85),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_15),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_68),
.B1(n_58),
.B2(n_9),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_90),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_96),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_7),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_19),
.C(n_24),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_101),
.B1(n_93),
.B2(n_20),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_101)
);

AOI321xp33_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_93),
.A3(n_95),
.B1(n_91),
.B2(n_92),
.C(n_23),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_106),
.C(n_107),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_14),
.B1(n_21),
.B2(n_22),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_102),
.C(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_102),
.C(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_35),
.Y(n_114)
);


endmodule