module fake_jpeg_32124_n_514 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_514);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_514;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_58),
.Y(n_109)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_59),
.B(n_62),
.Y(n_125)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_16),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_89),
.Y(n_157)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_77),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_86),
.Y(n_140)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_30),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_93),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_21),
.B(n_15),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_1),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_101),
.Y(n_160)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_98),
.Y(n_155)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_44),
.Y(n_99)
);

NAND2x1_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_103),
.Y(n_147)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_28),
.B1(n_48),
.B2(n_35),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_108),
.A2(n_110),
.B1(n_156),
.B2(n_159),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_28),
.B1(n_48),
.B2(n_35),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_39),
.B1(n_42),
.B2(n_25),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_111),
.A2(n_121),
.B1(n_135),
.B2(n_143),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_64),
.B(n_39),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_144),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_39),
.B1(n_42),
.B2(n_36),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_60),
.B(n_38),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_124),
.B(n_126),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_38),
.C(n_22),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_91),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_131),
.B1(n_78),
.B2(n_79),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_67),
.A2(n_28),
.B1(n_48),
.B2(n_35),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_72),
.A2(n_42),
.B1(n_36),
.B2(n_20),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_69),
.A2(n_26),
.B(n_47),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g212 ( 
.A(n_137),
.B(n_103),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_81),
.A2(n_36),
.B1(n_20),
.B2(n_48),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_20),
.C(n_35),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_92),
.A2(n_28),
.B1(n_49),
.B2(n_47),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_70),
.A2(n_41),
.B1(n_46),
.B2(n_51),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_97),
.A2(n_49),
.B1(n_51),
.B2(n_32),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_73),
.A2(n_46),
.B1(n_41),
.B2(n_45),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_32),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_163),
.B(n_166),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_61),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_165),
.B(n_171),
.CI(n_200),
.CON(n_257),
.SN(n_257)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_33),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_115),
.A2(n_80),
.B1(n_74),
.B2(n_83),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_167),
.A2(n_212),
.B1(n_71),
.B2(n_130),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_45),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_175),
.Y(n_220)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_33),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_170),
.B(n_180),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_34),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_176),
.Y(n_230)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_186),
.Y(n_250)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_109),
.B(n_34),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_181),
.A2(n_215),
.B1(n_148),
.B2(n_104),
.Y(n_255)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_112),
.A2(n_102),
.B1(n_63),
.B2(n_66),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_185),
.A2(n_211),
.B1(n_55),
.B2(n_57),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_56),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_188),
.B(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_195),
.Y(n_258)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_114),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_133),
.B(n_56),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_198),
.Y(n_259)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_114),
.Y(n_200)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g204 ( 
.A(n_153),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_150),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_100),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_127),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_153),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_134),
.A2(n_87),
.B1(n_76),
.B2(n_95),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_106),
.B(n_119),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_214),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_106),
.B(n_99),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_69),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_104),
.C(n_161),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_232),
.C(n_233),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_200),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_152),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_238),
.B1(n_240),
.B2(n_255),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_165),
.B(n_152),
.C(n_161),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_235),
.A2(n_206),
.B(n_202),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_136),
.B1(n_132),
.B2(n_130),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_136),
.B1(n_132),
.B2(n_112),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_193),
.B1(n_201),
.B2(n_183),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_181),
.A2(n_212),
.B1(n_164),
.B2(n_216),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_224),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_261),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_262),
.A2(n_270),
.B1(n_276),
.B2(n_288),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_165),
.B(n_195),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_242),
.B(n_247),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_168),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_268),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_173),
.B1(n_171),
.B2(n_211),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_267),
.A2(n_242),
.B1(n_225),
.B2(n_149),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_180),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_173),
.B1(n_175),
.B2(n_188),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_184),
.C(n_171),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_272),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_163),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_273),
.A2(n_286),
.B(n_230),
.Y(n_319)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_217),
.A2(n_146),
.B1(n_162),
.B2(n_142),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_223),
.B(n_192),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_277),
.B(n_284),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_169),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_281),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_279),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_251),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_280),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_177),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_210),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_176),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_227),
.A2(n_148),
.B1(n_190),
.B2(n_197),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_182),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_295),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_235),
.A2(n_257),
.B1(n_254),
.B2(n_234),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_259),
.A2(n_174),
.B1(n_189),
.B2(n_146),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_294),
.B1(n_225),
.B2(n_253),
.Y(n_317)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_228),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_297),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_187),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_256),
.B(n_252),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_254),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_257),
.A2(n_145),
.B1(n_149),
.B2(n_107),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_231),
.B(n_194),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_199),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_298),
.Y(n_325)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_229),
.B(n_208),
.Y(n_298)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_267),
.A2(n_196),
.B1(n_241),
.B2(n_145),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_302),
.A2(n_314),
.B1(n_320),
.B2(n_332),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_303),
.A2(n_319),
.B(n_286),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_247),
.C(n_219),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_274),
.Y(n_335)
);

AND2x2_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_243),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_305),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_307),
.B(n_327),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_323),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_256),
.C(n_252),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_273),
.C(n_276),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_317),
.A2(n_330),
.B1(n_266),
.B2(n_278),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_265),
.A2(n_205),
.B1(n_196),
.B2(n_218),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_293),
.B(n_222),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_288),
.B(n_237),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_331),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_298),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_268),
.B(n_253),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_329),
.B(n_289),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_270),
.A2(n_218),
.B1(n_245),
.B2(n_236),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_281),
.B(n_237),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_265),
.A2(n_245),
.B1(n_230),
.B2(n_221),
.Y(n_332)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_352),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_345),
.C(n_350),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_338),
.A2(n_319),
.B(n_314),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_346),
.Y(n_380)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_284),
.C(n_277),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_351),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_264),
.C(n_263),
.Y(n_345)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_348),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_294),
.C(n_292),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g351 ( 
.A(n_306),
.Y(n_351)
);

A2O1A1O1Ixp25_ASAP7_75t_L g352 ( 
.A1(n_306),
.A2(n_292),
.B(n_271),
.C(n_269),
.D(n_283),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_357),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_326),
.A2(n_262),
.B1(n_297),
.B2(n_291),
.Y(n_355)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_290),
.Y(n_356)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_296),
.C(n_280),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_309),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_358),
.B(n_362),
.Y(n_372)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_302),
.A2(n_279),
.B1(n_261),
.B2(n_295),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_361),
.A2(n_317),
.B1(n_330),
.B2(n_323),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_299),
.B(n_226),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_299),
.B(n_221),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_363),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_304),
.B(n_311),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_367),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_275),
.Y(n_366)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_366),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_311),
.B(n_226),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_303),
.B(n_308),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_377),
.A2(n_381),
.B(n_384),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_305),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_391),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_382),
.A2(n_386),
.B1(n_360),
.B2(n_361),
.Y(n_409)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_338),
.A2(n_316),
.B(n_301),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_331),
.C(n_324),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_388),
.C(n_393),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_364),
.A2(n_308),
.B1(n_332),
.B2(n_320),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_336),
.B(n_305),
.C(n_310),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_344),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_337),
.A2(n_343),
.B(n_308),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_392),
.B(n_360),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_305),
.C(n_310),
.Y(n_393)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_396),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_327),
.Y(n_399)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_399),
.Y(n_425)
);

OAI21xp33_ASAP7_75t_L g400 ( 
.A1(n_395),
.A2(n_354),
.B(n_352),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_400),
.Y(n_427)
);

FAx1_ASAP7_75t_SL g402 ( 
.A(n_397),
.B(n_344),
.CI(n_367),
.CON(n_402),
.SN(n_402)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_408),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_397),
.B(n_385),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_406),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_391),
.B(n_301),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_316),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_409),
.A2(n_418),
.B1(n_422),
.B2(n_387),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_325),
.C(n_312),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_412),
.C(n_416),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_312),
.C(n_315),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_414),
.Y(n_430)
);

AO21x1_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_282),
.B(n_2),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_315),
.C(n_333),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_370),
.C(n_393),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_417),
.A2(n_420),
.B(n_421),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_333),
.B1(n_322),
.B2(n_348),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_368),
.Y(n_419)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_419),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_322),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_381),
.A2(n_384),
.B1(n_396),
.B2(n_373),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_383),
.Y(n_423)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_423),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_414),
.A2(n_373),
.B1(n_371),
.B2(n_380),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_426),
.A2(n_429),
.B1(n_437),
.B2(n_440),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_421),
.A2(n_380),
.B1(n_392),
.B2(n_377),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_SL g432 ( 
.A1(n_413),
.A2(n_398),
.B(n_390),
.C(n_378),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_432),
.A2(n_434),
.B(n_439),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_433),
.A2(n_405),
.B1(n_401),
.B2(n_418),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_413),
.A2(n_398),
.B(n_378),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_424),
.A2(n_341),
.B1(n_342),
.B2(n_394),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_SL g438 ( 
.A(n_403),
.B(n_406),
.C(n_404),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_438),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_422),
.A2(n_341),
.B(n_321),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_410),
.A2(n_282),
.B1(n_2),
.B2(n_3),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_442),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_409),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_442)
);

OAI322xp33_ASAP7_75t_L g445 ( 
.A1(n_399),
.A2(n_43),
.A3(n_31),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_445)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_445),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_443),
.B(n_416),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_460),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_412),
.C(n_411),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_452),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_404),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_455),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_420),
.Y(n_454)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_417),
.C(n_407),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_426),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_459),
.Y(n_471)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_437),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_407),
.C(n_402),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_444),
.B(n_402),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_440),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_462),
.A2(n_439),
.B1(n_434),
.B2(n_431),
.Y(n_465)
);

XOR2x2_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_432),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_464),
.A2(n_452),
.B(n_450),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_472),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_460),
.B(n_436),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_473),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_449),
.A2(n_432),
.B1(n_441),
.B2(n_429),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_468),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_488)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_454),
.A2(n_432),
.B(n_428),
.Y(n_469)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_428),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_31),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_474),
.B(n_475),
.C(n_450),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_31),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_451),
.A2(n_2),
.B(n_5),
.Y(n_478)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_480),
.B(n_486),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_483),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_477),
.B(n_448),
.Y(n_483)
);

O2A1O1Ixp33_ASAP7_75t_SL g484 ( 
.A1(n_464),
.A2(n_468),
.B(n_471),
.C(n_463),
.Y(n_484)
);

O2A1O1Ixp33_ASAP7_75t_SL g495 ( 
.A1(n_484),
.A2(n_491),
.B(n_10),
.C(n_12),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_446),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_476),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_447),
.B(n_7),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_488),
.B(n_489),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_474),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_470),
.A2(n_10),
.B(n_12),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_466),
.C(n_475),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_494),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_495),
.A2(n_488),
.B(n_490),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_31),
.C(n_43),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_498),
.B(n_499),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_31),
.C(n_13),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_31),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_497),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_493),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_503),
.A2(n_496),
.B(n_486),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_496),
.A2(n_480),
.B(n_484),
.Y(n_504)
);

AO21x1_ASAP7_75t_L g509 ( 
.A1(n_504),
.A2(n_506),
.B(n_481),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_505),
.B(n_489),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_508),
.Y(n_511)
);

AO21x1_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_501),
.B(n_502),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_511),
.C(n_13),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_14),
.B(n_12),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_13),
.Y(n_514)
);


endmodule