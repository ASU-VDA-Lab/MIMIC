module fake_jpeg_10745_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_62),
.Y(n_71)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_40),
.B1(n_51),
.B2(n_48),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_71),
.B(n_52),
.C(n_68),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_50),
.B(n_46),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_11),
.B(n_12),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_90),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_42),
.B1(n_51),
.B2(n_45),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_88),
.B(n_10),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_85),
.B1(n_14),
.B2(n_17),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_0),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_52),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_89),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_70),
.B1(n_2),
.B2(n_4),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_4),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_5),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_13),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_5),
.B(n_7),
.C(n_9),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_107),
.B1(n_21),
.B2(n_23),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_115),
.B(n_114),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_97),
.B(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_104),
.C(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_119),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_120),
.B(n_109),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_109),
.A3(n_99),
.B1(n_116),
.B2(n_108),
.C1(n_93),
.C2(n_34),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_24),
.C(n_27),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_113),
.Y(n_127)
);


endmodule