module fake_jpeg_17083_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_27),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_25),
.B1(n_21),
.B2(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_2),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_51),
.Y(n_99)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_20),
.A2(n_3),
.B(n_5),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_52),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_11),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_5),
.B(n_6),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_55),
.B(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_23),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_7),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_10),
.C(n_11),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_72),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_30),
.B1(n_21),
.B2(n_23),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_67),
.A2(n_102),
.B(n_82),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_68),
.A2(n_88),
.B1(n_17),
.B2(n_99),
.Y(n_123)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_100),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_96),
.Y(n_128)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_39),
.A2(n_35),
.B1(n_34),
.B2(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_60),
.B1(n_35),
.B2(n_42),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_83),
.Y(n_120)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_19),
.B1(n_32),
.B2(n_34),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_24),
.Y(n_117)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_97),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_34),
.B1(n_35),
.B2(n_24),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_122),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_105),
.A2(n_123),
.B1(n_118),
.B2(n_125),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_24),
.B1(n_17),
.B2(n_10),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_73),
.B(n_75),
.Y(n_143)
);

OR2x4_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_29),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_112),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_45),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_110),
.B(n_117),
.Y(n_157)
);

FAx1_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_29),
.CI(n_16),
.CON(n_112),
.SN(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_10),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_121),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_16),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_133),
.B1(n_108),
.B2(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_64),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_130),
.Y(n_151)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_77),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_67),
.B1(n_92),
.B2(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_70),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_66),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_73),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_146),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_119),
.B(n_120),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_133),
.B1(n_105),
.B2(n_127),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_142),
.B1(n_139),
.B2(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_121),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_110),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_118),
.C(n_115),
.Y(n_174)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_111),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_157),
.B1(n_143),
.B2(n_151),
.C(n_160),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_138),
.B(n_150),
.Y(n_186)
);

NOR4xp25_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_149),
.C(n_158),
.D(n_136),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_136),
.B(n_156),
.C(n_157),
.D(n_140),
.Y(n_187)
);

XOR2x2_ASAP7_75t_SL g169 ( 
.A(n_153),
.B(n_118),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_103),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_125),
.C(n_122),
.Y(n_179)
);

NOR4xp25_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_130),
.C(n_159),
.D(n_152),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_169),
.B(n_164),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_120),
.C(n_122),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_155),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_183),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_198),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_187),
.B(n_189),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_180),
.A2(n_153),
.B1(n_147),
.B2(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

OAI22x1_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_197),
.B1(n_199),
.B2(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_177),
.C(n_172),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_167),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_161),
.B(n_104),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_171),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_174),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_205),
.C(n_206),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_177),
.C(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_209),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_176),
.B1(n_196),
.B2(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_171),
.C(n_165),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_162),
.C(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_185),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_176),
.Y(n_212)
);

AOI321xp33_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_176),
.A3(n_186),
.B1(n_180),
.B2(n_199),
.C(n_187),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_217),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_220),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_202),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_211),
.C(n_190),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_206),
.C(n_200),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_216),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_208),
.C(n_201),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_212),
.B(n_214),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_113),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_231),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_195),
.B(n_192),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_226),
.A2(n_113),
.B1(n_163),
.B2(n_222),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_233),
.A2(n_227),
.B(n_229),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_235),
.B(n_236),
.CI(n_233),
.CON(n_237),
.SN(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_228),
.C(n_232),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_236),
.Y(n_238)
);


endmodule