module fake_jpeg_21973_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_19),
.A2(n_22),
.B1(n_24),
.B2(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_6),
.B(n_7),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_9),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_33),
.B(n_35),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_32),
.B1(n_27),
.B2(n_29),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_21),
.B(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_15),
.B1(n_18),
.B2(n_7),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_26),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_42),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_44),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_31),
.B(n_29),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_20),
.B(n_7),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_49),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_50),
.B1(n_38),
.B2(n_42),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_54),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_48),
.B(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_55),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_34),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_53),
.C(n_43),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_60),
.C(n_41),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_41),
.C(n_46),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_56),
.B(n_34),
.Y(n_62)
);


endmodule