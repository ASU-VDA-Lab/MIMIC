module fake_jpeg_16428_n_213 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_213);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_52),
.B1(n_55),
.B2(n_19),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_18),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_20),
.B1(n_34),
.B2(n_17),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_60),
.Y(n_90)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_34),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_71),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_17),
.B1(n_34),
.B2(n_27),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_22),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_21),
.B1(n_32),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_84),
.B1(n_85),
.B2(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_82),
.B1(n_88),
.B2(n_92),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_22),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_26),
.B1(n_32),
.B2(n_23),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_93),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_30),
.B1(n_31),
.B2(n_19),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_43),
.C(n_45),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_19),
.C(n_30),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_30),
.B1(n_19),
.B2(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_53),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_19),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_24),
.B(n_6),
.C(n_7),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_115),
.B1(n_119),
.B2(n_109),
.Y(n_128)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_111),
.B(n_106),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_4),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_83),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_103),
.C(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_82),
.C(n_68),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_127),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_79),
.B1(n_96),
.B2(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_131),
.B1(n_137),
.B2(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_119),
.B1(n_102),
.B2(n_99),
.Y(n_145)
);

NAND2xp67_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_84),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_133),
.B(n_141),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_85),
.B1(n_75),
.B2(n_77),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_95),
.B(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_115),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_80),
.B1(n_89),
.B2(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_78),
.B(n_7),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_5),
.B1(n_7),
.B2(n_24),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_149),
.B1(n_158),
.B2(n_157),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_97),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_156),
.B(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_153),
.Y(n_162)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_116),
.C(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_104),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_143),
.A3(n_146),
.B1(n_152),
.B2(n_144),
.C1(n_148),
.C2(n_151),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_160),
.A2(n_133),
.B(n_122),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_169),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_138),
.B1(n_140),
.B2(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_173),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_140),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_160),
.A2(n_112),
.B(n_141),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_100),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_147),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g178 ( 
.A1(n_174),
.A2(n_147),
.B(n_150),
.Y(n_178)
);

OAI322xp33_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_179),
.A3(n_173),
.B1(n_169),
.B2(n_172),
.C1(n_171),
.C2(n_24),
.Y(n_190)
);

OA21x2_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_159),
.B(n_145),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_183),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_165),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_16),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_156),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_24),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_186),
.A2(n_167),
.B1(n_175),
.B2(n_170),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_161),
.B1(n_179),
.B2(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_183),
.Y(n_196)
);

AOI31xp33_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_181),
.A3(n_16),
.B(n_14),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_24),
.B(n_10),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_194),
.B(n_13),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_24),
.B1(n_10),
.B2(n_11),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_193),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_9),
.B(n_11),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_201),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_192),
.B(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_195),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.C(n_206),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_187),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_193),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_176),
.B1(n_182),
.B2(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_206),
.B(n_198),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_208),
.B(n_176),
.CI(n_198),
.CON(n_210),
.SN(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_209),
.B(n_211),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_210),
.Y(n_213)
);


endmodule