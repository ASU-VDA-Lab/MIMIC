module fake_netlist_1_11737_n_694 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_694);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_694;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_446;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_631;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_56), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_47), .Y(n_79) );
BUFx6f_ASAP7_75t_L g80 ( .A(n_6), .Y(n_80) );
INVx1_ASAP7_75t_SL g81 ( .A(n_3), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_36), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_29), .Y(n_83) );
OR2x2_ASAP7_75t_L g84 ( .A(n_65), .B(n_40), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_14), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_49), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_33), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_11), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_31), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_59), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_53), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_30), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g95 ( .A(n_4), .B(n_1), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_55), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_4), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_21), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_3), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_13), .Y(n_101) );
XNOR2xp5_ASAP7_75t_L g102 ( .A(n_22), .B(n_10), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_37), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_42), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_1), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_67), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_73), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_0), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_12), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_20), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_9), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_66), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_50), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_43), .Y(n_119) );
BUFx8_ASAP7_75t_SL g120 ( .A(n_51), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_34), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_28), .Y(n_122) );
BUFx5_ASAP7_75t_L g123 ( .A(n_58), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_25), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_111), .B(n_0), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_100), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_100), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
OR2x2_ASAP7_75t_L g129 ( .A(n_89), .B(n_2), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_123), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_82), .B(n_5), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_78), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_123), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_123), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_84), .B(n_39), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_103), .B(n_5), .Y(n_138) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_92), .B(n_77), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_103), .B(n_41), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_80), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_123), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_80), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_123), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_107), .B(n_6), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_120), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_119), .B(n_7), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_80), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_88), .B(n_8), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_90), .B(n_44), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_111), .B(n_8), .Y(n_158) );
CKINVDCx16_ASAP7_75t_R g159 ( .A(n_118), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_113), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_91), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_98), .B(n_10), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_97), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_123), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_104), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_116), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_122), .Y(n_169) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_125), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_157), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_131), .Y(n_173) );
NAND2xp33_ASAP7_75t_SL g174 ( .A(n_148), .B(n_124), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_159), .B(n_98), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_128), .B(n_113), .Y(n_180) );
OR2x6_ASAP7_75t_L g181 ( .A(n_129), .B(n_95), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_159), .B(n_110), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_128), .B(n_109), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_128), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_152), .B(n_114), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_131), .A2(n_105), .B1(n_86), .B2(n_117), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_131), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_152), .B(n_81), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
AND2x6_ASAP7_75t_L g192 ( .A(n_147), .B(n_115), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_152), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_147), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_151), .B(n_108), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
NOR2xp33_ASAP7_75t_SL g200 ( .A(n_139), .B(n_120), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_129), .B(n_106), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_132), .B(n_99), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_132), .B(n_94), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_151), .B(n_102), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_137), .B(n_124), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_151), .B(n_94), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_137), .B(n_112), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_142), .B(n_112), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_138), .B(n_101), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_142), .B(n_101), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_138), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_157), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_161), .B(n_46), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_161), .B(n_45), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_162), .B(n_11), .Y(n_220) );
BUFx4f_ASAP7_75t_L g221 ( .A(n_139), .Y(n_221) );
OAI22xp33_ASAP7_75t_SL g222 ( .A1(n_158), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_162), .B(n_168), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_164), .B(n_52), .Y(n_224) );
AO22x2_ASAP7_75t_L g225 ( .A1(n_164), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_166), .B(n_168), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_150), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_175), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_170), .B(n_166), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_172), .B(n_135), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_226), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_175), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_214), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_226), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_180), .B(n_135), .Y(n_235) );
INVxp67_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_181), .B(n_208), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_226), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_172), .B(n_135), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_192), .A2(n_157), .B1(n_167), .B2(n_156), .Y(n_241) );
NAND2x1_ASAP7_75t_L g242 ( .A(n_192), .B(n_157), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_192), .A2(n_157), .B1(n_167), .B2(n_163), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_172), .B(n_144), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_214), .B(n_144), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_220), .B(n_134), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_196), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_186), .B(n_157), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_204), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_200), .A2(n_157), .B1(n_169), .B2(n_155), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_186), .B(n_223), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_220), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
OAI22xp5_ASAP7_75t_SL g256 ( .A1(n_181), .A2(n_126), .B1(n_127), .B2(n_155), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_188), .B(n_126), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_190), .B(n_127), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_176), .A2(n_146), .B1(n_165), .B2(n_133), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_181), .B(n_178), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_224), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_173), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_192), .B(n_146), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_176), .A2(n_169), .B1(n_155), .B2(n_140), .Y(n_264) );
NOR2x2_ASAP7_75t_L g265 ( .A(n_174), .B(n_221), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_213), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_204), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_173), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_192), .A2(n_169), .B1(n_155), .B2(n_140), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_198), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_184), .B(n_169), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_198), .B(n_130), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_173), .B(n_130), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_198), .B(n_133), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_198), .B(n_149), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_179), .A2(n_149), .B(n_165), .Y(n_276) );
NOR2x2_ASAP7_75t_L g277 ( .A(n_174), .B(n_134), .Y(n_277) );
OR2x6_ASAP7_75t_L g278 ( .A(n_177), .B(n_169), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_213), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_187), .B(n_153), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_198), .A2(n_140), .B1(n_153), .B2(n_150), .Y(n_281) );
NOR2xp67_ASAP7_75t_L g282 ( .A(n_185), .B(n_145), .Y(n_282) );
CKINVDCx14_ASAP7_75t_R g283 ( .A(n_182), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_202), .B(n_140), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_202), .B(n_203), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_221), .A2(n_140), .B1(n_153), .B2(n_150), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_213), .A2(n_140), .B1(n_153), .B2(n_145), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_211), .B(n_153), .Y(n_288) );
NOR3xp33_ASAP7_75t_L g289 ( .A(n_205), .B(n_145), .C(n_143), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_188), .B(n_140), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_254), .A2(n_199), .B1(n_189), .B2(n_191), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_237), .B(n_210), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_235), .A2(n_197), .B(n_194), .C(n_215), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_244), .A2(n_193), .B(n_207), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_236), .B(n_205), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_260), .B(n_183), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_285), .A2(n_210), .B(n_207), .C(n_229), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_283), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_244), .A2(n_193), .B(n_216), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_253), .B(n_206), .Y(n_303) );
NOR2xp33_ASAP7_75t_SL g304 ( .A(n_270), .B(n_224), .Y(n_304) );
AO32x1_ASAP7_75t_L g305 ( .A1(n_259), .A2(n_225), .A3(n_218), .B1(n_219), .B2(n_224), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_283), .B(n_212), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_258), .A2(n_201), .B(n_222), .C(n_215), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_230), .A2(n_216), .B(n_218), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_270), .B(n_227), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_SL g310 ( .A1(n_242), .A2(n_224), .B(n_143), .C(n_141), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_235), .B(n_16), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_261), .B(n_227), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_234), .B(n_143), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_255), .A2(n_141), .B(n_225), .C(n_154), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_257), .B(n_225), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_230), .A2(n_227), .B(n_217), .Y(n_316) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_255), .A2(n_141), .B(n_154), .C(n_171), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_239), .A2(n_227), .B(n_217), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_257), .B(n_154), .Y(n_319) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_276), .A2(n_154), .B(n_217), .C(n_171), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_278), .B(n_154), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_257), .B(n_217), .Y(n_322) );
OAI21xp33_ASAP7_75t_L g323 ( .A1(n_238), .A2(n_171), .B(n_19), .Y(n_323) );
XOR2x2_ASAP7_75t_L g324 ( .A(n_289), .B(n_18), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_239), .A2(n_171), .B(n_24), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_278), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_247), .A2(n_23), .B(n_27), .C(n_32), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_262), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_278), .B(n_35), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_250), .A2(n_38), .B(n_48), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_268), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_290), .B(n_54), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_261), .B(n_57), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_290), .B(n_61), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_247), .A2(n_246), .B(n_273), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_290), .B(n_62), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_246), .A2(n_64), .B(n_68), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_266), .A2(n_69), .B(n_70), .C(n_72), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_268), .B(n_74), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_233), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_261), .B(n_75), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_279), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_282), .B(n_76), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_256), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_300), .A2(n_271), .B(n_280), .C(n_288), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_SL g346 ( .A1(n_314), .A2(n_284), .B(n_291), .C(n_252), .Y(n_346) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_303), .A2(n_273), .B(n_288), .C(n_271), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_SL g348 ( .A1(n_295), .A2(n_291), .B(n_275), .C(n_274), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_294), .B(n_261), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_316), .A2(n_286), .B(n_264), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_294), .A2(n_241), .B1(n_243), .B2(n_280), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_293), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_301), .Y(n_353) );
CKINVDCx6p67_ASAP7_75t_R g354 ( .A(n_343), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g355 ( .A1(n_307), .A2(n_263), .B(n_272), .C(n_269), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_318), .A2(n_233), .B(n_281), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_342), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_299), .A2(n_233), .B1(n_287), .B2(n_265), .Y(n_358) );
AO31x2_ASAP7_75t_L g359 ( .A1(n_315), .A2(n_228), .A3(n_232), .B(n_267), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_344), .B(n_233), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_297), .A2(n_277), .B1(n_232), .B2(n_240), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_311), .A2(n_228), .B(n_240), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_SL g364 ( .A1(n_338), .A2(n_245), .B(n_248), .C(n_249), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_313), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_308), .A2(n_267), .B(n_248), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_334), .A2(n_245), .B(n_249), .C(n_251), .Y(n_367) );
AO31x2_ASAP7_75t_L g368 ( .A1(n_320), .A2(n_251), .A3(n_319), .B(n_322), .Y(n_368) );
AO21x2_ASAP7_75t_L g369 ( .A1(n_323), .A2(n_332), .B(n_325), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_306), .B(n_326), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_298), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_331), .B(n_328), .Y(n_372) );
BUFx10_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
AO31x2_ASAP7_75t_L g374 ( .A1(n_292), .A2(n_336), .A3(n_330), .B(n_317), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_SL g375 ( .A1(n_333), .A2(n_341), .B(n_339), .C(n_312), .Y(n_375) );
NOR2xp67_ASAP7_75t_SL g376 ( .A(n_340), .B(n_331), .Y(n_376) );
BUFx12f_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
OA21x2_ASAP7_75t_L g378 ( .A1(n_350), .A2(n_337), .B(n_302), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_357), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_346), .A2(n_304), .B(n_310), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_364), .A2(n_304), .B(n_335), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_359), .Y(n_382) );
BUFx12f_ASAP7_75t_L g383 ( .A(n_377), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_352), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_348), .A2(n_305), .B(n_296), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_356), .A2(n_327), .B(n_309), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_361), .B(n_324), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_370), .B(n_292), .Y(n_388) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_365), .A2(n_305), .B(n_321), .C(n_358), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_359), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_359), .Y(n_392) );
CKINVDCx12_ASAP7_75t_R g393 ( .A(n_353), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_354), .B(n_305), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_373), .A2(n_360), .B1(n_349), .B2(n_351), .Y(n_395) );
AO31x2_ASAP7_75t_L g396 ( .A1(n_345), .A2(n_367), .A3(n_366), .B(n_368), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_360), .B(n_373), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_355), .A2(n_347), .B(n_368), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_368), .A2(n_369), .B(n_371), .Y(n_399) );
A2O1A1Ixp33_ASAP7_75t_L g400 ( .A1(n_363), .A2(n_372), .B(n_376), .C(n_362), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_375), .A2(n_369), .B(n_363), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_362), .B(n_372), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_362), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_374), .B(n_294), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_374), .B(n_294), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_388), .A2(n_387), .B1(n_379), .B2(n_384), .C(n_405), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_404), .B(n_391), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_379), .B(n_384), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_402), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_391), .B(n_392), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_401), .A2(n_398), .B(n_399), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_383), .A2(n_394), .B1(n_392), .B2(n_397), .Y(n_414) );
OR2x6_ASAP7_75t_L g415 ( .A(n_402), .B(n_400), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_399), .B(n_396), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_396), .B(n_398), .Y(n_417) );
OR2x6_ASAP7_75t_L g418 ( .A(n_380), .B(n_385), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_396), .B(n_403), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_403), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_390), .B(n_395), .Y(n_421) );
OA21x2_ASAP7_75t_L g422 ( .A1(n_381), .A2(n_386), .B(n_396), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_396), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_389), .A2(n_386), .B(n_378), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_390), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_378), .B(n_383), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_378), .B(n_393), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_378), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_382), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_391), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_379), .B(n_384), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
OR2x6_ASAP7_75t_L g435 ( .A(n_402), .B(n_382), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_391), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
OR2x6_ASAP7_75t_L g438 ( .A(n_402), .B(n_382), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_379), .B(n_384), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_407), .B(n_419), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_410), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_407), .B(n_419), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_435), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_435), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_432), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_406), .B(n_439), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_407), .B(n_412), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_432), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_436), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_411), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_430), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_412), .B(n_439), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_430), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_412), .B(n_408), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_429), .B(n_426), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_419), .B(n_416), .Y(n_460) );
INVx4_ASAP7_75t_L g461 ( .A(n_435), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_416), .B(n_417), .Y(n_462) );
OAI33xp33_ASAP7_75t_L g463 ( .A1(n_436), .A2(n_420), .A3(n_429), .B1(n_423), .B2(n_431), .B3(n_430), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_431), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_427), .B(n_426), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_429), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_427), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_408), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_433), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_416), .B(n_417), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_417), .B(n_420), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_406), .B(n_421), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_435), .B(n_438), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_423), .B(n_421), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_423), .B(n_428), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_428), .B(n_438), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_435), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_425), .A2(n_414), .B1(n_415), .B2(n_438), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_435), .B(n_438), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_438), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_438), .B(n_424), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_424), .B(n_415), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_437), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_409), .B(n_437), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_476), .B(n_415), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_440), .B(n_415), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_476), .B(n_415), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_460), .B(n_415), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_460), .B(n_409), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_441), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_460), .B(n_409), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_462), .B(n_409), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_447), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_444), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_470), .B(n_472), .Y(n_501) );
NOR3xp33_ASAP7_75t_SL g502 ( .A(n_475), .B(n_414), .C(n_425), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_440), .B(n_437), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_467), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_451), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_462), .B(n_434), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_476), .B(n_437), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_470), .B(n_434), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_461), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_440), .B(n_434), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_462), .B(n_434), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_473), .B(n_422), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_454), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_452), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_452), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_471), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_471), .B(n_422), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_459), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_456), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_448), .B(n_418), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_476), .B(n_418), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_473), .B(n_422), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_464), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_442), .B(n_450), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_461), .B(n_413), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_464), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_456), .Y(n_530) );
BUFx2_ASAP7_75t_L g531 ( .A(n_469), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_442), .B(n_422), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_442), .B(n_422), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_445), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_458), .Y(n_536) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_468), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_482), .B(n_418), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_445), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_450), .B(n_413), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_445), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_448), .B(n_418), .Y(n_542) );
INVx4_ASAP7_75t_L g543 ( .A(n_461), .Y(n_543) );
INVx4_ASAP7_75t_L g544 ( .A(n_461), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_543), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_518), .B(n_475), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_527), .B(n_458), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_520), .B(n_474), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_527), .B(n_466), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_530), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_522), .B(n_536), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_493), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_501), .B(n_474), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_493), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_531), .B(n_481), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_497), .B(n_477), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_521), .B(n_491), .Y(n_558) );
OR2x6_ASAP7_75t_L g559 ( .A(n_543), .B(n_443), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_499), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_491), .B(n_466), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_531), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_505), .B(n_477), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_533), .B(n_465), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_499), .B(n_478), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_500), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_533), .B(n_457), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_534), .B(n_457), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_492), .B(n_485), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_500), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_492), .B(n_485), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_494), .B(n_485), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_515), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_495), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_543), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_534), .B(n_457), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_504), .B(n_455), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_506), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_494), .B(n_484), .Y(n_581) );
OAI32xp33_ASAP7_75t_L g582 ( .A1(n_489), .A2(n_480), .A3(n_483), .B1(n_468), .B2(n_482), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_519), .Y(n_583) );
NAND2x1_ASAP7_75t_L g584 ( .A(n_544), .B(n_443), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_506), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_504), .B(n_455), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_512), .B(n_455), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_512), .B(n_449), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_498), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_540), .B(n_449), .Y(n_590) );
CKINVDCx16_ASAP7_75t_R g591 ( .A(n_544), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_498), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_502), .B(n_487), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_488), .B(n_483), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_544), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_540), .B(n_489), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_547), .B(n_525), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_549), .B(n_525), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_562), .B(n_542), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_581), .B(n_514), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_562), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_591), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_564), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_571), .B(n_514), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_545), .B(n_511), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_583), .B(n_523), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_563), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_573), .B(n_507), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_569), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_583), .B(n_508), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_550), .B(n_510), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_555), .A2(n_516), .B(n_517), .C(n_528), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_596), .B(n_508), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_546), .B(n_496), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_574), .B(n_496), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_570), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_566), .A2(n_537), .B(n_528), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_578), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_558), .B(n_516), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_556), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_546), .A2(n_513), .B1(n_507), .B2(n_488), .C(n_490), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_590), .B(n_513), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_561), .B(n_538), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_566), .B(n_529), .Y(n_624) );
OAI32xp33_ASAP7_75t_L g625 ( .A1(n_545), .A2(n_511), .A3(n_528), .B1(n_532), .B2(n_529), .Y(n_625) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_554), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_560), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_575), .B(n_526), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_568), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_575), .B(n_526), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_572), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_565), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_576), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_598), .B(n_551), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_602), .A2(n_593), .B(n_582), .C(n_577), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_624), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_609), .B(n_553), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_628), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_612), .A2(n_595), .B(n_563), .C(n_554), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_599), .A2(n_594), .B1(n_488), .B2(n_490), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_630), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_610), .Y(n_642) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_601), .A2(n_559), .B(n_511), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_621), .A2(n_594), .B1(n_490), .B2(n_548), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_613), .B(n_553), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_626), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_607), .A2(n_548), .B1(n_557), .B2(n_567), .C(n_580), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_610), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_606), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_603), .B(n_557), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_603), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_619), .A2(n_538), .B1(n_524), .B2(n_509), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_620), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_613), .Y(n_654) );
OAI21xp33_ASAP7_75t_SL g655 ( .A1(n_605), .A2(n_559), .B(n_567), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_598), .B(n_604), .Y(n_656) );
AO22x1_ASAP7_75t_L g657 ( .A1(n_655), .A2(n_617), .B1(n_604), .B2(n_600), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_653), .Y(n_658) );
AOI322xp5_ASAP7_75t_L g659 ( .A1(n_649), .A2(n_600), .A3(n_597), .B1(n_608), .B2(n_615), .C1(n_614), .C2(n_623), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_647), .B(n_629), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_644), .A2(n_611), .B1(n_623), .B2(n_524), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g662 ( .A1(n_636), .A2(n_620), .B1(n_629), .B2(n_627), .C1(n_631), .C2(n_625), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_637), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_645), .Y(n_664) );
NAND4xp75_ASAP7_75t_L g665 ( .A(n_640), .B(n_608), .C(n_615), .D(n_627), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_635), .A2(n_625), .B(n_584), .Y(n_666) );
AO21x1_ASAP7_75t_L g667 ( .A1(n_639), .A2(n_585), .B(n_622), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_635), .A2(n_524), .B1(n_616), .B2(n_618), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_638), .B(n_618), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_639), .A2(n_559), .B(n_616), .Y(n_670) );
AOI311xp33_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_641), .A3(n_646), .B(n_651), .C(n_648), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_657), .A2(n_643), .B(n_654), .C(n_652), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_667), .A2(n_642), .B1(n_650), .B2(n_656), .C(n_634), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_660), .A2(n_622), .B1(n_632), .B2(n_633), .C(n_552), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_666), .A2(n_633), .B1(n_632), .B2(n_592), .C(n_589), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_SL g676 ( .A1(n_668), .A2(n_486), .B(n_480), .C(n_532), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_659), .B(n_592), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_663), .A2(n_589), .B1(n_538), .B2(n_463), .C(n_509), .Y(n_678) );
NAND5xp2_ASAP7_75t_L g679 ( .A(n_671), .B(n_662), .C(n_661), .D(n_664), .E(n_665), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_672), .A2(n_662), .B1(n_669), .B2(n_658), .C(n_446), .Y(n_680) );
AND3x2_ASAP7_75t_L g681 ( .A(n_673), .B(n_446), .C(n_509), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_675), .A2(n_588), .B(n_587), .C(n_579), .Y(n_682) );
NOR2x1_ASAP7_75t_L g683 ( .A(n_677), .B(n_486), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_682), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_683), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_680), .A2(n_679), .B(n_678), .C(n_674), .Y(n_686) );
OA22x2_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_681), .B1(n_676), .B2(n_483), .Y(n_687) );
INVx4_ASAP7_75t_L g688 ( .A(n_685), .Y(n_688) );
BUFx2_ASAP7_75t_SL g689 ( .A(n_688), .Y(n_689) );
NAND4xp75_ASAP7_75t_L g690 ( .A(n_689), .B(n_684), .C(n_685), .D(n_687), .Y(n_690) );
AOI222xp33_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_463), .B1(n_487), .B2(n_484), .C1(n_479), .C2(n_468), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_691), .Y(n_692) );
AO221x1_ASAP7_75t_L g693 ( .A1(n_692), .A2(n_541), .B1(n_539), .B2(n_535), .C(n_453), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_487), .B(n_586), .Y(n_694) );
endmodule