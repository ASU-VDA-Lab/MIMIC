module real_jpeg_20018_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_304, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_304;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_299;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_244;
wire n_216;
wire n_133;
wire n_213;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_0),
.A2(n_47),
.B1(n_49),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_0),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_0),
.A2(n_63),
.B1(n_64),
.B2(n_142),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_142),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_0),
.A2(n_27),
.B1(n_35),
.B2(n_142),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_27),
.B1(n_35),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_1),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_114),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_1),
.A2(n_47),
.B1(n_49),
.B2(n_114),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_114),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_2),
.A2(n_49),
.B(n_59),
.C(n_128),
.D(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_46),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_2),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_2),
.A2(n_82),
.B(n_147),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_2),
.A2(n_32),
.B(n_43),
.C(n_179),
.D(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_32),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_2),
.B(n_116),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_2),
.A2(n_33),
.B(n_224),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_2),
.A2(n_27),
.B1(n_35),
.B2(n_161),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_47),
.B1(n_49),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_5),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_5),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_38),
.B1(n_47),
.B2(n_49),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_38),
.B1(n_63),
.B2(n_64),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_47),
.B1(n_49),
.B2(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_8),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_10),
.B(n_64),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_10),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_10),
.A2(n_83),
.B1(n_190),
.B2(n_207),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_27),
.B1(n_35),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_12),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_12),
.A2(n_47),
.B1(n_49),
.B2(n_92),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_92),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_92),
.Y(n_181)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_16),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_16),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_16),
.A2(n_36),
.B1(n_47),
.B2(n_49),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_94),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_70),
.B2(n_71),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_26),
.A2(n_113),
.B(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_26),
.A2(n_31),
.B1(n_113),
.B2(n_250),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_27),
.A2(n_29),
.B(n_161),
.C(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_29),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_31),
.A2(n_34),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_31),
.A2(n_90),
.B(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_44),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_56),
.B1(n_57),
.B2(n_69),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_42),
.A2(n_53),
.B1(n_201),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_42),
.A2(n_238),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_46),
.B1(n_51),
.B2(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_43),
.A2(n_46),
.B1(n_73),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_43),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_44),
.B(n_49),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_45),
.A2(n_47),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_53),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_53),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_53),
.A2(n_202),
.B(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_66),
.B(n_67),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_66),
.B1(n_76),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_58),
.A2(n_66),
.B1(n_87),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_58),
.A2(n_66),
.B1(n_141),
.B2(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_58),
.A2(n_177),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_58),
.A2(n_66),
.B1(n_108),
.B2(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_62),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_59),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_60),
.B(n_64),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_61),
.A2(n_63),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_64),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_66),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_66),
.A2(n_141),
.B(n_143),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_66),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_66),
.A2(n_143),
.B(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_72),
.B(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_88),
.B(n_89),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_80),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_88),
.B1(n_89),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_81),
.A2(n_86),
.B1(n_88),
.B2(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_85),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_82),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_82),
.A2(n_106),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_82),
.A2(n_105),
.B1(n_106),
.B2(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_83),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_83),
.B(n_148),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_84),
.A2(n_153),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_84),
.B(n_161),
.Y(n_167)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_86),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_93),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_95),
.Y(n_290)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_101),
.A2(n_102),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.C(n_111),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_103),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_104),
.B(n_107),
.Y(n_263)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_109),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_110),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI321xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_278),
.A3(n_291),
.B1(n_297),
.B2(n_302),
.C(n_304),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_244),
.C(n_274),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_216),
.B(n_243),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_195),
.B(n_215),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_171),
.B(n_194),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_149),
.B(n_170),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_135),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_128),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_129),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_140),
.C(n_145),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_158),
.B(n_169),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_156),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_164),
.B(n_168),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_173),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_184),
.B2(n_193),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_183),
.C(n_193),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_180),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_188),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_209),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_211),
.C(n_213),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_204),
.B2(n_208),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_205),
.C(n_206),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_204),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_218),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_232),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_231),
.C(n_232),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_226),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_260),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_260),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_256),
.C(n_259),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_259),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_272),
.B2(n_273),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_264),
.C(n_273),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_269),
.C(n_271),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_267),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.C(n_286),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_280),
.A2(n_281),
.B1(n_284),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);


endmodule