module fake_jpeg_15098_n_24 (n_3, n_2, n_1, n_0, n_4, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_0),
.A2(n_3),
.B1(n_5),
.B2(n_2),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_8),
.B(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_14),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_7),
.A2(n_0),
.B(n_1),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_13),
.C(n_3),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_1),
.C(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_9),
.B(n_10),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_21),
.B(n_18),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_9),
.B1(n_10),
.B2(n_16),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_22),
.B(n_21),
.Y(n_24)
);


endmodule