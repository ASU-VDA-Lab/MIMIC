module fake_netlist_6_3244_n_70 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_70);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_70;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_18;
wire n_24;
wire n_21;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_48;
wire n_47;
wire n_62;
wire n_29;
wire n_65;
wire n_31;
wire n_19;
wire n_40;
wire n_57;
wire n_25;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp67_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_13),
.B(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_4),
.B(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_3),
.B(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_27),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_26),
.B(n_20),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_28),
.B(n_26),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

OAI21x1_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_28),
.B(n_31),
.Y(n_40)
);

OAI21x1_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_28),
.B(n_31),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_18),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_31),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_38),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_46),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_48),
.B(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_49),
.Y(n_58)
);

OAI322xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_25),
.A3(n_24),
.B1(n_21),
.B2(n_23),
.C1(n_51),
.C2(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_56),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_61),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_59),
.C(n_25),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_23),
.Y(n_66)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_24),
.B1(n_19),
.B2(n_17),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_24),
.B1(n_19),
.B2(n_23),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_66),
.B1(n_23),
.B2(n_19),
.Y(n_69)
);

OR2x6_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_19),
.Y(n_70)
);


endmodule