module fake_jpeg_20709_n_112 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_112);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_20),
.C(n_23),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_30),
.B1(n_22),
.B2(n_19),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_18),
.B(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_23),
.B1(n_27),
.B2(n_11),
.Y(n_41)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_37),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_32),
.B1(n_22),
.B2(n_19),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_36),
.B1(n_22),
.B2(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_34),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.C(n_35),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_10),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_16),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_59),
.B1(n_43),
.B2(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_26),
.B1(n_21),
.B2(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_51),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_48),
.B1(n_11),
.B2(n_14),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_70),
.B1(n_72),
.B2(n_13),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_45),
.C(n_46),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_63),
.C(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_58),
.B1(n_59),
.B2(n_11),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_44),
.B(n_49),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_9),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_17),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.C(n_83),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_63),
.B1(n_17),
.B2(n_14),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_14),
.B1(n_20),
.B2(n_17),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_28),
.C(n_10),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_67),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g82 ( 
.A(n_69),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_28),
.C(n_9),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_68),
.C(n_71),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_75),
.B(n_68),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_82),
.B1(n_12),
.B2(n_7),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.C(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_8),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_85),
.B1(n_90),
.B2(n_15),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_90),
.C(n_8),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_102),
.B(n_5),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_5),
.A3(n_8),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_100),
.C2(n_101),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_1),
.C(n_4),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_103),
.C(n_108),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_107),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);


endmodule