module fake_netlist_6_3526_n_108 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_108);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_108;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_28),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_30),
.B1(n_31),
.B2(n_26),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_30),
.B1(n_31),
.B2(n_26),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_43),
.Y(n_54)
);

AOI21x1_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_38),
.B(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_41),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_41),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_46),
.Y(n_60)
);

NAND2x1_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_49),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_52),
.B1(n_50),
.B2(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_45),
.Y(n_65)
);

OAI21x1_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_22),
.B(n_21),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_52),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

AO21x2_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_66),
.B(n_63),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_62),
.B(n_45),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_68),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_22),
.B1(n_35),
.B2(n_33),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_33),
.B1(n_35),
.B2(n_53),
.Y(n_85)
);

AOI211x1_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_73),
.B(n_2),
.C(n_3),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_71),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_83),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

OAI211xp5_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_83),
.B(n_93),
.C(n_92),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_52),
.B1(n_50),
.B2(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_72),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_1),
.Y(n_103)
);

AOI22x1_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_100),
.B1(n_50),
.B2(n_3),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_100),
.B1(n_2),
.B2(n_5),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_1),
.B(n_6),
.C(n_8),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_104),
.B1(n_53),
.B2(n_71),
.Y(n_107)
);

OR5x1_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_9),
.C(n_11),
.D(n_13),
.E(n_17),
.Y(n_108)
);


endmodule