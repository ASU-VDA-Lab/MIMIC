module fake_jpeg_24140_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_15),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_24),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_38),
.B1(n_37),
.B2(n_30),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_23),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_38),
.B1(n_18),
.B2(n_37),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_47),
.B1(n_52),
.B2(n_45),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_30),
.B1(n_36),
.B2(n_39),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_14),
.B(n_25),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_17),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_26),
.B(n_23),
.C(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_39),
.Y(n_89)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_27),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_0),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_0),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_79),
.B(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_76),
.B1(n_81),
.B2(n_83),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_45),
.B1(n_17),
.B2(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_82),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_35),
.B1(n_39),
.B2(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_53),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_14),
.B1(n_25),
.B2(n_27),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_68),
.B(n_57),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_20),
.B(n_26),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_100),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_26),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_63),
.B1(n_60),
.B2(n_35),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_107),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_60),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_79),
.B(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_118),
.B1(n_102),
.B2(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_64),
.C(n_70),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_113),
.C(n_117),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_64),
.C(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_62),
.B1(n_28),
.B2(n_19),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_102),
.B1(n_104),
.B2(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_73),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_62),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_62),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_55),
.C(n_77),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_96),
.C(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_134),
.B1(n_130),
.B2(n_124),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_127),
.C(n_128),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_96),
.C(n_93),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_100),
.C(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_109),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_106),
.C(n_104),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_119),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_13),
.A3(n_12),
.B1(n_11),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_118),
.B(n_110),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_137),
.B(n_143),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_108),
.B(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_35),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_1),
.Y(n_146)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_1),
.B(n_2),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_2),
.CI(n_3),
.CON(n_150),
.SN(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_13),
.B1(n_12),
.B2(n_5),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_3),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_8),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_142),
.B1(n_136),
.B2(n_7),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_158),
.B1(n_149),
.B2(n_146),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_136),
.B(n_6),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_156),
.C(n_150),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_3),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_10),
.B1(n_154),
.B2(n_109),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_147),
.C(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_161),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_150),
.C(n_9),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_168),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_165),
.Y(n_170)
);


endmodule