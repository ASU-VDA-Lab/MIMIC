module fake_jpeg_16414_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_3),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_22),
.Y(n_25)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_11),
.A2(n_8),
.B1(n_15),
.B2(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_17),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_21),
.B1(n_18),
.B2(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_36),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_0),
.B(n_3),
.Y(n_46)
);

A2O1A1O1Ixp25_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_24),
.B(n_27),
.C(n_26),
.D(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_29),
.B1(n_27),
.B2(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_15),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_42),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_6),
.A3(n_10),
.B1(n_20),
.B2(n_27),
.C1(n_29),
.C2(n_48),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);


endmodule