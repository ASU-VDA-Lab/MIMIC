module fake_jpeg_28243_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_25),
.B1(n_23),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_25),
.B1(n_22),
.B2(n_15),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_62),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_66),
.B1(n_72),
.B2(n_42),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_38),
.B1(n_35),
.B2(n_20),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_70),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_39),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_78),
.B(n_26),
.Y(n_105)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_39),
.CI(n_36),
.CON(n_70),
.SN(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_15),
.B(n_22),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_18),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_29),
.C(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_36),
.B(n_39),
.C(n_56),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_111),
.B(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_42),
.B1(n_52),
.B2(n_46),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_89),
.B1(n_101),
.B2(n_60),
.Y(n_119)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_88),
.A2(n_98),
.B1(n_104),
.B2(n_99),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_53),
.B1(n_56),
.B2(n_30),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_53),
.B1(n_15),
.B2(n_22),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_102),
.B1(n_78),
.B2(n_16),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_16),
.B1(n_28),
.B2(n_21),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_105),
.B1(n_21),
.B2(n_61),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_83),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_21),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_21),
.B(n_29),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_109),
.A2(n_69),
.B1(n_80),
.B2(n_77),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_114),
.B(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_72),
.B1(n_74),
.B2(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_120),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_119),
.B(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_78),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_68),
.B1(n_74),
.B2(n_79),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_119),
.B1(n_134),
.B2(n_140),
.Y(n_150)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_128),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_129),
.B1(n_132),
.B2(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_62),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_85),
.A2(n_88),
.B1(n_92),
.B2(n_111),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_90),
.B1(n_108),
.B2(n_102),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_81),
.C(n_17),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_101),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_89),
.B1(n_110),
.B2(n_99),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_151),
.B1(n_164),
.B2(n_17),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_166),
.B1(n_7),
.B2(n_3),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_110),
.B1(n_84),
.B2(n_91),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_84),
.B1(n_91),
.B2(n_103),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_154),
.B(n_123),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_103),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_165),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_94),
.B1(n_21),
.B2(n_19),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_94),
.B1(n_21),
.B2(n_17),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_0),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_0),
.Y(n_179)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_19),
.A3(n_17),
.B1(n_9),
.B2(n_14),
.C1(n_13),
.C2(n_11),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_8),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_123),
.B1(n_121),
.B2(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_182),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_179),
.B(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_135),
.C(n_94),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_180),
.C(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_17),
.C(n_19),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_159),
.Y(n_181)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_14),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_11),
.C(n_10),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_0),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_142),
.C(n_147),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_192),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_9),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_9),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_149),
.B(n_8),
.Y(n_194)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_1),
.B(n_3),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_170),
.B1(n_160),
.B2(n_161),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_1),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_170),
.B(n_141),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_223),
.B(n_179),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_141),
.B1(n_166),
.B2(n_145),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_149),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_145),
.B(n_167),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_175),
.A2(n_171),
.B1(n_156),
.B2(n_165),
.Y(n_225)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_178),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_211),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_212),
.B(n_201),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_176),
.C(n_191),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_235),
.C(n_240),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_198),
.B(n_199),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_222),
.B(n_216),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_177),
.C(n_183),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_180),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_202),
.C(n_193),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_187),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_245),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_217),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_202),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_248),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_255),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_258),
.B(n_213),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_207),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_210),
.B1(n_209),
.B2(n_225),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_184),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_260),
.B(n_246),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_212),
.B1(n_210),
.B2(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_241),
.B1(n_224),
.B2(n_239),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g263 ( 
.A(n_261),
.B(n_235),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_271),
.B(n_273),
.Y(n_280)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_231),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_269),
.Y(n_285)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_228),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_270),
.A2(n_257),
.B1(n_218),
.B2(n_205),
.Y(n_286)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_219),
.B1(n_224),
.B2(n_227),
.C(n_205),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_275),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_240),
.B(n_219),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_242),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_250),
.C(n_249),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_267),
.C(n_269),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_220),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_287),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_214),
.B(n_258),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_214),
.B(n_266),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_266),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_282),
.B1(n_278),
.B2(n_248),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_220),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_291),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_207),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_292),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_294),
.B(n_295),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_188),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_280),
.B1(n_253),
.B2(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_253),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_293),
.B(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_285),
.B(n_152),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_301),
.B(n_298),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_152),
.B(n_182),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_3),
.Y(n_303)
);

A2O1A1O1Ixp25_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_305),
.B(n_297),
.C(n_5),
.D(n_7),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_304),
.B(n_4),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_4),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_7),
.C(n_253),
.Y(n_311)
);


endmodule