module fake_jpeg_341_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_12),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_51),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_48),
.B1(n_51),
.B2(n_42),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_48),
.B1(n_59),
.B2(n_39),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_40),
.B1(n_46),
.B2(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_84),
.Y(n_87)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_76),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_79),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_43),
.C(n_48),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_80),
.C(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_53),
.Y(n_79)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_57),
.B1(n_39),
.B2(n_20),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_89),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_5),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_90),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_2),
.B(n_3),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_99),
.B(n_93),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_92),
.B1(n_89),
.B2(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_110),
.B1(n_112),
.B2(n_7),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_113),
.C(n_110),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_22),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_9),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_35),
.B(n_23),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_130),
.B(n_25),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_9),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_24),
.B(n_32),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_10),
.B(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_117),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_21),
.C(n_13),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_135),
.C(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_137),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_27),
.C(n_14),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_122),
.B1(n_139),
.B2(n_121),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_136),
.B(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_127),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_129),
.B1(n_142),
.B2(n_134),
.Y(n_148)
);

OAI311xp33_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_17),
.A3(n_29),
.B1(n_30),
.C1(n_31),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_129),
.B(n_34),
.Y(n_150)
);


endmodule