module fake_jpeg_5530_n_196 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_196);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_29),
.Y(n_52)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_58),
.B1(n_75),
.B2(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_24),
.B1(n_28),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_49),
.A2(n_53),
.B1(n_67),
.B2(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_52),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_27),
.B1(n_19),
.B2(n_16),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_27),
.B1(n_19),
.B2(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_14),
.B1(n_15),
.B2(n_28),
.Y(n_69)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_35),
.B(n_14),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_82),
.Y(n_84)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_37),
.A2(n_22),
.B1(n_28),
.B2(n_4),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_11),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_105),
.B1(n_106),
.B2(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_54),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_3),
.C(n_5),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_99),
.B(n_96),
.C(n_105),
.D(n_87),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_102),
.B(n_91),
.C(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_74),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_7),
.B(n_9),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_74),
.B(n_81),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_7),
.B1(n_10),
.B2(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_47),
.B1(n_76),
.B2(n_70),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_118),
.B1(n_127),
.B2(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_53),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_116),
.Y(n_151)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_123),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_81),
.B(n_48),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_64),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_59),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_84),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_65),
.B1(n_72),
.B2(n_90),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_92),
.B1(n_100),
.B2(n_85),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_108),
.C(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_139),
.Y(n_162)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_108),
.C(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_144),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_104),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_150),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_112),
.C(n_114),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_156),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_135),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_165),
.C(n_140),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_126),
.B(n_111),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_160),
.B(n_149),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_121),
.B(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_113),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_163),
.B(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_139),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_157),
.A2(n_150),
.B1(n_135),
.B2(n_133),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_176),
.B1(n_164),
.B2(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_155),
.C(n_166),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_150),
.B1(n_127),
.B2(n_130),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_180),
.A2(n_174),
.B1(n_172),
.B2(n_177),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_161),
.B(n_166),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_171),
.B(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_187),
.A2(n_180),
.B1(n_182),
.B2(n_181),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_187),
.B(n_182),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_190),
.B(n_109),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_191),
.B(n_189),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_188),
.C(n_169),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_185),
.Y(n_196)
);


endmodule