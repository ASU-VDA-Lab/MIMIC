module fake_netlist_6_661_n_1868 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1868);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1868;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_792;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1805;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_326),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_493),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_221),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_318),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_44),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_4),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_0),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_22),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_212),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_33),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_451),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_495),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_195),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_87),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_376),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_469),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_319),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_259),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_54),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_296),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_307),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_461),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_194),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_381),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_482),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_261),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_281),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_36),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_84),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_246),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_489),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_15),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_449),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_499),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_418),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_290),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_385),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_176),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_257),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_435),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_370),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_321),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_111),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_400),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_353),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_464),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_405),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_124),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_335),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_397),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_308),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_207),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_209),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_116),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_344),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_439),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_456),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_325),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_434),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g564 ( 
.A(n_234),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_336),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_172),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_96),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_309),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_317),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_229),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_128),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_46),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_425),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_351),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_190),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_24),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_19),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_306),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_21),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_275),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_80),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_82),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_109),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_328),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_458),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_199),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_260),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_297),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_231),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_192),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_448),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_178),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_382),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_189),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_250),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_205),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_267),
.Y(n_598)
);

BUFx2_ASAP7_75t_SL g599 ( 
.A(n_92),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_41),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_60),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_39),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_220),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_411),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_394),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_32),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_161),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_311),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_274),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_60),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_348),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_18),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_76),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_484),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_94),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_211),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_338),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_230),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_466),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_310),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_280),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_475),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_453),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_144),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_480),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_471),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_371),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_300),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_81),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_258),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_9),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_227),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_83),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_286),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_369),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_299),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_440),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_2),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_43),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_223),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_406),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_119),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_28),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_270),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_82),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_58),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_17),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_65),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_305),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_155),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_146),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_249),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_180),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_410),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_95),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_191),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_412),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_17),
.Y(n_658)
);

BUFx5_ASAP7_75t_L g659 ( 
.A(n_302),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_375),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_152),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_462),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_483),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_383),
.Y(n_664)
);

BUFx5_ASAP7_75t_L g665 ( 
.A(n_153),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_188),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_151),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_95),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_173),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_481),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_183),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_77),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_43),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_320),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_122),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_105),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_175),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_284),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_166),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_143),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_20),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_174),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_277),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_295),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_428),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_264),
.Y(n_686)
);

INVxp67_ASAP7_75t_SL g687 ( 
.A(n_301),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_19),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_163),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_157),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_392),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_426),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_215),
.Y(n_693)
);

BUFx10_ASAP7_75t_L g694 ( 
.A(n_387),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_98),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_49),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_479),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_85),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_30),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_437),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_433),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_10),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_255),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_145),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_206),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_331),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_143),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_333),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_219),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_151),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_22),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_73),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_498),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_494),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_665),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_638),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_665),
.Y(n_717)
);

CKINVDCx14_ASAP7_75t_R g718 ( 
.A(n_541),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_505),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_708),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_612),
.B(n_0),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_569),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_555),
.Y(n_723)
);

INVxp33_ASAP7_75t_L g724 ( 
.A(n_510),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_615),
.Y(n_725)
);

CKINVDCx16_ASAP7_75t_R g726 ( 
.A(n_507),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_535),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_508),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_665),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_506),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_512),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_665),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_535),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_665),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_665),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_665),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_513),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_515),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_516),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_519),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_555),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_520),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_521),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_581),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_523),
.Y(n_745)
);

BUFx6f_ASAP7_75t_SL g746 ( 
.A(n_664),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_564),
.B(n_1),
.Y(n_747)
);

NOR2xp67_ASAP7_75t_L g748 ( 
.A(n_642),
.B(n_1),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_513),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_509),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_582),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_582),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_629),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_524),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_629),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_647),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_564),
.B(n_2),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_531),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_527),
.Y(n_759)
);

INVxp33_ASAP7_75t_L g760 ( 
.A(n_517),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_528),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_529),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_531),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_642),
.B(n_3),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_607),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_511),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_607),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_706),
.B(n_3),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_581),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_581),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_581),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_522),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_566),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_647),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_659),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_577),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_532),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_624),
.B(n_4),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_659),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_676),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_546),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_530),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_648),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_571),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_655),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_533),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_671),
.B(n_5),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_667),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_659),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_534),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_537),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_672),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_549),
.B(n_5),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_690),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_549),
.B(n_6),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_698),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_552),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_676),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_702),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_538),
.Y(n_801)
);

CKINVDCx16_ASAP7_75t_R g802 ( 
.A(n_507),
.Y(n_802)
);

BUFx8_ASAP7_75t_L g803 ( 
.A(n_746),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_728),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_744),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_744),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_716),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_736),
.Y(n_808)
);

BUFx8_ASAP7_75t_L g809 ( 
.A(n_746),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_736),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_750),
.Y(n_811)
);

XNOR2xp5_ASAP7_75t_L g812 ( 
.A(n_727),
.B(n_548),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_723),
.B(n_671),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_728),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_719),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_715),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_730),
.B(n_568),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_744),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_717),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_769),
.B(n_568),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_729),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_731),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_741),
.B(n_675),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_732),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_734),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_738),
.B(n_623),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_735),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_770),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_775),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_771),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_739),
.B(n_623),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_740),
.B(n_575),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_741),
.B(n_575),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_766),
.B(n_558),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_749),
.B(n_675),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_775),
.B(n_580),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_747),
.A2(n_578),
.B1(n_628),
.B2(n_548),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_779),
.B(n_580),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_772),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_773),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_776),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_757),
.B(n_599),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_779),
.Y(n_843)
);

XNOR2xp5_ASAP7_75t_L g844 ( 
.A(n_727),
.B(n_578),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_790),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_758),
.B(n_664),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_763),
.B(n_664),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_790),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_781),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_748),
.B(n_595),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_766),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_765),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_784),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_786),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_789),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_793),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_742),
.B(n_595),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_777),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_743),
.B(n_598),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_721),
.A2(n_621),
.B(n_598),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_795),
.Y(n_861)
);

AND3x1_ASAP7_75t_L g862 ( 
.A(n_768),
.B(n_796),
.C(n_794),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_797),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_829),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_832),
.B(n_777),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_857),
.B(n_745),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_819),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_808),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_811),
.B(n_798),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_813),
.B(n_514),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_829),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_859),
.B(n_754),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_808),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_817),
.B(n_782),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_815),
.B(n_628),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_860),
.A2(n_504),
.B(n_503),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_862),
.A2(n_720),
.B1(n_718),
.B2(n_722),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_819),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_808),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_836),
.B(n_838),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_826),
.B(n_759),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_829),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_831),
.B(n_761),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_807),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_824),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_836),
.B(n_621),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_829),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_824),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_829),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_829),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_814),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_852),
.B(n_782),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_852),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_813),
.B(n_762),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_810),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_820),
.B(n_783),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_812),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_820),
.B(n_787),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_850),
.A2(n_778),
.B1(n_788),
.B2(n_764),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_843),
.Y(n_900)
);

OR2x6_ASAP7_75t_L g901 ( 
.A(n_842),
.B(n_725),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_852),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_839),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_810),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_820),
.B(n_791),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_820),
.B(n_800),
.Y(n_906)
);

OAI22xp33_ASAP7_75t_SL g907 ( 
.A1(n_842),
.A2(n_707),
.B1(n_712),
.B2(n_711),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_839),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_836),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_850),
.A2(n_606),
.B1(n_525),
.B2(n_536),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_837),
.B(n_785),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_846),
.B(n_792),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_840),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_836),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_840),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_816),
.B(n_801),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_846),
.B(n_746),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_810),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_823),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_822),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_843),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_843),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_L g923 ( 
.A(n_837),
.B(n_802),
.C(n_726),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_843),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_816),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_816),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_841),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_821),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_841),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_804),
.B(n_737),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_849),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_821),
.B(n_518),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_849),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_853),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_847),
.B(n_724),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_853),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_847),
.B(n_760),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_821),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_825),
.B(n_827),
.Y(n_939)
);

AND2x6_ASAP7_75t_L g940 ( 
.A(n_838),
.B(n_657),
.Y(n_940)
);

OAI22xp33_ASAP7_75t_L g941 ( 
.A1(n_842),
.A2(n_646),
.B1(n_567),
.B2(n_576),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_825),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_856),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_842),
.B(n_767),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_825),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_804),
.B(n_615),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_930),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_899),
.B(n_827),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_865),
.B(n_851),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_869),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_903),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_L g952 ( 
.A(n_881),
.B(n_659),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_900),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_900),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_899),
.B(n_827),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_914),
.B(n_860),
.Y(n_956)
);

XOR2xp5_ASAP7_75t_L g957 ( 
.A(n_911),
.B(n_812),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_897),
.B(n_851),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_914),
.B(n_838),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_919),
.A2(n_834),
.B(n_842),
.C(n_823),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_935),
.B(n_858),
.Y(n_961)
);

BUFx8_ASAP7_75t_L g962 ( 
.A(n_891),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_908),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_910),
.A2(n_838),
.B1(n_850),
.B2(n_833),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_865),
.A2(n_858),
.B1(n_714),
.B2(n_554),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_914),
.B(n_845),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_935),
.B(n_835),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_912),
.B(n_803),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_900),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_874),
.B(n_803),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_913),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_874),
.B(n_833),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_905),
.A2(n_894),
.B1(n_937),
.B2(n_892),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_937),
.B(n_803),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_884),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_866),
.B(n_833),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_946),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_870),
.B(n_803),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_872),
.B(n_833),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_870),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_910),
.A2(n_855),
.B(n_850),
.C(n_539),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_921),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_883),
.B(n_916),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_915),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_905),
.A2(n_685),
.B1(n_687),
.B2(n_550),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_867),
.B(n_845),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_892),
.B(n_809),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_878),
.B(n_845),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_875),
.Y(n_989)
);

INVxp33_ASAP7_75t_L g990 ( 
.A(n_923),
.Y(n_990)
);

BUFx5_ASAP7_75t_L g991 ( 
.A(n_940),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_896),
.B(n_844),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_893),
.B(n_855),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_898),
.B(n_844),
.Y(n_994)
);

O2A1O1Ixp5_ASAP7_75t_L g995 ( 
.A1(n_880),
.A2(n_855),
.B(n_540),
.C(n_542),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_L g996 ( 
.A(n_877),
.B(n_855),
.C(n_856),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_941),
.B(n_733),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_921),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_907),
.B(n_809),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_927),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_921),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_906),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_917),
.B(n_809),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_929),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_917),
.B(n_809),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_906),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_902),
.B(n_845),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_920),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_920),
.B(n_835),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_920),
.B(n_854),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_931),
.Y(n_1011)
);

OAI221xp5_ASAP7_75t_L g1012 ( 
.A1(n_933),
.A2(n_544),
.B1(n_637),
.B2(n_630),
.C(n_556),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_906),
.A2(n_944),
.B1(n_880),
.B2(n_901),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_885),
.B(n_848),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_944),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_922),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_934),
.B(n_854),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_936),
.A2(n_543),
.B(n_545),
.C(n_526),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_943),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_901),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_932),
.B(n_922),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_922),
.B(n_848),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_909),
.B(n_685),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_888),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_909),
.B(n_547),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_886),
.B(n_666),
.C(n_579),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_924),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_939),
.B(n_848),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_924),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_901),
.B(n_854),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_909),
.B(n_551),
.Y(n_1031)
);

NOR2xp67_ASAP7_75t_L g1032 ( 
.A(n_924),
.B(n_828),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_882),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_925),
.B(n_848),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_925),
.B(n_805),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_926),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_926),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_928),
.B(n_828),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_944),
.B(n_861),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_909),
.B(n_557),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_928),
.B(n_805),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_938),
.B(n_806),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_938),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_945),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_942),
.B(n_945),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_864),
.B(n_806),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_868),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_873),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_942),
.B(n_818),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_886),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_864),
.B(n_818),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_876),
.B(n_861),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_882),
.B(n_559),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_873),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_882),
.B(n_560),
.Y(n_1055)
);

OR2x6_ASAP7_75t_SL g1056 ( 
.A(n_879),
.B(n_572),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_L g1057 ( 
.A(n_879),
.B(n_593),
.C(n_583),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_864),
.B(n_733),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_882),
.B(n_561),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_871),
.B(n_553),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_895),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_895),
.A2(n_863),
.B(n_861),
.C(n_563),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_871),
.B(n_751),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_889),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_904),
.B(n_863),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_876),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_904),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_918),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_918),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_940),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_871),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_890),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_890),
.B(n_751),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_890),
.B(n_601),
.C(n_600),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_940),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_889),
.B(n_562),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_889),
.B(n_573),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_983),
.A2(n_570),
.B(n_574),
.C(n_565),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_1006),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_972),
.B(n_889),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_956),
.A2(n_830),
.B(n_589),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_959),
.A2(n_887),
.B(n_590),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_956),
.A2(n_863),
.B(n_830),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_973),
.B(n_1006),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_959),
.A2(n_887),
.B(n_592),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_948),
.A2(n_940),
.B1(n_604),
.B2(n_620),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_950),
.B(n_752),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_967),
.B(n_887),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1052),
.A2(n_940),
.B(n_622),
.Y(n_1089)
);

INVx11_ASAP7_75t_L g1090 ( 
.A(n_962),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_982),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1002),
.B(n_587),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_966),
.A2(n_632),
.B(n_625),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_976),
.B(n_636),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_979),
.B(n_649),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_966),
.A2(n_662),
.B(n_654),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_1006),
.B(n_584),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1050),
.A2(n_985),
.B1(n_955),
.B2(n_948),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1017),
.B(n_663),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_951),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_963),
.B(n_670),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_971),
.B(n_674),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_955),
.A2(n_683),
.B(n_684),
.C(n_678),
.Y(n_1103)
);

AND2x2_ASAP7_75t_SL g1104 ( 
.A(n_997),
.B(n_752),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1021),
.A2(n_693),
.B(n_686),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_984),
.B(n_700),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1028),
.A2(n_701),
.B(n_657),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1028),
.A2(n_657),
.B(n_586),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_993),
.A2(n_657),
.B(n_588),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_950),
.B(n_753),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_982),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_947),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_949),
.B(n_753),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1045),
.A2(n_1007),
.B(n_1022),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1013),
.A2(n_756),
.B1(n_774),
.B2(n_755),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1045),
.A2(n_964),
.B(n_1033),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1000),
.B(n_585),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1033),
.A2(n_594),
.B(n_591),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1004),
.B(n_596),
.Y(n_1119)
);

OAI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_1019),
.A2(n_610),
.B(n_602),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1033),
.A2(n_603),
.B(n_597),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_981),
.A2(n_756),
.B(n_774),
.C(n_755),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_961),
.B(n_605),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1029),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1064),
.A2(n_609),
.B(n_608),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_965),
.B(n_780),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1009),
.B(n_799),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_958),
.B(n_780),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1065),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1064),
.A2(n_1051),
.B(n_1046),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1011),
.B(n_611),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1010),
.B(n_614),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1064),
.A2(n_617),
.B(n_616),
.Y(n_1133)
);

AOI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_992),
.A2(n_799),
.B(n_631),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1029),
.A2(n_619),
.B(n_618),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_977),
.B(n_626),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_996),
.B(n_627),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1024),
.B(n_634),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1066),
.A2(n_640),
.B(n_635),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_975),
.B(n_989),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1039),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_994),
.B(n_990),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1039),
.B(n_641),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1065),
.Y(n_1144)
);

INVx4_ASAP7_75t_L g1145 ( 
.A(n_1008),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_953),
.A2(n_652),
.B(n_644),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_980),
.B(n_613),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_954),
.A2(n_998),
.B(n_969),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1030),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1036),
.B(n_656),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1035),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1035),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1037),
.B(n_660),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1058),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1001),
.A2(n_692),
.B(n_691),
.Y(n_1155)
);

AO21x1_ASAP7_75t_L g1156 ( 
.A1(n_952),
.A2(n_659),
.B(n_694),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1026),
.B(n_1074),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1012),
.A2(n_697),
.B(n_705),
.C(n_703),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1016),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1043),
.B(n_1044),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1032),
.A2(n_659),
.B(n_709),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1070),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1027),
.A2(n_713),
.B(n_643),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1054),
.B(n_659),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_1075),
.B(n_694),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_L g1166 ( 
.A(n_1057),
.B(n_645),
.C(n_633),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1034),
.A2(n_651),
.B(n_650),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1061),
.B(n_653),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1034),
.A2(n_661),
.B(n_658),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_987),
.B(n_186),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_986),
.A2(n_669),
.B(n_668),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_986),
.A2(n_679),
.B(n_677),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1063),
.B(n_680),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_988),
.A2(n_682),
.B(n_681),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1020),
.B(n_694),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1047),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_1072),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_995),
.A2(n_689),
.B(n_695),
.C(n_688),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1071),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1067),
.B(n_1068),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1069),
.B(n_696),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_988),
.A2(n_1014),
.B(n_1041),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1060),
.A2(n_193),
.B(n_187),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_957),
.B(n_699),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1014),
.A2(n_710),
.B(n_704),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1048),
.B(n_6),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1041),
.A2(n_197),
.B(n_196),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1042),
.B(n_7),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1042),
.B(n_7),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1049),
.A2(n_200),
.B(n_198),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1023),
.A2(n_202),
.B1(n_203),
.B2(n_201),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1049),
.B(n_1038),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1053),
.A2(n_208),
.B(n_204),
.Y(n_1193)
);

OAI321xp33_ASAP7_75t_L g1194 ( 
.A1(n_1073),
.A2(n_673),
.A3(n_615),
.B1(n_10),
.B2(n_12),
.C(n_8),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1055),
.A2(n_213),
.B(n_210),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_991),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_978),
.B(n_673),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1015),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1062),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1059),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_970),
.A2(n_673),
.B(n_11),
.C(n_8),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_962),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_999),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1076),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_974),
.B(n_9),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1077),
.B(n_11),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1025),
.B(n_12),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_991),
.B(n_214),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1025),
.B(n_13),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_991),
.B(n_13),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_991),
.B(n_216),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1056),
.B(n_14),
.Y(n_1212)
);

AOI222xp33_ASAP7_75t_L g1213 ( 
.A1(n_968),
.A2(n_16),
.B1(n_20),
.B2(n_14),
.C1(n_15),
.C2(n_18),
.Y(n_1213)
);

CKINVDCx10_ASAP7_75t_R g1214 ( 
.A(n_1003),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1031),
.A2(n_218),
.B(n_217),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_1005),
.A2(n_1040),
.B(n_991),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1018),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_983),
.B(n_16),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_983),
.B(n_21),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_975),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_973),
.B(n_222),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_983),
.B(n_23),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_L g1223 ( 
.A(n_991),
.B(n_224),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_951),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_983),
.B(n_23),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_983),
.B(n_24),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_983),
.B(n_25),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_959),
.A2(n_226),
.B(n_225),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_973),
.B(n_228),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_983),
.B(n_25),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_973),
.B(n_232),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_983),
.B(n_26),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1008),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_983),
.B(n_26),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_951),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_975),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_983),
.B(n_27),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_SL g1238 ( 
.A(n_1008),
.B(n_27),
.Y(n_1238)
);

NOR3xp33_ASAP7_75t_L g1239 ( 
.A(n_992),
.B(n_28),
.C(n_29),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_950),
.B(n_29),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_956),
.A2(n_235),
.B(n_233),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_959),
.A2(n_237),
.B(n_236),
.Y(n_1242)
);

AOI21xp33_ASAP7_75t_L g1243 ( 
.A1(n_985),
.A2(n_30),
.B(n_31),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_960),
.A2(n_31),
.B(n_32),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_956),
.A2(n_239),
.B(n_238),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_983),
.B(n_33),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_959),
.A2(n_241),
.B(n_240),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_983),
.A2(n_243),
.B1(n_244),
.B2(n_242),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1006),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_973),
.A2(n_247),
.B1(n_248),
.B2(n_245),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1006),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_959),
.A2(n_252),
.B(n_251),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1006),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_973),
.A2(n_254),
.B1(n_256),
.B2(n_253),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_983),
.B(n_34),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1006),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_983),
.B(n_34),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_959),
.A2(n_263),
.B(n_262),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_983),
.B(n_35),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1079),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1225),
.A2(n_266),
.B1(n_268),
.B2(n_265),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1142),
.B(n_35),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1110),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1080),
.A2(n_271),
.B(n_269),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1141),
.B(n_272),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1151),
.B(n_36),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1089),
.A2(n_276),
.B(n_273),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1152),
.B(n_37),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1257),
.B(n_37),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1088),
.A2(n_279),
.B(n_278),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1084),
.A2(n_283),
.B1(n_285),
.B2(n_282),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1079),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1100),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1182),
.A2(n_288),
.B(n_287),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_L g1275 ( 
.A(n_1173),
.B(n_38),
.C(n_39),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1083),
.A2(n_291),
.B(n_289),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1218),
.A2(n_293),
.B1(n_294),
.B2(n_292),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1098),
.A2(n_303),
.B1(n_304),
.B2(n_298),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1127),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1219),
.A2(n_313),
.B1(n_314),
.B2(n_312),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1116),
.A2(n_316),
.B(n_315),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1087),
.B(n_38),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1141),
.B(n_322),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1176),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1192),
.A2(n_324),
.B(n_323),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1141),
.B(n_327),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1114),
.A2(n_330),
.B(n_329),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1259),
.B(n_40),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1149),
.B(n_332),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1198),
.B(n_334),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1222),
.B(n_40),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1226),
.B(n_41),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1227),
.B(n_42),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1154),
.B(n_337),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1079),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1230),
.B(n_42),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1243),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1297)
);

AOI33xp33_ASAP7_75t_L g1298 ( 
.A1(n_1212),
.A2(n_45),
.A3(n_47),
.B1(n_48),
.B2(n_49),
.B3(n_50),
.Y(n_1298)
);

O2A1O1Ixp5_ASAP7_75t_L g1299 ( 
.A1(n_1157),
.A2(n_1234),
.B(n_1237),
.C(n_1232),
.Y(n_1299)
);

NOR2x1_ASAP7_75t_L g1300 ( 
.A(n_1145),
.B(n_339),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1246),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1224),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1255),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1303)
);

NOR3xp33_ASAP7_75t_SL g1304 ( 
.A(n_1115),
.B(n_51),
.C(n_52),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1154),
.B(n_53),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1128),
.B(n_54),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1251),
.B(n_340),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1112),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1130),
.A2(n_342),
.B(n_341),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1129),
.B(n_55),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1205),
.A2(n_345),
.B1(n_346),
.B2(n_343),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1134),
.B(n_55),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1144),
.A2(n_349),
.B1(n_350),
.B2(n_347),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1094),
.A2(n_354),
.B(n_352),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1104),
.B(n_56),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1235),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1095),
.A2(n_356),
.B1(n_357),
.B2(n_355),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1221),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1318)
);

OAI21xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1241),
.A2(n_57),
.B(n_59),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1240),
.B(n_59),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1223),
.A2(n_359),
.B(n_358),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1113),
.B(n_61),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1123),
.B(n_61),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1132),
.B(n_360),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1229),
.A2(n_362),
.B(n_361),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1220),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1233),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1162),
.B(n_1251),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1126),
.B(n_62),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1231),
.A2(n_364),
.B(n_363),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1184),
.B(n_62),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1236),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1188),
.B(n_1189),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1213),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1124),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1124),
.A2(n_372),
.B1(n_373),
.B2(n_368),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1159),
.Y(n_1338)
);

O2A1O1Ixp5_ASAP7_75t_L g1339 ( 
.A1(n_1139),
.A2(n_377),
.B(n_378),
.C(n_374),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1200),
.B(n_63),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1148),
.A2(n_380),
.B(n_379),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1201),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1180),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1091),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1090),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1082),
.A2(n_386),
.B(n_384),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1179),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1162),
.A2(n_502),
.B1(n_501),
.B2(n_500),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1085),
.A2(n_389),
.B(n_388),
.Y(n_1349)
);

AOI21xp33_ASAP7_75t_L g1350 ( 
.A1(n_1122),
.A2(n_64),
.B(n_66),
.Y(n_1350)
);

OAI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1197),
.A2(n_66),
.B(n_67),
.Y(n_1351)
);

AND2x2_ASAP7_75t_SL g1352 ( 
.A(n_1238),
.B(n_67),
.Y(n_1352)
);

AND2x6_ASAP7_75t_L g1353 ( 
.A(n_1196),
.B(n_390),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1162),
.B(n_393),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_SL g1355 ( 
.A(n_1202),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1111),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1131),
.B(n_395),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1194),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1203),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1099),
.A2(n_398),
.B(n_396),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1186),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_SL g1362 ( 
.A(n_1175),
.B(n_68),
.C(n_69),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1204),
.B(n_70),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1147),
.B(n_71),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1249),
.B(n_71),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1092),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1097),
.A2(n_401),
.B(n_399),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1249),
.B(n_1253),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1179),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1253),
.B(n_402),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1092),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1179),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1245),
.A2(n_404),
.B(n_403),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1208),
.A2(n_408),
.B(n_407),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1140),
.B(n_72),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1117),
.B(n_72),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1244),
.A2(n_1217),
.B1(n_1239),
.B2(n_1206),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1101),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1145),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1177),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1078),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1256),
.B(n_409),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1238),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1211),
.A2(n_1138),
.B(n_1137),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1102),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1256),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1143),
.A2(n_414),
.B(n_413),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1170),
.A2(n_74),
.B(n_75),
.C(n_76),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1086),
.A2(n_497),
.B1(n_496),
.B2(n_492),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1177),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1158),
.A2(n_77),
.B(n_78),
.C(n_79),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1136),
.A2(n_416),
.B(n_415),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1119),
.B(n_1175),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1120),
.B(n_78),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1106),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1120),
.B(n_1168),
.Y(n_1396)
);

AOI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1161),
.A2(n_419),
.B(n_417),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1181),
.B(n_79),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1171),
.B(n_80),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1217),
.A2(n_491),
.B1(n_490),
.B2(n_488),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1150),
.A2(n_421),
.B(n_420),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1153),
.A2(n_423),
.B(n_422),
.Y(n_1402)
);

CKINVDCx14_ASAP7_75t_R g1403 ( 
.A(n_1191),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1081),
.A2(n_427),
.B(n_424),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1199),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1167),
.B(n_81),
.Y(n_1406)
);

OAI22x1_ASAP7_75t_L g1407 ( 
.A1(n_1214),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_1407)
);

O2A1O1Ixp5_ASAP7_75t_SL g1408 ( 
.A1(n_1250),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1165),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1103),
.A2(n_86),
.B(n_88),
.C(n_89),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1164),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1215),
.A2(n_487),
.B(n_486),
.Y(n_1412)
);

NOR3xp33_ASAP7_75t_L g1413 ( 
.A(n_1166),
.B(n_89),
.C(n_90),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1207),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1169),
.B(n_90),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1166),
.B(n_91),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1172),
.B(n_91),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1210),
.A2(n_485),
.B(n_478),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1209),
.Y(n_1419)
);

NOR3xp33_ASAP7_75t_L g1420 ( 
.A(n_1254),
.B(n_92),
.C(n_93),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1248),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1174),
.B(n_97),
.Y(n_1422)
);

NOR3xp33_ASAP7_75t_L g1423 ( 
.A(n_1185),
.B(n_97),
.C(n_98),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1216),
.B(n_429),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1178),
.B(n_430),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1135),
.B(n_99),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1093),
.B(n_99),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1118),
.B(n_100),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1121),
.B(n_100),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1228),
.A2(n_477),
.B(n_476),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1096),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1125),
.B(n_101),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1105),
.B(n_101),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1107),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1183),
.Y(n_1435)
);

INVx6_ASAP7_75t_L g1436 ( 
.A(n_1165),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1165),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1156),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1273),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1263),
.B(n_1108),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1302),
.Y(n_1441)
);

NOR2xp67_ASAP7_75t_L g1442 ( 
.A(n_1326),
.B(n_1419),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1364),
.A2(n_1396),
.B(n_1329),
.C(n_1299),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1341),
.A2(n_1258),
.B(n_1252),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1403),
.A2(n_1163),
.B1(n_1109),
.B2(n_1247),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1315),
.B(n_1165),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1383),
.B(n_1133),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1287),
.A2(n_1242),
.B(n_1190),
.Y(n_1448)
);

BUFx4f_ASAP7_75t_L g1449 ( 
.A(n_1295),
.Y(n_1449)
);

AOI221x1_ASAP7_75t_L g1450 ( 
.A1(n_1420),
.A2(n_1187),
.B1(n_1193),
.B2(n_1195),
.C(n_1155),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1435),
.A2(n_1146),
.A3(n_474),
.B(n_473),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1332),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1379),
.B(n_431),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1345),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1327),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1262),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1336),
.B(n_102),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1343),
.B(n_1378),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1276),
.A2(n_472),
.B(n_470),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1279),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1322),
.B(n_103),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1308),
.B(n_104),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1359),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1384),
.A2(n_468),
.B(n_467),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1333),
.A2(n_465),
.B(n_463),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1312),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_1466)
);

NOR2xp67_ASAP7_75t_L g1467 ( 
.A(n_1323),
.B(n_460),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1385),
.B(n_1395),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1334),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1281),
.A2(n_459),
.B(n_457),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1295),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1414),
.B(n_108),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1376),
.A2(n_1334),
.B(n_1373),
.C(n_1319),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_SL g1474 ( 
.A(n_1352),
.B(n_432),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1269),
.A2(n_109),
.B(n_110),
.C(n_111),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1319),
.A2(n_110),
.B(n_112),
.C(n_113),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1316),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1431),
.A2(n_454),
.B(n_452),
.Y(n_1478)
);

AO32x2_ASAP7_75t_L g1479 ( 
.A1(n_1421),
.A2(n_112),
.A3(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1295),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1412),
.A2(n_450),
.B(n_447),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1267),
.A2(n_446),
.B(n_445),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1393),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1438),
.A2(n_444),
.B(n_443),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1434),
.A2(n_441),
.B(n_438),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1290),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1282),
.B(n_1361),
.Y(n_1487)
);

AOI21xp33_ASAP7_75t_L g1488 ( 
.A1(n_1377),
.A2(n_114),
.B(n_115),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1351),
.A2(n_116),
.B(n_117),
.C(n_118),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1405),
.B(n_117),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1290),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1366),
.B(n_118),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1354),
.B(n_436),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1320),
.B(n_1371),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1354),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1266),
.B(n_185),
.Y(n_1496)
);

AOI221x1_ASAP7_75t_L g1497 ( 
.A1(n_1351),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.C(n_122),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1274),
.A2(n_123),
.B(n_124),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1268),
.B(n_1288),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1411),
.A2(n_125),
.B(n_126),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1291),
.B(n_184),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1284),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1394),
.A2(n_126),
.B(n_127),
.C(n_128),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1309),
.A2(n_127),
.B(n_129),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1321),
.A2(n_129),
.B(n_130),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1260),
.Y(n_1506)
);

AO31x2_ASAP7_75t_L g1507 ( 
.A1(n_1391),
.A2(n_1410),
.A3(n_1292),
.B(n_1293),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1397),
.A2(n_130),
.B(n_131),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1296),
.A2(n_131),
.B(n_132),
.Y(n_1509)
);

O2A1O1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1306),
.A2(n_132),
.B(n_133),
.C(n_134),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1424),
.A2(n_133),
.B(n_134),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1324),
.A2(n_135),
.B(n_136),
.Y(n_1512)
);

AOI31xp67_ASAP7_75t_L g1513 ( 
.A1(n_1278),
.A2(n_135),
.A3(n_136),
.B(n_137),
.Y(n_1513)
);

AO32x2_ASAP7_75t_L g1514 ( 
.A1(n_1271),
.A2(n_137),
.A3(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1422),
.A2(n_138),
.B(n_139),
.C(n_140),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1338),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1289),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1398),
.A2(n_141),
.B(n_142),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1390),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_1519)
);

AO31x2_ASAP7_75t_L g1520 ( 
.A1(n_1430),
.A2(n_184),
.A3(n_146),
.B(n_147),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1305),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1416),
.A2(n_145),
.B(n_147),
.C(n_148),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1331),
.B(n_148),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1418),
.A2(n_149),
.B(n_150),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1390),
.B(n_149),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1390),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1404),
.A2(n_150),
.B(n_152),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1310),
.A2(n_183),
.B(n_154),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1272),
.Y(n_1529)
);

NOR2xp67_ASAP7_75t_L g1530 ( 
.A(n_1344),
.B(n_153),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1340),
.B(n_182),
.Y(n_1531)
);

AO31x2_ASAP7_75t_L g1532 ( 
.A1(n_1388),
.A2(n_154),
.A3(n_155),
.B(n_156),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1375),
.B(n_156),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1407),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1426),
.A2(n_158),
.B(n_159),
.C(n_160),
.Y(n_1535)
);

NOR2xp67_ASAP7_75t_L g1536 ( 
.A(n_1356),
.B(n_160),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1289),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1369),
.Y(n_1538)
);

OAI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1417),
.A2(n_161),
.B(n_162),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1406),
.A2(n_182),
.B(n_163),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1437),
.A2(n_162),
.B(n_164),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1425),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1357),
.A2(n_165),
.B(n_167),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1380),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1270),
.A2(n_168),
.B(n_169),
.Y(n_1545)
);

NAND2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1260),
.B(n_170),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1318),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_1547)
);

BUFx8_ASAP7_75t_L g1548 ( 
.A(n_1355),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1363),
.B(n_1372),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1304),
.B(n_1413),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1328),
.B(n_1335),
.Y(n_1551)
);

AO32x2_ASAP7_75t_L g1552 ( 
.A1(n_1277),
.A2(n_171),
.A3(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1365),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1325),
.A2(n_1330),
.B(n_1402),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1264),
.A2(n_176),
.B(n_177),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1358),
.B(n_181),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1401),
.A2(n_1360),
.B(n_1346),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1425),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_1558)
);

AO31x2_ASAP7_75t_L g1559 ( 
.A1(n_1303),
.A2(n_179),
.A3(n_180),
.B(n_181),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1272),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_L g1561 ( 
.A(n_1347),
.B(n_1335),
.Y(n_1561)
);

CKINVDCx11_ASAP7_75t_R g1562 ( 
.A(n_1307),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1347),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1368),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1339),
.A2(n_1415),
.B(n_1427),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1349),
.A2(n_1285),
.B(n_1314),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1370),
.Y(n_1567)
);

AO31x2_ASAP7_75t_L g1568 ( 
.A1(n_1280),
.A2(n_1317),
.A3(n_1389),
.B(n_1313),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1294),
.A2(n_1428),
.B1(n_1429),
.B2(n_1432),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1298),
.B(n_1370),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1399),
.B(n_1386),
.Y(n_1571)
);

AO31x2_ASAP7_75t_L g1572 ( 
.A1(n_1400),
.A2(n_1261),
.A3(n_1433),
.B(n_1337),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1386),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1307),
.Y(n_1574)
);

AO31x2_ASAP7_75t_L g1575 ( 
.A1(n_1374),
.A2(n_1348),
.A3(n_1367),
.B(n_1387),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1300),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1382),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1392),
.A2(n_1265),
.B(n_1286),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1301),
.B(n_1350),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1342),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1362),
.A2(n_1297),
.B(n_1423),
.C(n_1381),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1408),
.A2(n_1278),
.B(n_1275),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1311),
.B(n_1283),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1353),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1353),
.B(n_1311),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1353),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1460),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1455),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1562),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1439),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1441),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1474),
.A2(n_1409),
.B1(n_1436),
.B2(n_1355),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1533),
.B(n_1353),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1526),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1527),
.A2(n_1409),
.B(n_1508),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1550),
.A2(n_1469),
.B1(n_1569),
.B2(n_1583),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1454),
.Y(n_1597)
);

BUFx8_ASAP7_75t_SL g1598 ( 
.A(n_1483),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1477),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1443),
.A2(n_1521),
.B1(n_1473),
.B2(n_1491),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1463),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1452),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1519),
.A2(n_1509),
.B1(n_1518),
.B2(n_1547),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1548),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1449),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1502),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1495),
.Y(n_1607)
);

OAI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1542),
.A2(n_1558),
.B1(n_1456),
.B2(n_1556),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1487),
.B(n_1461),
.Y(n_1609)
);

CKINVDCx11_ASAP7_75t_R g1610 ( 
.A(n_1486),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1458),
.A2(n_1585),
.B1(n_1468),
.B2(n_1570),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1564),
.Y(n_1612)
);

INVx6_ASAP7_75t_L g1613 ( 
.A(n_1526),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1534),
.A2(n_1539),
.B1(n_1540),
.B2(n_1528),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1488),
.A2(n_1579),
.B1(n_1524),
.B2(n_1580),
.Y(n_1615)
);

CKINVDCx6p67_ASAP7_75t_R g1616 ( 
.A(n_1453),
.Y(n_1616)
);

BUFx4_ASAP7_75t_R g1617 ( 
.A(n_1529),
.Y(n_1617)
);

INVx6_ASAP7_75t_L g1618 ( 
.A(n_1486),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1506),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1446),
.A2(n_1493),
.B1(n_1576),
.B2(n_1499),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1517),
.A2(n_1537),
.B1(n_1574),
.B2(n_1567),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1544),
.A2(n_1462),
.B1(n_1457),
.B2(n_1501),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1553),
.B(n_1494),
.Y(n_1623)
);

CKINVDCx6p67_ASAP7_75t_R g1624 ( 
.A(n_1453),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1516),
.Y(n_1625)
);

CKINVDCx11_ASAP7_75t_R g1626 ( 
.A(n_1493),
.Y(n_1626)
);

INVx4_ASAP7_75t_L g1627 ( 
.A(n_1577),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1471),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1549),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1582),
.A2(n_1512),
.B1(n_1543),
.B2(n_1440),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1442),
.A2(n_1531),
.B1(n_1496),
.B2(n_1571),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1538),
.Y(n_1632)
);

INVx6_ASAP7_75t_L g1633 ( 
.A(n_1577),
.Y(n_1633)
);

OAI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1497),
.A2(n_1472),
.B1(n_1484),
.B2(n_1546),
.Y(n_1634)
);

INVx6_ASAP7_75t_L g1635 ( 
.A(n_1480),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1560),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1445),
.A2(n_1505),
.B1(n_1504),
.B2(n_1498),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1584),
.A2(n_1586),
.B1(n_1551),
.B2(n_1490),
.Y(n_1638)
);

CKINVDCx6p67_ASAP7_75t_R g1639 ( 
.A(n_1525),
.Y(n_1639)
);

CKINVDCx16_ASAP7_75t_R g1640 ( 
.A(n_1573),
.Y(n_1640)
);

INVx6_ASAP7_75t_L g1641 ( 
.A(n_1561),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1545),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1511),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1541),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1513),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1500),
.A2(n_1481),
.B1(n_1482),
.B2(n_1479),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1555),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1492),
.B(n_1507),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1581),
.B(n_1467),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1563),
.Y(n_1650)
);

INVx4_ASAP7_75t_L g1651 ( 
.A(n_1565),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1489),
.B(n_1447),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1530),
.A2(n_1536),
.B1(n_1503),
.B2(n_1522),
.Y(n_1653)
);

NAND2x1p5_ASAP7_75t_L g1654 ( 
.A(n_1578),
.B(n_1470),
.Y(n_1654)
);

INVx6_ASAP7_75t_L g1655 ( 
.A(n_1510),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1565),
.A2(n_1465),
.B1(n_1478),
.B2(n_1485),
.Y(n_1656)
);

OAI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1450),
.A2(n_1479),
.B1(n_1557),
.B2(n_1554),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1451),
.Y(n_1658)
);

INVx3_ASAP7_75t_SL g1659 ( 
.A(n_1532),
.Y(n_1659)
);

INVx6_ASAP7_75t_L g1660 ( 
.A(n_1535),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1476),
.A2(n_1515),
.B1(n_1466),
.B2(n_1475),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1566),
.A2(n_1479),
.B1(n_1572),
.B2(n_1568),
.Y(n_1662)
);

INVx3_ASAP7_75t_SL g1663 ( 
.A(n_1520),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1464),
.A2(n_1444),
.B1(n_1448),
.B2(n_1459),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1514),
.A2(n_1568),
.B1(n_1552),
.B2(n_1572),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1514),
.A2(n_1552),
.B1(n_1559),
.B2(n_1575),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_SL g1667 ( 
.A1(n_1514),
.A2(n_1552),
.B1(n_1559),
.B2(n_1575),
.Y(n_1667)
);

INVx6_ASAP7_75t_L g1668 ( 
.A(n_1520),
.Y(n_1668)
);

BUFx12f_ASAP7_75t_L g1669 ( 
.A(n_1451),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1562),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1454),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1449),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1523),
.A2(n_1329),
.B1(n_1104),
.B2(n_1126),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1439),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1449),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1474),
.A2(n_875),
.B1(n_1334),
.B2(n_1175),
.Y(n_1676)
);

OAI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1474),
.A2(n_875),
.B1(n_1334),
.B2(n_1175),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1455),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1455),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1562),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1460),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1474),
.A2(n_1104),
.B1(n_1329),
.B2(n_1352),
.Y(n_1682)
);

INVx3_ASAP7_75t_SL g1683 ( 
.A(n_1460),
.Y(n_1683)
);

INVx3_ASAP7_75t_SL g1684 ( 
.A(n_1460),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1673),
.A2(n_1614),
.B(n_1649),
.Y(n_1685)
);

INVx6_ASAP7_75t_SL g1686 ( 
.A(n_1617),
.Y(n_1686)
);

AO21x2_ASAP7_75t_L g1687 ( 
.A1(n_1657),
.A2(n_1645),
.B(n_1658),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1590),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1603),
.A2(n_1622),
.B(n_1682),
.C(n_1653),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_SL g1690 ( 
.A1(n_1648),
.A2(n_1611),
.B(n_1600),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1665),
.B(n_1659),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1629),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1632),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1590),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1591),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1601),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1667),
.B(n_1666),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1609),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1651),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1588),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1591),
.Y(n_1701)
);

AO21x2_ASAP7_75t_L g1702 ( 
.A1(n_1647),
.A2(n_1644),
.B(n_1662),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1668),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1663),
.B(n_1612),
.Y(n_1704)
);

AOI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1652),
.A2(n_1642),
.B(n_1661),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1587),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1596),
.A2(n_1615),
.B1(n_1655),
.B2(n_1637),
.C(n_1630),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1668),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1664),
.A2(n_1654),
.B(n_1656),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1650),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1669),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1674),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1623),
.B(n_1631),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1620),
.B(n_1606),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1643),
.A2(n_1595),
.B(n_1638),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1660),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1599),
.Y(n_1717)
);

CKINVDCx20_ASAP7_75t_R g1718 ( 
.A(n_1598),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1640),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1635),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1625),
.B(n_1593),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1660),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1635),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1636),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1646),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1627),
.B(n_1628),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1608),
.B(n_1655),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1621),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1616),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1681),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1715),
.A2(n_1634),
.B(n_1676),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1716),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1721),
.B(n_1678),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1721),
.B(n_1594),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1712),
.B(n_1679),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1727),
.B(n_1677),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1701),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_R g1739 ( 
.A(n_1719),
.B(n_1626),
.Y(n_1739)
);

OA21x2_ASAP7_75t_L g1740 ( 
.A1(n_1715),
.A2(n_1592),
.B(n_1639),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1690),
.B(n_1627),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1689),
.A2(n_1624),
.B(n_1594),
.C(n_1675),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1709),
.A2(n_1641),
.B(n_1633),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1744)
);

NOR2x1_ASAP7_75t_L g1745 ( 
.A(n_1713),
.B(n_1619),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1726),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1685),
.A2(n_1641),
.B1(n_1607),
.B2(n_1602),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.B(n_1684),
.Y(n_1748)
);

AO32x2_ASAP7_75t_L g1749 ( 
.A1(n_1697),
.A2(n_1672),
.A3(n_1619),
.B1(n_1610),
.B2(n_1633),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_L g1750 ( 
.A(n_1716),
.B(n_1675),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1704),
.B(n_1618),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1691),
.B(n_1618),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1690),
.B(n_1675),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1698),
.B(n_1719),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1707),
.A2(n_1605),
.B(n_1604),
.C(n_1680),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1725),
.A2(n_1605),
.B(n_1589),
.C(n_1670),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1694),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1693),
.B(n_1597),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1708),
.B(n_1672),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1716),
.B(n_1605),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1725),
.A2(n_1613),
.B1(n_1671),
.B2(n_1697),
.C(n_1728),
.Y(n_1761)
);

BUFx4f_ASAP7_75t_SL g1762 ( 
.A(n_1686),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1695),
.B(n_1613),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1738),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1734),
.Y(n_1765)
);

AND2x4_ASAP7_75t_SL g1766 ( 
.A(n_1741),
.B(n_1711),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1736),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1752),
.B(n_1699),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1743),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1741),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1730),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1743),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1754),
.B(n_1696),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1717),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1757),
.B(n_1687),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1763),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1731),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1763),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_SL g1779 ( 
.A(n_1762),
.B(n_1718),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1746),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1746),
.Y(n_1781)
);

BUFx2_ASAP7_75t_L g1782 ( 
.A(n_1769),
.Y(n_1782)
);

OAI222xp33_ASAP7_75t_L g1783 ( 
.A1(n_1774),
.A2(n_1737),
.B1(n_1753),
.B2(n_1741),
.C1(n_1745),
.C2(n_1748),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1767),
.B(n_1761),
.C(n_1731),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1776),
.B(n_1744),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1768),
.B(n_1752),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1771),
.A2(n_1731),
.B1(n_1741),
.B2(n_1753),
.Y(n_1787)
);

OR2x6_ASAP7_75t_L g1788 ( 
.A(n_1770),
.B(n_1711),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1765),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1765),
.Y(n_1790)
);

INVxp67_ASAP7_75t_SL g1791 ( 
.A(n_1775),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1775),
.B(n_1687),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1778),
.A2(n_1747),
.B1(n_1716),
.B2(n_1722),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1780),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1778),
.B(n_1687),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1776),
.B(n_1702),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1780),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1773),
.A2(n_1716),
.B1(n_1722),
.B2(n_1711),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1789),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1788),
.B(n_1770),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1789),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1790),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1790),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1795),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1785),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1788),
.B(n_1770),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1805),
.B(n_1784),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1800),
.B(n_1785),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1804),
.B(n_1791),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1800),
.B(n_1797),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1799),
.Y(n_1811)
);

OAI211xp5_ASAP7_75t_L g1812 ( 
.A1(n_1807),
.A2(n_1742),
.B(n_1787),
.C(n_1755),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1808),
.B(n_1786),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1811),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1810),
.B(n_1809),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1809),
.B(n_1803),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1811),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_L g1818 ( 
.A(n_1814),
.B(n_1755),
.C(n_1742),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1815),
.B(n_1739),
.Y(n_1819)
);

OAI222xp33_ASAP7_75t_L g1820 ( 
.A1(n_1816),
.A2(n_1788),
.B1(n_1806),
.B2(n_1782),
.C1(n_1798),
.C2(n_1793),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1818),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1819),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1821),
.A2(n_1820),
.B1(n_1812),
.B2(n_1817),
.C1(n_1783),
.C2(n_1756),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1823),
.B(n_1822),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1824),
.A2(n_1756),
.B1(n_1782),
.B2(n_1700),
.C(n_1706),
.Y(n_1825)
);

NOR3xp33_ASAP7_75t_L g1826 ( 
.A(n_1824),
.B(n_1729),
.C(n_1758),
.Y(n_1826)
);

O2A1O1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1729),
.B(n_1804),
.C(n_1813),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1825),
.A2(n_1779),
.B(n_1729),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1827),
.Y(n_1829)
);

NOR2xp67_ASAP7_75t_SL g1830 ( 
.A(n_1828),
.B(n_1720),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1828),
.A2(n_1806),
.B1(n_1760),
.B2(n_1788),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1830),
.B(n_1801),
.Y(n_1832)
);

OAI21xp33_ASAP7_75t_SL g1833 ( 
.A1(n_1831),
.A2(n_1802),
.B(n_1801),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1829),
.A2(n_1720),
.B(n_1723),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1834),
.B(n_1802),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_R g1836 ( 
.A(n_1832),
.B(n_1686),
.Y(n_1836)
);

AO22x2_ASAP7_75t_L g1837 ( 
.A1(n_1833),
.A2(n_1723),
.B1(n_1806),
.B2(n_1726),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1832),
.A2(n_1760),
.B1(n_1726),
.B2(n_1750),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1832),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1832),
.Y(n_1840)
);

OA22x2_ASAP7_75t_L g1841 ( 
.A1(n_1832),
.A2(n_1726),
.B1(n_1724),
.B2(n_1766),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1839),
.A2(n_1750),
.B1(n_1751),
.B2(n_1770),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1840),
.A2(n_1797),
.B1(n_1724),
.B2(n_1716),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1837),
.A2(n_1711),
.B1(n_1794),
.B2(n_1759),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1838),
.A2(n_1686),
.B1(n_1711),
.B2(n_1772),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1835),
.A2(n_1711),
.B1(n_1759),
.B2(n_1733),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1841),
.A2(n_1759),
.B1(n_1766),
.B2(n_1769),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1836),
.A2(n_1766),
.B1(n_1772),
.B2(n_1769),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1839),
.Y(n_1849)
);

NOR4xp25_ASAP7_75t_L g1850 ( 
.A(n_1849),
.B(n_1795),
.C(n_1792),
.D(n_1686),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1842),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1845),
.A2(n_1772),
.B1(n_1732),
.B2(n_1740),
.Y(n_1852)
);

XNOR2xp5_ASAP7_75t_L g1853 ( 
.A(n_1846),
.B(n_1735),
.Y(n_1853)
);

NAND2xp33_ASAP7_75t_L g1854 ( 
.A(n_1843),
.B(n_1732),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1844),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1848),
.A2(n_1792),
.B1(n_1796),
.B2(n_1777),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1847),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1796),
.B1(n_1781),
.B2(n_1777),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1855),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1851),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_L g1861 ( 
.A(n_1859),
.B(n_1854),
.C(n_1853),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1860),
.A2(n_1850),
.B(n_1856),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1862),
.B(n_1858),
.Y(n_1863)
);

AOI21xp33_ASAP7_75t_L g1864 ( 
.A1(n_1863),
.A2(n_1861),
.B(n_1852),
.Y(n_1864)
);

AND3x4_ASAP7_75t_L g1865 ( 
.A(n_1864),
.B(n_1749),
.C(n_1777),
.Y(n_1865)
);

OAI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1864),
.A2(n_1732),
.B1(n_1714),
.B2(n_1781),
.Y(n_1866)
);

OAI221xp5_ASAP7_75t_R g1867 ( 
.A1(n_1866),
.A2(n_1749),
.B1(n_1740),
.B2(n_1732),
.C(n_1705),
.Y(n_1867)
);

AOI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1867),
.A2(n_1865),
.B(n_1703),
.C(n_1764),
.Y(n_1868)
);


endmodule