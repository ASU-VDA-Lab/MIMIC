module fake_aes_8810_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVxp67_ASAP7_75t_SL g4 ( .A(n_1), .Y(n_4) );
BUFx6f_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
INVx5_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AOI22xp33_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_4), .B1(n_1), .B2(n_0), .Y(n_8) );
INVx2_ASAP7_75t_SL g9 ( .A(n_7), .Y(n_9) );
AOI22xp33_ASAP7_75t_L g10 ( .A1(n_8), .A2(n_4), .B1(n_6), .B2(n_5), .Y(n_10) );
NAND3xp33_ASAP7_75t_L g11 ( .A(n_10), .B(n_7), .C(n_5), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_9), .B1(n_7), .B2(n_6), .Y(n_12) );
OAI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_2), .B(n_11), .Y(n_13) );
endmodule