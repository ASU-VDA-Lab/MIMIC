module fake_jpeg_5141_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_8),
.B1(n_3),
.B2(n_5),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_1),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_15),
.B1(n_10),
.B2(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_15),
.B1(n_10),
.B2(n_13),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_27),
.B1(n_33),
.B2(n_26),
.Y(n_38)
);

AO22x1_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_0),
.B1(n_14),
.B2(n_4),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_28),
.B(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.C(n_3),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_34),
.C(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_31),
.B(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_16),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_40),
.B(n_39),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_27),
.B1(n_34),
.B2(n_30),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

AOI21x1_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_45),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_35),
.A3(n_37),
.B1(n_39),
.B2(n_40),
.C1(n_44),
.C2(n_42),
.Y(n_47)
);


endmodule