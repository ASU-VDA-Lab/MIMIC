module fake_jpeg_31449_n_423 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_423);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_423;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_11),
.B(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_14),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_51),
.B(n_26),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_61),
.Y(n_128)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_0),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_67),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_72),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_1),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_86),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_16),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_32),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_18),
.B(n_21),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_84),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_2),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_85),
.B(n_87),
.Y(n_130)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_42),
.B1(n_31),
.B2(n_15),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_93),
.A2(n_102),
.B1(n_113),
.B2(n_125),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_31),
.B1(n_42),
.B2(n_41),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_107),
.B1(n_114),
.B2(n_120),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_2),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_53),
.A2(n_31),
.B1(n_41),
.B2(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_23),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_112),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_34),
.B1(n_25),
.B2(n_39),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_129),
.B1(n_131),
.B2(n_54),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_25),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_62),
.A2(n_40),
.B1(n_28),
.B2(n_38),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_58),
.A2(n_41),
.B1(n_20),
.B2(n_39),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_30),
.B(n_3),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_100),
.C(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_37),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_75),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_47),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_30),
.B1(n_33),
.B2(n_22),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_48),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_52),
.A2(n_22),
.B1(n_33),
.B2(n_5),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_72),
.A2(n_33),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_132),
.B1(n_61),
.B2(n_45),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_57),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_139),
.B(n_150),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_93),
.A2(n_60),
.B1(n_68),
.B2(n_71),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_140),
.A2(n_96),
.B1(n_88),
.B2(n_135),
.Y(n_214)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_143),
.B(n_148),
.Y(n_223)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_145),
.A2(n_149),
.B1(n_158),
.B2(n_170),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_46),
.C(n_79),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_162),
.C(n_128),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_94),
.A2(n_81),
.B1(n_64),
.B2(n_59),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_100),
.B(n_75),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_154),
.Y(n_190)
);

NAND2x1p5_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_115),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_155),
.A2(n_132),
.B(n_97),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_157),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_59),
.B1(n_56),
.B2(n_65),
.Y(n_158)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_56),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_76),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_98),
.B(n_63),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_55),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_172),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_116),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_121),
.A2(n_4),
.B1(n_7),
.B2(n_10),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_173),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_174),
.A2(n_88),
.B1(n_123),
.B2(n_137),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_7),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_12),
.Y(n_201)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_129),
.B(n_131),
.Y(n_187)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_183),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_13),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_11),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_185),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_106),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_187),
.A2(n_159),
.B(n_148),
.Y(n_247)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_130),
.A3(n_108),
.B1(n_128),
.B2(n_122),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_189),
.B(n_161),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_153),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_201),
.B(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_122),
.C(n_101),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_195),
.C(n_147),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_121),
.B1(n_96),
.B2(n_135),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_181),
.B1(n_156),
.B2(n_177),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_117),
.B(n_90),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_216),
.B(n_162),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_214),
.A2(n_152),
.B1(n_137),
.B2(n_179),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_146),
.B(n_117),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_155),
.A2(n_132),
.B(n_90),
.C(n_97),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_150),
.Y(n_245)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_159),
.B1(n_174),
.B2(n_180),
.Y(n_251)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_182),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_132),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_157),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_230),
.B(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_232),
.C(n_236),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_220),
.A2(n_204),
.B(n_208),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_233),
.A2(n_240),
.B(n_245),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_138),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_234),
.B(n_253),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_235),
.A2(n_251),
.B1(n_254),
.B2(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_138),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_238),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_176),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_239),
.B(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_247),
.A2(n_198),
.B1(n_207),
.B2(n_213),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_194),
.A2(n_141),
.B1(n_185),
.B2(n_179),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_139),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_260),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_187),
.A2(n_178),
.B1(n_142),
.B2(n_144),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_178),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_259),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_200),
.A2(n_218),
.B(n_189),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_190),
.B(n_201),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_188),
.B(n_178),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_199),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_199),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_222),
.Y(n_284)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_186),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_160),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_263),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_229),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_292),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_203),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_277),
.C(n_280),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_198),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_190),
.C(n_226),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_187),
.B1(n_217),
.B2(n_214),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_281),
.A2(n_289),
.B1(n_295),
.B2(n_228),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_286),
.B(n_296),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_284),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_244),
.A2(n_217),
.B(n_187),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_234),
.B(n_224),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_287),
.B(n_197),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_215),
.B1(n_210),
.B2(n_205),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_213),
.B1(n_205),
.B2(n_152),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_238),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_246),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_224),
.C(n_197),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_242),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_235),
.A2(n_205),
.B1(n_215),
.B2(n_210),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_258),
.A2(n_227),
.B1(n_197),
.B2(n_196),
.Y(n_296)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_SL g298 ( 
.A(n_267),
.B(n_240),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_317),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_271),
.B(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_233),
.B(n_239),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_300),
.A2(n_303),
.B(n_309),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_237),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_301),
.B(n_307),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_247),
.B(n_261),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_237),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_267),
.A2(n_260),
.B(n_228),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_241),
.Y(n_310)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_250),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_313),
.C(n_274),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_288),
.B1(n_275),
.B2(n_277),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_230),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_314),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_265),
.B(n_249),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_321),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_255),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_318),
.A2(n_289),
.B1(n_295),
.B2(n_275),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_262),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_322),
.B1(n_264),
.B2(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_222),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_269),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_268),
.A2(n_243),
.B(n_206),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_270),
.C(n_222),
.Y(n_347)
);

OAI21x1_ASAP7_75t_SL g324 ( 
.A1(n_300),
.A2(n_283),
.B(n_281),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_339),
.B1(n_346),
.B2(n_310),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_327),
.A2(n_341),
.B1(n_343),
.B2(n_344),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_333),
.C(n_342),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_266),
.C(n_287),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_338),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_302),
.A2(n_268),
.B1(n_291),
.B2(n_280),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_303),
.B1(n_309),
.B2(n_299),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_266),
.C(n_291),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_305),
.A2(n_279),
.B1(n_278),
.B2(n_282),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_307),
.A2(n_279),
.B1(n_278),
.B2(n_282),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_270),
.B1(n_193),
.B2(n_196),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_347),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_311),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_354),
.Y(n_367)
);

INVx11_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_352),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_297),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_358),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_298),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_355),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_314),
.Y(n_357)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_357),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_315),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_332),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_363),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_313),
.C(n_317),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_317),
.C(n_320),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_329),
.Y(n_361)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_298),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_366),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_336),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_340),
.B1(n_310),
.B2(n_327),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_301),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_365),
.B(n_331),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_320),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_350),
.A2(n_337),
.B1(n_325),
.B2(n_349),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_370),
.A2(n_375),
.B1(n_379),
.B2(n_381),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_345),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_373),
.C(n_360),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_325),
.B1(n_334),
.B2(n_345),
.Y(n_375)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_349),
.A2(n_322),
.B1(n_347),
.B2(n_323),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_382),
.B(n_383),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_356),
.C(n_351),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_363),
.C(n_321),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_387),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_375),
.A2(n_357),
.B(n_348),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_386),
.A2(n_390),
.B(n_371),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_368),
.B(n_352),
.Y(n_387)
);

AO22x1_ASAP7_75t_L g388 ( 
.A1(n_381),
.A2(n_348),
.B1(n_362),
.B2(n_366),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_373),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_359),
.B(n_343),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_354),
.C(n_344),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_392),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_376),
.B(n_319),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_374),
.B(n_316),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_393),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_370),
.Y(n_394)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_394),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_389),
.A2(n_369),
.B1(n_359),
.B2(n_355),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_386),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_318),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_308),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_391),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_367),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_403),
.A2(n_377),
.B(n_306),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_407),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_396),
.A2(n_397),
.B(n_402),
.Y(n_405)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_405),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_383),
.C(n_382),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_409),
.B(n_410),
.Y(n_412)
);

AOI322xp5_ASAP7_75t_L g414 ( 
.A1(n_411),
.A2(n_401),
.A3(n_395),
.B1(n_306),
.B2(n_398),
.C1(n_377),
.C2(n_193),
.Y(n_414)
);

AOI221xp5_ASAP7_75t_L g418 ( 
.A1(n_414),
.A2(n_416),
.B1(n_407),
.B2(n_175),
.C(n_12),
.Y(n_418)
);

AOI322xp5_ASAP7_75t_L g416 ( 
.A1(n_408),
.A2(n_160),
.A3(n_175),
.B1(n_209),
.B2(n_97),
.C1(n_166),
.C2(n_206),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_406),
.C(n_404),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_417),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_418),
.A2(n_419),
.B(n_175),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_413),
.Y(n_419)
);

AO21x1_ASAP7_75t_L g422 ( 
.A1(n_421),
.A2(n_415),
.B(n_412),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_420),
.Y(n_423)
);


endmodule