module real_jpeg_2814_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_0),
.B(n_24),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_0),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_0),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_0),
.B(n_55),
.C(n_65),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_0),
.A2(n_35),
.B1(n_37),
.B2(n_92),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_0),
.B(n_52),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_0),
.B(n_102),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_0),
.A2(n_24),
.B(n_77),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_4),
.A2(n_27),
.B1(n_88),
.B2(n_91),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_4),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_4),
.A2(n_27),
.B1(n_54),
.B2(n_55),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_41),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_146)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_60),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_35),
.B1(n_37),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_73),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_83),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_62),
.C(n_74),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_20),
.B(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_42),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_44),
.C(n_49),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_23),
.A2(n_29),
.B1(n_34),
.B2(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_24),
.A2(n_26),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_24),
.A2(n_31),
.A3(n_35),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_47),
.C(n_91),
.Y(n_114)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_26),
.A2(n_48),
.B(n_90),
.C(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_29),
.A2(n_34),
.B1(n_40),
.B2(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OA22x2_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_34),
.B(n_92),
.Y(n_126)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_37),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_35),
.B(n_133),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_87),
.B1(n_93),
.B2(n_95),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_94),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_48),
.B1(n_88),
.B2(n_91),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B(n_58),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_51),
.B(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_51),
.A2(n_80),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_59),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_61),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_52),
.A2(n_61),
.B1(n_92),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_52),
.A2(n_61),
.B1(n_143),
.B2(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_55),
.B(n_141),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_62),
.B(n_74),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B(n_71),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_63),
.A2(n_102),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_102),
.B1(n_128),
.B2(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_67),
.A2(n_69),
.B1(n_99),
.B2(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_75),
.B(n_79),
.Y(n_160)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_103),
.B2(n_104),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_85),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_96),
.CI(n_98),
.CON(n_85),
.SN(n_85)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_167),
.B(n_171),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_156),
.B(n_166),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_137),
.B(n_155),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_130),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_130),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_127),
.C(n_158),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_149),
.B(n_154),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_144),
.B(n_148),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_147),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_153),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_159),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_170),
.Y(n_171)
);


endmodule