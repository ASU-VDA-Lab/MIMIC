module fake_ibex_133_n_873 (n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_873);

input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_873;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_698;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_641;
wire n_557;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_589;
wire n_229;
wire n_209;
wire n_472;
wire n_571;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_741;
wire n_807;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_23),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_28),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_50),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_30),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_55),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_86),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_40),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_48),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_77),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_87),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_52),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_89),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_116),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_63),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_65),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_69),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_62),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_16),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_57),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_97),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_51),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_24),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_94),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_141),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_49),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_68),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_99),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_36),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_39),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_70),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_14),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_44),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_71),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_100),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_84),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_45),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_78),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_112),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_33),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_23),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_13),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_81),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_123),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_106),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_54),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_21),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_24),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_137),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_61),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_128),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_59),
.B(n_43),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_36),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_145),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_120),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_5),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_73),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_133),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_15),
.B(n_76),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_58),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_121),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_66),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_118),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_33),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_131),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_126),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_16),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_188),
.B(n_0),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_183),
.A2(n_231),
.B(n_189),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_194),
.B(n_224),
.Y(n_264)
);

BUFx8_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_214),
.Y(n_266)
);

CKINVDCx6p67_ASAP7_75t_R g267 ( 
.A(n_173),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_180),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_160),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_214),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_180),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_180),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_150),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_199),
.B(n_3),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_4),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_199),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_193),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_164),
.Y(n_282)
);

OAI22x1_ASAP7_75t_R g283 ( 
.A1(n_151),
.A2(n_163),
.B1(n_230),
.B2(n_158),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_152),
.B(n_6),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_154),
.B(n_6),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_193),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_67),
.B(n_149),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_155),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_156),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_245),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_157),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_159),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_151),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_153),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_161),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_162),
.A2(n_166),
.B(n_165),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_167),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_198),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_158),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_163),
.B(n_7),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_152),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_168),
.B(n_8),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_230),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_198),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_175),
.Y(n_309)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_169),
.A2(n_72),
.B(n_148),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_237),
.B(n_10),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_185),
.B(n_12),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_170),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_171),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_198),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_198),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_237),
.B(n_14),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_258),
.B(n_15),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_172),
.A2(n_83),
.B(n_147),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_178),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_174),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_178),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_238),
.B(n_17),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_176),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_164),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_179),
.A2(n_82),
.B(n_146),
.Y(n_326)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_164),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_164),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_184),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_265),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_267),
.Y(n_333)
);

OR2x6_ASAP7_75t_L g334 ( 
.A(n_270),
.B(n_195),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_276),
.B(n_191),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_264),
.B(n_238),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_276),
.B(n_192),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

AND3x1_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_207),
.C(n_202),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_300),
.B(n_196),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_232),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_290),
.B(n_201),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_306),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_263),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_284),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_268),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_300),
.B(n_203),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_267),
.B(n_277),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_262),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_232),
.Y(n_356)
);

NOR3xp33_ASAP7_75t_L g357 ( 
.A(n_307),
.B(n_219),
.C(n_215),
.Y(n_357)
);

OR2x6_ASAP7_75t_L g358 ( 
.A(n_270),
.B(n_208),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_233),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_272),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_233),
.Y(n_362)
);

NAND3x1_ASAP7_75t_L g363 ( 
.A(n_277),
.B(n_229),
.C(n_228),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_312),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_268),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_268),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_273),
.Y(n_367)
);

NOR2x1p5_ASAP7_75t_L g368 ( 
.A(n_292),
.B(n_234),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_312),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_269),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_273),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_284),
.A2(n_223),
.B1(n_204),
.B2(n_225),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_290),
.B(n_205),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_260),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_275),
.B(n_246),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_261),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_273),
.Y(n_382)
);

OR2x6_ASAP7_75t_L g383 ( 
.A(n_296),
.B(n_255),
.Y(n_383)
);

BUFx4f_ASAP7_75t_L g384 ( 
.A(n_291),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_269),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_273),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_283),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_280),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_280),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_278),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_278),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_279),
.B(n_235),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_294),
.B(n_206),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_305),
.A2(n_190),
.B1(n_204),
.B2(n_223),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_278),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_295),
.A2(n_257),
.B1(n_256),
.B2(n_254),
.Y(n_396)
);

AND2x6_ASAP7_75t_L g397 ( 
.A(n_274),
.B(n_212),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_281),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_281),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_281),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_322),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_287),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_281),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_299),
.B(n_213),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_281),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_286),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_286),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_286),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_286),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_272),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_289),
.Y(n_411)
);

AND3x2_ASAP7_75t_L g412 ( 
.A(n_285),
.B(n_250),
.C(n_217),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_320),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_298),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_309),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_299),
.A2(n_221),
.B1(n_253),
.B2(n_252),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_293),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_293),
.Y(n_418)
);

A2O1A1Ixp33_ASAP7_75t_L g419 ( 
.A1(n_347),
.A2(n_313),
.B(n_314),
.C(n_311),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_369),
.A2(n_314),
.B1(n_317),
.B2(n_323),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_346),
.B(n_216),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_336),
.B(n_322),
.Y(n_423)
);

AND2x6_ASAP7_75t_SL g424 ( 
.A(n_383),
.B(n_266),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_384),
.B(n_220),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_344),
.B(n_177),
.Y(n_426)
);

OAI22xp33_ASAP7_75t_L g427 ( 
.A1(n_383),
.A2(n_190),
.B1(n_225),
.B2(n_320),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_356),
.B(n_181),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_384),
.B(n_222),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_353),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_359),
.B(n_182),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_362),
.B(n_186),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_346),
.B(n_226),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_330),
.B(n_187),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_346),
.B(n_236),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_335),
.A2(n_288),
.B(n_310),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_363),
.A2(n_240),
.B1(n_241),
.B2(n_244),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_334),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_355),
.B(n_200),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_333),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_355),
.B(n_209),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_331),
.A2(n_340),
.B1(n_357),
.B2(n_332),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_392),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_339),
.B(n_266),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_332),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_368),
.A2(n_210),
.B1(n_248),
.B2(n_249),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_218),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_348),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_369),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_339),
.B(n_271),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_247),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_360),
.B(n_211),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_379),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_364),
.B(n_288),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_354),
.B(n_271),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_371),
.B(n_288),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_372),
.B(n_377),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_413),
.B(n_394),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_335),
.B(n_338),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_373),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

AOI221xp5_ASAP7_75t_L g466 ( 
.A1(n_347),
.A2(n_282),
.B1(n_325),
.B2(n_328),
.C(n_315),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_401),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_338),
.B(n_310),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_380),
.B(n_18),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_358),
.Y(n_471)
);

AND2x4_ASAP7_75t_SL g472 ( 
.A(n_358),
.B(n_282),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_358),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_342),
.B(n_242),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_342),
.B(n_319),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_342),
.B(n_326),
.Y(n_476)
);

NOR3xp33_ASAP7_75t_L g477 ( 
.A(n_378),
.B(n_18),
.C(n_19),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_361),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_402),
.B(n_20),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_329),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_411),
.B(n_376),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_412),
.B(n_272),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_376),
.A2(n_327),
.B1(n_328),
.B2(n_325),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_418),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_396),
.B(n_308),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_416),
.B(n_308),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_341),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_345),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_416),
.B(n_397),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_345),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_401),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_490),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_440),
.B(n_404),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_457),
.A2(n_349),
.B(n_343),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_387),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_430),
.B(n_387),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_349),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_420),
.B(n_446),
.Y(n_503)
);

NOR3xp33_ASAP7_75t_L g504 ( 
.A(n_427),
.B(n_404),
.C(n_352),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_453),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_458),
.B(n_383),
.Y(n_507)
);

NAND2x1p5_ASAP7_75t_L g508 ( 
.A(n_478),
.B(n_361),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_421),
.B(n_462),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_427),
.B(n_20),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_480),
.A2(n_327),
.B1(n_308),
.B2(n_328),
.Y(n_511)
);

CKINVDCx10_ASAP7_75t_R g512 ( 
.A(n_424),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_470),
.Y(n_513)
);

AO21x1_ASAP7_75t_L g514 ( 
.A1(n_468),
.A2(n_405),
.B(n_365),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_456),
.B(n_22),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_461),
.B(n_25),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_468),
.A2(n_325),
.B(n_328),
.C(n_315),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_464),
.B(n_25),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_455),
.B(n_26),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_472),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

O2A1O1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_419),
.A2(n_408),
.B(n_366),
.C(n_374),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_455),
.B(n_26),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_445),
.A2(n_327),
.B1(n_308),
.B2(n_328),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_475),
.A2(n_480),
.B(n_460),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_434),
.B(n_407),
.C(n_374),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_493),
.A2(n_325),
.B1(n_361),
.B2(n_410),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_452),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_478),
.Y(n_532)
);

BUFx12f_ASAP7_75t_L g533 ( 
.A(n_467),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

AO32x1_ASAP7_75t_L g535 ( 
.A1(n_463),
.A2(n_403),
.A3(n_386),
.B1(n_390),
.B2(n_391),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_471),
.B(n_27),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_469),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_435),
.B(n_27),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_473),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_425),
.A2(n_398),
.B(n_395),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_28),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_429),
.A2(n_403),
.B(n_399),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_429),
.A2(n_405),
.B(n_400),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_422),
.B(n_29),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_442),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_426),
.A2(n_406),
.B(n_409),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_428),
.A2(n_432),
.B(n_431),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_439),
.B(n_31),
.Y(n_548)
);

O2A1O1Ixp33_ASAP7_75t_L g549 ( 
.A1(n_488),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_449),
.B(n_32),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_R g551 ( 
.A(n_482),
.B(n_35),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_433),
.B(n_436),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_433),
.B(n_37),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_436),
.A2(n_297),
.B(n_302),
.C(n_315),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_487),
.A2(n_302),
.B1(n_315),
.B2(n_316),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_484),
.Y(n_556)
);

O2A1O1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_477),
.A2(n_38),
.B(n_41),
.C(n_42),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_481),
.B(n_41),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_450),
.A2(n_454),
.B(n_438),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_486),
.B(n_42),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_491),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_479),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_441),
.B(n_302),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_489),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_444),
.A2(n_382),
.B(n_370),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_477),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_485),
.A2(n_466),
.B1(n_316),
.B2(n_315),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_532),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g570 ( 
.A1(n_552),
.A2(n_523),
.B(n_519),
.Y(n_570)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_559),
.A2(n_370),
.B(n_367),
.C(n_351),
.Y(n_571)
);

OAI21x1_ASAP7_75t_SL g572 ( 
.A1(n_509),
.A2(n_46),
.B(n_47),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_527),
.A2(n_337),
.B(n_56),
.Y(n_573)
);

NAND3x1_ASAP7_75t_L g574 ( 
.A(n_512),
.B(n_53),
.C(n_60),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_534),
.B(n_537),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_541),
.A2(n_544),
.B(n_553),
.C(n_538),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_516),
.A2(n_510),
.B1(n_518),
.B2(n_515),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_548),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_560),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_525),
.A2(n_111),
.B(n_113),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

AOI21xp33_ASAP7_75t_L g582 ( 
.A1(n_549),
.A2(n_558),
.B(n_522),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_562),
.A2(n_124),
.B(n_129),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_502),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_513),
.B(n_507),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_566),
.A2(n_546),
.B(n_540),
.Y(n_586)
);

OA21x2_ASAP7_75t_L g587 ( 
.A1(n_554),
.A2(n_543),
.B(n_542),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_497),
.B(n_505),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_497),
.B(n_550),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_502),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g591 ( 
.A(n_520),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_500),
.B(n_530),
.Y(n_592)
);

AO31x2_ASAP7_75t_L g593 ( 
.A1(n_568),
.A2(n_555),
.A3(n_563),
.B(n_531),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_495),
.B(n_539),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_524),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_512),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_501),
.A2(n_506),
.B1(n_536),
.B2(n_561),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_532),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_565),
.A2(n_535),
.B(n_496),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_502),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_496),
.A2(n_526),
.B1(n_564),
.B2(n_545),
.Y(n_601)
);

NOR2x1_ASAP7_75t_SL g602 ( 
.A(n_532),
.B(n_521),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_506),
.B(n_496),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_508),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_551),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_535),
.A2(n_320),
.B1(n_322),
.B2(n_375),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_535),
.B(n_503),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_503),
.B(n_420),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_503),
.B(n_430),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_503),
.B(n_420),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_498),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_430),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_498),
.B(n_503),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_498),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_430),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_527),
.A2(n_499),
.B(n_468),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_503),
.B(n_447),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

AO22x2_ASAP7_75t_L g619 ( 
.A1(n_510),
.A2(n_413),
.B1(n_516),
.B2(n_513),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

AO32x2_ASAP7_75t_L g621 ( 
.A1(n_568),
.A2(n_529),
.A3(n_279),
.B1(n_511),
.B2(n_556),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_498),
.Y(n_622)
);

AOI211x1_ASAP7_75t_L g623 ( 
.A1(n_509),
.A2(n_552),
.B(n_541),
.C(n_544),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_533),
.Y(n_624)
);

O2A1O1Ixp5_ASAP7_75t_L g625 ( 
.A1(n_514),
.A2(n_474),
.B(n_517),
.C(n_519),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_498),
.B(n_503),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_498),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_503),
.B(n_420),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_499),
.A2(n_476),
.B(n_459),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_498),
.B(n_503),
.Y(n_630)
);

AOI221x1_ASAP7_75t_L g631 ( 
.A1(n_517),
.A2(n_504),
.B1(n_528),
.B2(n_477),
.C(n_437),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_499),
.A2(n_476),
.B(n_459),
.Y(n_632)
);

AOI221x1_ASAP7_75t_L g633 ( 
.A1(n_517),
.A2(n_504),
.B1(n_528),
.B2(n_477),
.C(n_437),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_503),
.B(n_430),
.Y(n_634)
);

O2A1O1Ixp5_ASAP7_75t_L g635 ( 
.A1(n_514),
.A2(n_474),
.B(n_517),
.C(n_519),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_527),
.A2(n_499),
.B(n_468),
.Y(n_636)
);

INVx6_ASAP7_75t_L g637 ( 
.A(n_533),
.Y(n_637)
);

AOI221x1_ASAP7_75t_L g638 ( 
.A1(n_517),
.A2(n_504),
.B1(n_528),
.B2(n_477),
.C(n_437),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_SL g640 ( 
.A(n_551),
.B(n_401),
.C(n_467),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_498),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_503),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_503),
.B(n_420),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_500),
.B(n_434),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_521),
.Y(n_645)
);

AO22x2_ASAP7_75t_L g646 ( 
.A1(n_510),
.A2(n_413),
.B1(n_516),
.B2(n_513),
.Y(n_646)
);

OAI21x1_ASAP7_75t_SL g647 ( 
.A1(n_509),
.A2(n_547),
.B(n_518),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_503),
.B(n_420),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_532),
.Y(n_649)
);

OAI21x1_ASAP7_75t_SL g650 ( 
.A1(n_602),
.A2(n_583),
.B(n_580),
.Y(n_650)
);

OA21x2_ASAP7_75t_L g651 ( 
.A1(n_631),
.A2(n_638),
.B(n_633),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_598),
.B(n_604),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_598),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_608),
.B(n_610),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_611),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_614),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_628),
.B(n_643),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_618),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_598),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_648),
.B(n_609),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_576),
.A2(n_625),
.B(n_635),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_SL g662 ( 
.A1(n_619),
.A2(n_646),
.B1(n_605),
.B2(n_601),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_612),
.B(n_615),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_570),
.A2(n_592),
.B(n_607),
.Y(n_664)
);

OA21x2_ASAP7_75t_L g665 ( 
.A1(n_616),
.A2(n_636),
.B(n_586),
.Y(n_665)
);

BUFx2_ASAP7_75t_SL g666 ( 
.A(n_581),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_642),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_634),
.B(n_613),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_620),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_644),
.B(n_626),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_577),
.A2(n_619),
.B1(n_646),
.B2(n_589),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_594),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_569),
.B(n_649),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_570),
.A2(n_632),
.B(n_629),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_630),
.B(n_617),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_591),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_639),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_595),
.B(n_645),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_585),
.B(n_588),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_622),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_627),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_587),
.Y(n_682)
);

OAI21xp33_ASAP7_75t_L g683 ( 
.A1(n_577),
.A2(n_582),
.B(n_578),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_575),
.B(n_641),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_597),
.B(n_623),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_623),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_601),
.A2(n_578),
.B1(n_605),
.B2(n_606),
.Y(n_687)
);

BUFx2_ASAP7_75t_SL g688 ( 
.A(n_620),
.Y(n_688)
);

OAI21x1_ASAP7_75t_SL g689 ( 
.A1(n_579),
.A2(n_590),
.B(n_600),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_640),
.A2(n_603),
.B1(n_600),
.B2(n_584),
.Y(n_690)
);

NAND2x1_ASAP7_75t_L g691 ( 
.A(n_637),
.B(n_574),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_621),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_621),
.A2(n_593),
.B(n_624),
.Y(n_693)
);

AO21x2_ASAP7_75t_L g694 ( 
.A1(n_596),
.A2(n_607),
.B(n_599),
.Y(n_694)
);

BUFx2_ASAP7_75t_R g695 ( 
.A(n_596),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_576),
.A2(n_552),
.B(n_527),
.Y(n_696)
);

AO31x2_ASAP7_75t_L g697 ( 
.A1(n_631),
.A2(n_638),
.A3(n_633),
.B(n_514),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_598),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_642),
.B(n_447),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_570),
.A2(n_576),
.B(n_557),
.C(n_582),
.Y(n_700)
);

OAI21x1_ASAP7_75t_SL g701 ( 
.A1(n_602),
.A2(n_583),
.B(n_580),
.Y(n_701)
);

CKINVDCx6p67_ASAP7_75t_R g702 ( 
.A(n_624),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_598),
.Y(n_703)
);

NOR2x1_ASAP7_75t_SL g704 ( 
.A(n_598),
.B(n_532),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_608),
.B(n_610),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_609),
.B(n_612),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_598),
.B(n_602),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_609),
.B(n_612),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_598),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_576),
.A2(n_552),
.B(n_527),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_608),
.B(n_610),
.Y(n_711)
);

AOI22x1_ASAP7_75t_L g712 ( 
.A1(n_647),
.A2(n_572),
.B1(n_573),
.B2(n_547),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_576),
.A2(n_570),
.B(n_571),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_611),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_577),
.A2(n_510),
.B1(n_567),
.B2(n_619),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_642),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_707),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_655),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_660),
.B(n_706),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_706),
.B(n_663),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_658),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_700),
.A2(n_696),
.B(n_710),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_682),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_708),
.B(n_654),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_686),
.Y(n_726)
);

AO21x2_ASAP7_75t_L g727 ( 
.A1(n_661),
.A2(n_713),
.B(n_674),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_677),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_668),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_677),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_657),
.B(n_705),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_665),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_680),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_667),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_681),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_707),
.B(n_703),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_716),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_714),
.Y(n_738)
);

INVxp33_ASAP7_75t_L g739 ( 
.A(n_652),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_666),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_715),
.A2(n_671),
.B1(n_662),
.B2(n_711),
.Y(n_741)
);

INVxp33_ASAP7_75t_L g742 ( 
.A(n_652),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_652),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_675),
.B(n_715),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_684),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_670),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_671),
.B(n_699),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_659),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_659),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_709),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_692),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_685),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_650),
.B(n_701),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_664),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_691),
.B(n_689),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_679),
.B(n_672),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_687),
.A2(n_683),
.B1(n_709),
.B2(n_690),
.Y(n_757)
);

INVxp33_ASAP7_75t_L g758 ( 
.A(n_704),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_698),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_653),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_693),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_673),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_753),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_723),
.B(n_754),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_751),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_754),
.B(n_651),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_752),
.B(n_700),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_744),
.B(n_697),
.Y(n_768)
);

BUFx12f_ASAP7_75t_L g769 ( 
.A(n_748),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_724),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_731),
.B(n_678),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_748),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_728),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_753),
.B(n_694),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_727),
.B(n_732),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_730),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_749),
.Y(n_777)
);

NOR2x1_ASAP7_75t_L g778 ( 
.A(n_755),
.B(n_688),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_741),
.A2(n_702),
.B1(n_669),
.B2(n_690),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_753),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_771),
.B(n_746),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_764),
.B(n_761),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_771),
.B(n_747),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_764),
.B(n_718),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_772),
.B(n_769),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_765),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_764),
.B(n_766),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_778),
.B(n_717),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_767),
.B(n_726),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_767),
.B(n_745),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_765),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_766),
.B(n_761),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_772),
.B(n_717),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_768),
.B(n_719),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_777),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_770),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_777),
.B(n_721),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_787),
.B(n_775),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_787),
.B(n_773),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_782),
.B(n_792),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_784),
.B(n_773),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_786),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_786),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_794),
.B(n_768),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_782),
.B(n_775),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_790),
.B(n_776),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_790),
.B(n_776),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_795),
.Y(n_808)
);

NAND4xp25_ASAP7_75t_L g809 ( 
.A(n_783),
.B(n_779),
.C(n_778),
.D(n_725),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_791),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_792),
.B(n_774),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_794),
.B(n_768),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_796),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_802),
.Y(n_814)
);

AOI32xp33_ASAP7_75t_SL g815 ( 
.A1(n_808),
.A2(n_797),
.A3(n_720),
.B1(n_781),
.B2(n_750),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_809),
.B(n_740),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_813),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_799),
.B(n_796),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_802),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_813),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_803),
.Y(n_821)
);

NAND3x1_ASAP7_75t_SL g822 ( 
.A(n_800),
.B(n_702),
.C(n_769),
.Y(n_822)
);

OAI21xp33_ASAP7_75t_L g823 ( 
.A1(n_806),
.A2(n_779),
.B(n_734),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_803),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_810),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_816),
.B(n_695),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_817),
.A2(n_793),
.B1(n_755),
.B2(n_763),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_818),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_817),
.B(n_800),
.Y(n_829)
);

AOI322xp5_ASAP7_75t_L g830 ( 
.A1(n_823),
.A2(n_798),
.A3(n_805),
.B1(n_812),
.B2(n_811),
.C1(n_807),
.C2(n_801),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_820),
.B(n_769),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_823),
.A2(n_811),
.B1(n_805),
.B2(n_804),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_814),
.B(n_798),
.Y(n_833)
);

AOI31xp33_ASAP7_75t_L g834 ( 
.A1(n_822),
.A2(n_785),
.A3(n_788),
.B(n_758),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_815),
.A2(n_793),
.B(n_737),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_819),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_825),
.B(n_804),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_837),
.Y(n_838)
);

AOI21xp33_ASAP7_75t_L g839 ( 
.A1(n_835),
.A2(n_760),
.B(n_759),
.Y(n_839)
);

AOI21xp33_ASAP7_75t_L g840 ( 
.A1(n_826),
.A2(n_755),
.B(n_772),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_834),
.A2(n_755),
.B(n_811),
.Y(n_841)
);

OAI221xp5_ASAP7_75t_L g842 ( 
.A1(n_832),
.A2(n_763),
.B1(n_824),
.B2(n_821),
.C(n_788),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_833),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_838),
.B(n_830),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_L g845 ( 
.A(n_839),
.B(n_834),
.C(n_836),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_843),
.B(n_828),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_844),
.B(n_842),
.Y(n_847)
);

AOI32xp33_ASAP7_75t_L g848 ( 
.A1(n_846),
.A2(n_829),
.A3(n_827),
.B1(n_763),
.B2(n_736),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_848),
.B(n_845),
.Y(n_849)
);

NAND4xp75_ASAP7_75t_L g850 ( 
.A(n_847),
.B(n_841),
.C(n_831),
.D(n_840),
.Y(n_850)
);

NOR2x1p5_ASAP7_75t_L g851 ( 
.A(n_850),
.B(n_676),
.Y(n_851)
);

AOI32xp33_ASAP7_75t_L g852 ( 
.A1(n_849),
.A2(n_676),
.A3(n_742),
.B1(n_739),
.B2(n_757),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_851),
.B(n_810),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_852),
.B(n_669),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_853),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_854),
.Y(n_856)
);

AO22x2_ASAP7_75t_L g857 ( 
.A1(n_854),
.A2(n_762),
.B1(n_731),
.B2(n_756),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_856),
.B(n_729),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_855),
.B(n_719),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_857),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_857),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_861),
.A2(n_860),
.B(n_858),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_859),
.B(n_789),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_858),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_860),
.A2(n_736),
.B(n_722),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_861),
.A2(n_673),
.B(n_735),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_858),
.A2(n_717),
.B1(n_743),
.B2(n_780),
.Y(n_867)
);

OAI31xp33_ASAP7_75t_SL g868 ( 
.A1(n_862),
.A2(n_733),
.A3(n_738),
.B(n_712),
.Y(n_868)
);

OAI21x1_ASAP7_75t_L g869 ( 
.A1(n_864),
.A2(n_756),
.B(n_788),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_863),
.B(n_865),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_870),
.B(n_866),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_871),
.B(n_869),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_872),
.A2(n_867),
.B1(n_868),
.B2(n_743),
.Y(n_873)
);


endmodule