module fake_jpeg_12225_n_197 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_14),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_11),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_68),
.Y(n_96)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_84),
.B1(n_67),
.B2(n_71),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_101),
.C(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_65),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_69),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_60),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_67),
.B1(n_71),
.B2(n_55),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

OR2x2_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_76),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_55),
.B1(n_81),
.B2(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_93),
.B1(n_91),
.B2(n_57),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_121),
.B1(n_30),
.B2(n_53),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_78),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_115),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_63),
.B(n_72),
.C(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_117),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_123),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_57),
.B1(n_81),
.B2(n_76),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_109),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_61),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_127),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_75),
.Y(n_127)
);

HAxp5_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_77),
.CON(n_137),
.SN(n_137)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_82),
.Y(n_136)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_56),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_153),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_13),
.B(n_14),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_118),
.B(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_26),
.B(n_42),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_66),
.C(n_73),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_142),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_79),
.B1(n_64),
.B2(n_62),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_147),
.B1(n_150),
.B2(n_7),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_70),
.B1(n_1),
.B2(n_2),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_151),
.B1(n_15),
.B2(n_16),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_7),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_27),
.B1(n_51),
.B2(n_45),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_163),
.B(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_161),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_160),
.B(n_169),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_9),
.B(n_10),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_32),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_133),
.C(n_31),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_132),
.B(n_13),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_167),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_170),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_15),
.B(n_17),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_21),
.B(n_22),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_139),
.A3(n_140),
.B1(n_154),
.B2(n_134),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_157),
.B1(n_169),
.B2(n_159),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_175),
.B(n_176),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_133),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_156),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_184),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_181),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_186),
.C(n_180),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_157),
.B(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_176),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_189),
.C(n_175),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_177),
.B(n_184),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_187),
.B1(n_178),
.B2(n_179),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_182),
.C(n_165),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_25),
.B(n_33),
.C(n_34),
.D(n_35),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_41),
.Y(n_197)
);


endmodule