module fake_netlist_6_836_n_1702 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1702);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1702;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_14),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_27),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_77),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_30),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_93),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_66),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_67),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_49),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_96),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_74),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_118),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_5),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_51),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_45),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_20),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_41),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_35),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_44),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_58),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_60),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_46),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_57),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_92),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_89),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_111),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_62),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_59),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_17),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_141),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_87),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_46),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_25),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_0),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_134),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_161),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_112),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_119),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_53),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_45),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_12),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_11),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_129),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_81),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_21),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_36),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_6),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_68),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_128),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_6),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_54),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_100),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_28),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_36),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_104),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_27),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_65),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_39),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_102),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_144),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_32),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_122),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_22),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_23),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_8),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_56),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_88),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_95),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_37),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_108),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_40),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_132),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_78),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_35),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_5),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_30),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_135),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_103),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_53),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_15),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_85),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_70),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_72),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_75),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_32),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_105),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_33),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_16),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_13),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_116),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_42),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_99),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_101),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_114),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_48),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_94),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_33),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_130),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_71),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_98),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_84),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_20),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_109),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_41),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_113),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_138),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_73),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_26),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_10),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_51),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_25),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_133),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_159),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_1),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_79),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_139),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_12),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_48),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_54),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_34),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_49),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_37),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_146),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_147),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_154),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_7),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_17),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_14),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_160),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_39),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_258),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_163),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_165),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_165),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_211),
.B(n_1),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_184),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_165),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_165),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_164),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_165),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_250),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_165),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_166),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_165),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_168),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_169),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_190),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_170),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_190),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_190),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_190),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_190),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_190),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_166),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_190),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_171),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_194),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_194),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_251),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_251),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_251),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_183),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_220),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_251),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_175),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_249),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_188),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_215),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_251),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_220),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_251),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_251),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_249),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_189),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_191),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_222),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_211),
.B(n_3),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_180),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_203),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_203),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_203),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_203),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_225),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_225),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_225),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_225),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_234),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_234),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_222),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_234),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_234),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_285),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_192),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_246),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_244),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_193),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_248),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_198),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_248),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_285),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_181),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_274),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_244),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_244),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_200),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_321),
.B(n_290),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_322),
.B(n_323),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_335),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_356),
.B(n_236),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_322),
.A2(n_326),
.B(n_323),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_329),
.B(n_368),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_336),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_290),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_346),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_355),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_374),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_357),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_374),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_173),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_236),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_333),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_282),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_174),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_344),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_328),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_347),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_364),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_330),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g437 ( 
.A(n_331),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_365),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_331),
.B(n_274),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_348),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_330),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_380),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_352),
.B(n_183),
.Y(n_449)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_332),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_353),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_360),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_332),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_386),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_366),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_325),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_379),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_177),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_384),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_R g464 ( 
.A(n_391),
.B(n_178),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_387),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_R g466 ( 
.A(n_395),
.B(n_202),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_390),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_396),
.B(n_327),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_176),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_389),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_407),
.B(n_324),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_422),
.Y(n_475)
);

BUFx4f_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_417),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_405),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_416),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_416),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_385),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_450),
.B(n_176),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_431),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_367),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_401),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_431),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

INVx4_ASAP7_75t_SL g489 ( 
.A(n_455),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_403),
.B(n_418),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_418),
.B(n_393),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_431),
.B(n_394),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

NAND3x1_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_172),
.C(n_167),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_450),
.B(n_415),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_450),
.B(n_415),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_446),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_404),
.A2(n_282),
.B1(n_182),
.B2(n_187),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_446),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_334),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_404),
.A2(n_247),
.B1(n_185),
.B2(n_273),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_450),
.B(n_334),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_455),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_411),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_455),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_176),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_464),
.B(n_207),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_411),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_400),
.A2(n_179),
.B1(n_178),
.B2(n_240),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

OAI22xp33_ASAP7_75t_L g516 ( 
.A1(n_450),
.A2(n_306),
.B1(n_319),
.B2(n_262),
.Y(n_516)
);

BUFx6f_ASAP7_75t_SL g517 ( 
.A(n_415),
.Y(n_517)
);

BUFx4f_ASAP7_75t_L g518 ( 
.A(n_404),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_450),
.B(n_176),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_441),
.B(n_197),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_406),
.B(n_337),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_446),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_415),
.B(n_268),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_413),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_337),
.Y(n_525)
);

INVx4_ASAP7_75t_SL g526 ( 
.A(n_398),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_428),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_410),
.A2(n_179),
.B1(n_240),
.B2(n_313),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_398),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_398),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_399),
.B(n_339),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_399),
.B(n_409),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_428),
.B(n_268),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_409),
.B(n_339),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_340),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_428),
.A2(n_201),
.B1(n_204),
.B2(n_199),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

INVx6_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_425),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_397),
.B(n_340),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_426),
.B(n_268),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_414),
.B(n_341),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_466),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_426),
.A2(n_292),
.B1(n_218),
.B2(n_230),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_443),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_414),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_436),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_397),
.B(n_268),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_434),
.B(n_196),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_440),
.B(n_223),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_456),
.B(n_341),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_419),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_421),
.B(n_342),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_421),
.B(n_342),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_398),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_427),
.B(n_343),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_436),
.B(n_235),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_423),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_452),
.B(n_343),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_437),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_430),
.B(n_345),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_452),
.B(n_252),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_452),
.B(n_264),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_437),
.B(n_208),
.C(n_186),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_435),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_435),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_398),
.B(n_265),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_438),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_398),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_402),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_438),
.B(n_345),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_439),
.A2(n_275),
.B1(n_216),
.B2(n_299),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_402),
.B(n_349),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_439),
.Y(n_585)
);

INVx8_ASAP7_75t_L g586 ( 
.A(n_429),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_465),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_445),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_445),
.B(n_349),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_447),
.B(n_350),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_402),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_447),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_402),
.B(n_350),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_448),
.Y(n_595)
);

BUFx4f_ASAP7_75t_L g596 ( 
.A(n_451),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_459),
.A2(n_232),
.B1(n_318),
.B2(n_314),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_402),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_432),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_459),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_402),
.B(n_351),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_460),
.B(n_244),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_443),
.B(n_351),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_444),
.B(n_281),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_453),
.B(n_296),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_454),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_457),
.B(n_284),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_461),
.B(n_361),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_463),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_416),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_491),
.B(n_287),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_468),
.B(n_195),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_473),
.B(n_293),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_473),
.B(n_294),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_498),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_468),
.B(n_209),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_490),
.B(n_295),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_476),
.B(n_300),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_480),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_476),
.A2(n_518),
.B(n_502),
.C(n_505),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_531),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_512),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_467),
.B(n_481),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_512),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_505),
.B(n_305),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_467),
.B(n_312),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_518),
.B(n_205),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_568),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_467),
.B(n_612),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_601),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_544),
.Y(n_636)
);

BUFx8_ASAP7_75t_L g637 ( 
.A(n_608),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_521),
.B(n_362),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_502),
.B(n_206),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_525),
.B(n_210),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_475),
.B(n_392),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_544),
.Y(n_642)
);

O2A1O1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_567),
.A2(n_317),
.B(n_316),
.C(n_315),
.Y(n_643)
);

INVx6_ASAP7_75t_L g644 ( 
.A(n_595),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_540),
.B(n_213),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_559),
.B(n_214),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_469),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_491),
.B(n_217),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_514),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_499),
.Y(n_650)
);

INVxp33_ASAP7_75t_L g651 ( 
.A(n_472),
.Y(n_651)
);

BUFx8_ASAP7_75t_L g652 ( 
.A(n_608),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_567),
.A2(n_315),
.B(n_308),
.C(n_291),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_499),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_491),
.B(n_221),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_514),
.B(n_224),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_508),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_506),
.B(n_228),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_469),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_L g660 ( 
.A1(n_541),
.A2(n_219),
.B1(n_310),
.B2(n_309),
.C(n_307),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_508),
.B(n_524),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_524),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_477),
.B(n_311),
.C(n_227),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_554),
.B(n_231),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_527),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_527),
.B(n_229),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_484),
.A2(n_241),
.B1(n_304),
.B2(n_243),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_550),
.B(n_207),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_511),
.B(n_238),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_469),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_529),
.B(n_237),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_541),
.A2(n_551),
.B1(n_590),
.B2(n_562),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_595),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_543),
.B(n_226),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_610),
.B(n_215),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_605),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_599),
.A2(n_270),
.B(n_303),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_579),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_586),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_605),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_605),
.Y(n_683)
);

BUFx5_ASAP7_75t_L g684 ( 
.A(n_483),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_551),
.A2(n_308),
.B1(n_263),
.B2(n_233),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_577),
.B(n_239),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_536),
.A2(n_283),
.B(n_271),
.C(n_297),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_588),
.B(n_242),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_600),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_520),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_478),
.B(n_215),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_568),
.B(n_254),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_471),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_562),
.A2(n_263),
.B1(n_226),
.B2(n_291),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_543),
.B(n_571),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_478),
.B(n_233),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_520),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_573),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_469),
.B(n_255),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_592),
.B(n_259),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_594),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_597),
.B(n_260),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_471),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_485),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_604),
.B(n_261),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_487),
.B(n_266),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_562),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_497),
.B(n_276),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_557),
.B(n_245),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_557),
.B(n_253),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_590),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_484),
.A2(n_277),
.B1(n_301),
.B2(n_289),
.Y(n_712)
);

CKINVDCx11_ASAP7_75t_R g713 ( 
.A(n_586),
.Y(n_713)
);

AND2x2_ASAP7_75t_SL g714 ( 
.A(n_583),
.B(n_590),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_501),
.B(n_278),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_495),
.A2(n_500),
.B(n_584),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_485),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_586),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_486),
.Y(n_719)
);

AO221x1_ASAP7_75t_L g720 ( 
.A1(n_516),
.A2(n_183),
.B1(n_212),
.B2(n_267),
.C(n_9),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_596),
.B(n_503),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_591),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_478),
.B(n_269),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_484),
.A2(n_286),
.B1(n_280),
.B2(n_212),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_558),
.B(n_576),
.Y(n_725)
);

INVxp33_ASAP7_75t_SL g726 ( 
.A(n_569),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_522),
.B(n_302),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_532),
.B(n_288),
.C(n_279),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_486),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_558),
.B(n_513),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_SL g731 ( 
.A(n_552),
.B(n_587),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_563),
.B(n_272),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_488),
.Y(n_733)
);

BUFx6f_ASAP7_75t_SL g734 ( 
.A(n_607),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_520),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_560),
.B(n_267),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_511),
.B(n_256),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_530),
.Y(n_738)
);

NOR3xp33_ASAP7_75t_L g739 ( 
.A(n_606),
.B(n_257),
.C(n_267),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_575),
.A2(n_212),
.B1(n_7),
.B2(n_8),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_572),
.B(n_61),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_488),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_606),
.B(n_4),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_560),
.B(n_561),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_561),
.Y(n_745)
);

OAI221xp5_ASAP7_75t_L g746 ( 
.A1(n_583),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.C(n_18),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_582),
.B(n_82),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_493),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_561),
.B(n_69),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_537),
.B(n_83),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_537),
.B(n_536),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_539),
.B(n_63),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_591),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_493),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_496),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_591),
.Y(n_756)
);

AO22x1_ASAP7_75t_L g757 ( 
.A1(n_470),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_530),
.Y(n_758)
);

AND3x1_ASAP7_75t_L g759 ( 
.A(n_611),
.B(n_19),
.C(n_23),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_565),
.B(n_24),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_565),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_603),
.B(n_106),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_SL g763 ( 
.A1(n_539),
.A2(n_97),
.B(n_153),
.C(n_152),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_548),
.B(n_90),
.Y(n_764)
);

NOR2x1p5_ASAP7_75t_L g765 ( 
.A(n_611),
.B(n_24),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_609),
.B(n_28),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_609),
.B(n_607),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_470),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_565),
.B(n_29),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_517),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_504),
.B(n_117),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_598),
.B(n_482),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_470),
.A2(n_31),
.B1(n_38),
.B2(n_42),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_517),
.B(n_38),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_548),
.B(n_589),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_533),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_628),
.A2(n_625),
.B(n_661),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_615),
.B(n_607),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_751),
.B(n_566),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_615),
.A2(n_766),
.B(n_743),
.C(n_730),
.Y(n_780)
);

NOR2x1_ASAP7_75t_L g781 ( 
.A(n_745),
.B(n_500),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_775),
.B(n_566),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_641),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_625),
.A2(n_495),
.B1(n_494),
.B2(n_538),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_638),
.B(n_589),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_676),
.B(n_538),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_714),
.B(n_591),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_632),
.A2(n_519),
.B(n_546),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_730),
.A2(n_519),
.B1(n_580),
.B2(n_581),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_621),
.B(n_725),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_716),
.A2(n_534),
.B(n_509),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_635),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_613),
.B(n_581),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_636),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_672),
.A2(n_580),
.B1(n_578),
.B2(n_492),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_617),
.B(n_470),
.Y(n_796)
);

AOI21xp33_ASAP7_75t_L g797 ( 
.A1(n_621),
.A2(n_578),
.B(n_602),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_623),
.A2(n_593),
.B(n_549),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_714),
.B(n_564),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_623),
.A2(n_474),
.B(n_507),
.Y(n_800)
);

AO32x1_ASAP7_75t_L g801 ( 
.A1(n_620),
.A2(n_553),
.A3(n_555),
.B1(n_545),
.B2(n_542),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_664),
.B(n_574),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_632),
.A2(n_528),
.B(n_570),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_633),
.A2(n_474),
.B(n_507),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_634),
.A2(n_474),
.B(n_515),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_630),
.B(n_564),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_709),
.A2(n_535),
.B(n_496),
.C(n_556),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_619),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_630),
.B(n_535),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_721),
.A2(n_507),
.B(n_515),
.Y(n_810)
);

AND2x2_ASAP7_75t_SL g811 ( 
.A(n_762),
.B(n_510),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_741),
.A2(n_526),
.B(n_489),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_619),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_747),
.A2(n_526),
.B(n_489),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_709),
.A2(n_573),
.B(n_523),
.C(n_489),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_689),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_636),
.Y(n_817)
);

O2A1O1Ixp5_ASAP7_75t_L g818 ( 
.A1(n_622),
.A2(n_573),
.B(n_523),
.C(n_547),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_750),
.A2(n_523),
.B(n_573),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_627),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_639),
.A2(n_573),
.B(n_523),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_722),
.A2(n_523),
.B(n_547),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_710),
.B(n_43),
.C(n_44),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_707),
.A2(n_547),
.B1(n_136),
.B2(n_140),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_691),
.B(n_47),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_710),
.A2(n_47),
.B(n_50),
.C(n_52),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_743),
.B(n_766),
.C(n_685),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_643),
.A2(n_50),
.B(n_52),
.C(n_55),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_669),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_772),
.A2(n_711),
.B1(n_642),
.B2(n_683),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_746),
.A2(n_110),
.B(n_121),
.C(n_124),
.Y(n_831)
);

AOI21xp33_ASAP7_75t_L g832 ( 
.A1(n_737),
.A2(n_125),
.B(n_143),
.Y(n_832)
);

AND2x4_ASAP7_75t_SL g833 ( 
.A(n_745),
.B(n_145),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_752),
.A2(n_148),
.B(n_150),
.C(n_155),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_756),
.A2(n_683),
.B(n_681),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_636),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_677),
.A2(n_681),
.B(n_692),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_639),
.A2(n_764),
.B(n_649),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_679),
.B(n_682),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_629),
.A2(n_649),
.B(n_631),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_693),
.A2(n_717),
.B(n_703),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_650),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_701),
.B(n_761),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_677),
.A2(n_658),
.B(n_656),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_L g845 ( 
.A(n_636),
.B(n_670),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_654),
.A2(n_675),
.B1(n_665),
.B2(n_657),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_613),
.A2(n_626),
.B1(n_662),
.B2(n_761),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_R g848 ( 
.A(n_713),
.B(n_674),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_626),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_732),
.B(n_640),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_645),
.B(n_646),
.Y(n_851)
);

AO22x1_ASAP7_75t_L g852 ( 
.A1(n_739),
.A2(n_769),
.B1(n_774),
.B2(n_760),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_753),
.A2(n_671),
.B(n_666),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_693),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_753),
.A2(n_708),
.B(n_706),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_723),
.B(n_673),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_624),
.B(n_614),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_651),
.B(n_744),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_703),
.A2(n_742),
.B(n_704),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_685),
.B(n_644),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_753),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_768),
.A2(n_773),
.B1(n_648),
.B2(n_655),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_753),
.A2(n_715),
.B(n_670),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_738),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_614),
.B(n_776),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_684),
.B(n_749),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_687),
.B(n_769),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_690),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_653),
.A2(n_724),
.B(n_727),
.C(n_712),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_644),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_644),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_647),
.A2(n_659),
.B(n_699),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_667),
.B(n_740),
.C(n_736),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_647),
.A2(n_659),
.B(n_699),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_717),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_768),
.A2(n_773),
.B1(n_762),
.B2(n_705),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_700),
.A2(n_702),
.B(n_688),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_719),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_719),
.B(n_742),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_767),
.B(n_668),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_694),
.B(n_696),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_686),
.A2(n_771),
.B(n_698),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_697),
.B(n_735),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_729),
.B(n_754),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_729),
.A2(n_733),
.B(n_755),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_733),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_748),
.B(n_755),
.Y(n_888)
);

NOR2x1p5_ASAP7_75t_SL g889 ( 
.A(n_684),
.B(n_748),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_774),
.A2(n_660),
.B(n_728),
.C(n_694),
.Y(n_890)
);

NOR2x1_ASAP7_75t_R g891 ( 
.A(n_680),
.B(n_718),
.Y(n_891)
);

NOR2x1_ASAP7_75t_L g892 ( 
.A(n_680),
.B(n_718),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_684),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_695),
.B(n_731),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_765),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_763),
.A2(n_678),
.B(n_663),
.C(n_720),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_757),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_759),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_726),
.B(n_770),
.Y(n_899)
);

NOR2x1_ASAP7_75t_L g900 ( 
.A(n_770),
.B(n_637),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_637),
.A2(n_652),
.B(n_734),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_652),
.Y(n_902)
);

OAI321xp33_ASAP7_75t_L g903 ( 
.A1(n_734),
.A2(n_615),
.A3(n_766),
.B1(n_743),
.B2(n_746),
.C(n_621),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_689),
.B(n_477),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_625),
.A2(n_518),
.B(n_476),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_L g906 ( 
.A(n_615),
.B(n_621),
.C(n_511),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_615),
.A2(n_621),
.B(n_730),
.C(n_473),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_632),
.A2(n_661),
.B(n_721),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_615),
.A2(n_730),
.B1(n_621),
.B2(n_714),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_650),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_618),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_751),
.B(n_775),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_751),
.B(n_775),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_625),
.B(n_714),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_628),
.A2(n_518),
.B(n_476),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_632),
.A2(n_661),
.B(n_721),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_L g917 ( 
.A(n_615),
.B(n_621),
.C(n_511),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_751),
.B(n_775),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_618),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_615),
.A2(n_616),
.B(n_617),
.C(n_687),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_725),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_615),
.B(n_621),
.C(n_468),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_751),
.B(n_775),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_636),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_636),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_615),
.A2(n_766),
.B(n_743),
.C(n_730),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_751),
.B(n_775),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_751),
.B(n_775),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_625),
.A2(n_518),
.B(n_476),
.Y(n_929)
);

CKINVDCx6p67_ASAP7_75t_R g930 ( 
.A(n_713),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_630),
.A2(n_746),
.B1(n_615),
.B2(n_768),
.Y(n_931)
);

AO21x1_ASAP7_75t_L g932 ( 
.A1(n_790),
.A2(n_909),
.B(n_920),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_904),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_816),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_819),
.A2(n_853),
.B(n_863),
.Y(n_936)
);

CKINVDCx11_ASAP7_75t_R g937 ( 
.A(n_930),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_837),
.A2(n_855),
.B(n_859),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_873),
.A2(n_875),
.B(n_844),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_842),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_922),
.B(n_790),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_910),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_901),
.B(n_900),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_887),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_912),
.B(n_913),
.Y(n_945)
);

OA22x2_ASAP7_75t_L g946 ( 
.A1(n_882),
.A2(n_898),
.B1(n_921),
.B2(n_860),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_794),
.Y(n_947)
);

OAI22x1_ASAP7_75t_L g948 ( 
.A1(n_827),
.A2(n_778),
.B1(n_881),
.B2(n_921),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_867),
.A2(n_845),
.B(n_878),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_918),
.B(n_923),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_916),
.A2(n_883),
.B(n_840),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_794),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_895),
.B(n_871),
.Y(n_953)
);

AO31x2_ASAP7_75t_L g954 ( 
.A1(n_780),
.A2(n_926),
.A3(n_907),
.B(n_784),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_778),
.B(n_783),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_927),
.B(n_928),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_881),
.B(n_856),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_780),
.A2(n_926),
.B(n_777),
.Y(n_958)
);

BUFx8_ASAP7_75t_L g959 ( 
.A(n_902),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_782),
.B(n_779),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_810),
.A2(n_888),
.B(n_885),
.Y(n_961)
);

AOI222xp33_ASAP7_75t_L g962 ( 
.A1(n_931),
.A2(n_903),
.B1(n_877),
.B2(n_890),
.C1(n_914),
.C2(n_823),
.Y(n_962)
);

AO31x2_ASAP7_75t_L g963 ( 
.A1(n_795),
.A2(n_789),
.A3(n_862),
.B(n_807),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_905),
.A2(n_851),
.B(n_785),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_861),
.Y(n_965)
);

AOI221xp5_ASAP7_75t_L g966 ( 
.A1(n_931),
.A2(n_890),
.B1(n_906),
.B2(n_917),
.C(n_874),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_880),
.A2(n_821),
.B(n_798),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_835),
.A2(n_787),
.B(n_806),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_812),
.A2(n_814),
.B(n_800),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_L g970 ( 
.A(n_829),
.B(n_872),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_811),
.A2(n_914),
.B1(n_868),
.B2(n_831),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_803),
.A2(n_805),
.B(n_818),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_887),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_850),
.B(n_802),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_809),
.A2(n_799),
.B(n_797),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_796),
.A2(n_865),
.B(n_893),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_818),
.A2(n_804),
.B(n_919),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_781),
.A2(n_857),
.B(n_843),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_792),
.B(n_825),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_786),
.B(n_811),
.Y(n_980)
);

OAI22x1_ASAP7_75t_L g981 ( 
.A1(n_894),
.A2(n_897),
.B1(n_858),
.B2(n_869),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_839),
.A2(n_793),
.B(n_815),
.Y(n_982)
);

OAI21xp33_ASAP7_75t_SL g983 ( 
.A1(n_894),
.A2(n_846),
.B(n_830),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_869),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_870),
.B(n_820),
.Y(n_985)
);

AO21x1_ASAP7_75t_L g986 ( 
.A1(n_896),
.A2(n_874),
.B(n_832),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_831),
.A2(n_834),
.B(n_876),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_834),
.A2(n_854),
.B(n_879),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_808),
.B(n_813),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_911),
.A2(n_828),
.B(n_864),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_828),
.A2(n_826),
.B1(n_792),
.B2(n_849),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_866),
.B(n_852),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_793),
.A2(n_861),
.B(n_847),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_858),
.A2(n_889),
.B(n_884),
.C(n_833),
.Y(n_994)
);

AND3x4_ASAP7_75t_L g995 ( 
.A(n_892),
.B(n_848),
.C(n_891),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_822),
.A2(n_824),
.B(n_817),
.Y(n_996)
);

BUFx8_ASAP7_75t_L g997 ( 
.A(n_849),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_794),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_849),
.B(n_794),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_849),
.B(n_836),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_836),
.B(n_924),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_899),
.A2(n_836),
.B(n_924),
.C(n_925),
.Y(n_1002)
);

AND2x6_ASAP7_75t_L g1003 ( 
.A(n_836),
.B(n_925),
.Y(n_1003)
);

OA22x2_ASAP7_75t_L g1004 ( 
.A1(n_848),
.A2(n_801),
.B1(n_924),
.B2(n_925),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_801),
.A2(n_924),
.B(n_925),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_861),
.A2(n_790),
.B(n_907),
.C(n_909),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_861),
.A2(n_907),
.B(n_780),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_915),
.A2(n_625),
.B(n_518),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_915),
.A2(n_625),
.B(n_518),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_790),
.A2(n_907),
.B(n_909),
.C(n_922),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_842),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_861),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_907),
.A2(n_926),
.B(n_780),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_816),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_912),
.B(n_913),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_790),
.B(n_912),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_904),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_790),
.A2(n_922),
.B(n_909),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_790),
.A2(n_907),
.B(n_909),
.C(n_922),
.Y(n_1020)
);

AOI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_790),
.A2(n_922),
.B(n_909),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_915),
.A2(n_625),
.B(n_518),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_790),
.B(n_477),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_912),
.B(n_913),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_907),
.A2(n_926),
.B(n_780),
.Y(n_1025)
);

AO31x2_ASAP7_75t_L g1026 ( 
.A1(n_780),
.A2(n_926),
.A3(n_907),
.B(n_784),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_931),
.A2(n_909),
.B1(n_907),
.B2(n_780),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_922),
.B(n_790),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_788),
.A2(n_632),
.B(n_908),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_912),
.B(n_913),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_790),
.B(n_922),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_912),
.B(n_913),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_907),
.A2(n_926),
.B(n_780),
.Y(n_1035)
);

INVx6_ASAP7_75t_SL g1036 ( 
.A(n_793),
.Y(n_1036)
);

NAND2x1_ASAP7_75t_L g1037 ( 
.A(n_794),
.B(n_642),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_790),
.A2(n_909),
.B1(n_922),
.B2(n_917),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_915),
.A2(n_625),
.B(n_518),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_816),
.Y(n_1040)
);

AO31x2_ASAP7_75t_L g1041 ( 
.A1(n_780),
.A2(n_926),
.A3(n_907),
.B(n_784),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_788),
.A2(n_632),
.B(n_908),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_887),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_915),
.A2(n_625),
.B(n_518),
.Y(n_1044)
);

OA21x2_ASAP7_75t_L g1045 ( 
.A1(n_905),
.A2(n_929),
.B(n_838),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_907),
.A2(n_926),
.B(n_780),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_907),
.A2(n_926),
.B(n_780),
.Y(n_1047)
);

AOI211x1_ASAP7_75t_L g1048 ( 
.A1(n_827),
.A2(n_922),
.B(n_928),
.C(n_927),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_1049)
);

AO21x1_ASAP7_75t_L g1050 ( 
.A1(n_790),
.A2(n_909),
.B(n_920),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_794),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_931),
.A2(n_909),
.B1(n_907),
.B2(n_780),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_887),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_907),
.A2(n_926),
.B(n_780),
.Y(n_1055)
);

O2A1O1Ixp5_ASAP7_75t_L g1056 ( 
.A1(n_907),
.A2(n_790),
.B(n_926),
.C(n_780),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_915),
.A2(n_625),
.B(n_518),
.Y(n_1057)
);

OAI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_790),
.A2(n_615),
.B(n_621),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_790),
.B(n_912),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_788),
.A2(n_632),
.B(n_908),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_841),
.A2(n_886),
.B(n_791),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_788),
.A2(n_632),
.B(n_908),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_790),
.B(n_477),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_895),
.B(n_871),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_931),
.A2(n_909),
.B1(n_907),
.B2(n_780),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_816),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_887),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_940),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_1051),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_1040),
.B(n_935),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1017),
.B(n_1060),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_974),
.B(n_1023),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_953),
.B(n_1065),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_945),
.B(n_950),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_948),
.B(n_974),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_937),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_964),
.A2(n_949),
.B(n_945),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_1014),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_953),
.B(n_1065),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1058),
.B(n_1064),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_950),
.B(n_956),
.Y(n_1082)
);

CKINVDCx11_ASAP7_75t_R g1083 ( 
.A(n_1018),
.Y(n_1083)
);

AND2x6_ASAP7_75t_L g1084 ( 
.A(n_980),
.B(n_965),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_956),
.Y(n_1085)
);

BUFx4_ASAP7_75t_SL g1086 ( 
.A(n_943),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1015),
.B(n_1024),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1015),
.B(n_1024),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1031),
.B(n_1034),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1067),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_955),
.B(n_957),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_965),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_966),
.B(n_1028),
.C(n_941),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_960),
.B(n_1048),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_942),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_933),
.B(n_1033),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_979),
.B(n_1038),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_946),
.B(n_984),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1011),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1027),
.A2(n_1066),
.B1(n_1052),
.B2(n_980),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_943),
.Y(n_1101)
);

OAI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1019),
.A2(n_1021),
.B1(n_992),
.B2(n_946),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_970),
.B(n_943),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1019),
.B(n_1021),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_944),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_981),
.B(n_1010),
.Y(n_1106)
);

O2A1O1Ixp5_ASAP7_75t_L g1107 ( 
.A1(n_986),
.A2(n_1035),
.B(n_1025),
.C(n_1046),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1036),
.Y(n_1108)
);

NAND2x1_ASAP7_75t_L g1109 ( 
.A(n_1003),
.B(n_1051),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1020),
.B(n_992),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1008),
.A2(n_1022),
.B(n_1009),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_997),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_962),
.B(n_1006),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_997),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_971),
.A2(n_1013),
.B1(n_1046),
.B2(n_1047),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1013),
.B(n_1047),
.Y(n_1116)
);

AO21x2_ASAP7_75t_L g1117 ( 
.A1(n_958),
.A2(n_1055),
.B(n_987),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_1003),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_999),
.B(n_982),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1002),
.B(n_994),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_999),
.B(n_993),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_1003),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_962),
.B(n_932),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1036),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1056),
.A2(n_971),
.B(n_991),
.C(n_983),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_954),
.B(n_1026),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1050),
.B(n_954),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_995),
.B(n_985),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_958),
.A2(n_1007),
.B1(n_985),
.B2(n_975),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_973),
.B(n_1068),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1000),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1043),
.B(n_1054),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1045),
.A2(n_978),
.B1(n_1004),
.B2(n_968),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_959),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_SL g1135 ( 
.A(n_990),
.B(n_987),
.C(n_1057),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_998),
.Y(n_1136)
);

AND2x6_ASAP7_75t_L g1137 ( 
.A(n_1012),
.B(n_952),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1039),
.A2(n_1044),
.B1(n_1004),
.B2(n_990),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_947),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_989),
.A2(n_1001),
.B1(n_996),
.B2(n_1037),
.Y(n_1140)
);

OR2x2_ASAP7_75t_SL g1141 ( 
.A(n_959),
.B(n_1041),
.Y(n_1141)
);

OR2x2_ASAP7_75t_SL g1142 ( 
.A(n_954),
.B(n_1026),
.Y(n_1142)
);

CKINVDCx14_ASAP7_75t_R g1143 ( 
.A(n_1026),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_1030),
.A2(n_1063),
.B(n_1042),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1041),
.B(n_963),
.Y(n_1145)
);

OAI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_996),
.A2(n_988),
.B(n_976),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1041),
.B(n_963),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_963),
.B(n_988),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_1005),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_977),
.B(n_961),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_967),
.A2(n_938),
.B1(n_951),
.B2(n_972),
.Y(n_1151)
);

OR2x2_ASAP7_75t_SL g1152 ( 
.A(n_1061),
.B(n_936),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_969),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_939),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1029),
.B(n_1062),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1032),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1049),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1053),
.B(n_1059),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1058),
.B(n_922),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1058),
.A2(n_907),
.B(n_926),
.C(n_780),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_953),
.B(n_1065),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1023),
.B(n_1064),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_953),
.B(n_1065),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1017),
.B(n_1060),
.Y(n_1164)
);

INVx3_ASAP7_75t_SL g1165 ( 
.A(n_935),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1014),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_953),
.B(n_1065),
.Y(n_1167)
);

O2A1O1Ixp5_ASAP7_75t_L g1168 ( 
.A1(n_986),
.A2(n_907),
.B(n_790),
.C(n_922),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1017),
.B(n_1060),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_SL g1170 ( 
.A(n_1058),
.B(n_726),
.Y(n_1170)
);

CKINVDCx6p67_ASAP7_75t_R g1171 ( 
.A(n_937),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1058),
.B(n_922),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1040),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1023),
.B(n_1064),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_953),
.B(n_1065),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1017),
.B(n_1060),
.Y(n_1176)
);

NAND2x1p5_ASAP7_75t_L g1177 ( 
.A(n_1040),
.B(n_935),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_940),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1058),
.A2(n_907),
.B(n_926),
.C(n_780),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1017),
.B(n_1060),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_986),
.A2(n_907),
.B(n_790),
.C(n_922),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_940),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1023),
.B(n_1064),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_964),
.A2(n_949),
.B(n_625),
.Y(n_1184)
);

O2A1O1Ixp5_ASAP7_75t_SL g1185 ( 
.A1(n_1013),
.A2(n_1035),
.B(n_1046),
.C(n_1025),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1023),
.B(n_1064),
.Y(n_1186)
);

BUFx12f_ASAP7_75t_L g1187 ( 
.A(n_937),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_953),
.B(n_1065),
.Y(n_1188)
);

INVx5_ASAP7_75t_L g1189 ( 
.A(n_1003),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_974),
.B(n_904),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1058),
.A2(n_790),
.B1(n_909),
.B2(n_922),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1017),
.A2(n_922),
.B1(n_909),
.B2(n_668),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1040),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1017),
.A2(n_909),
.B1(n_790),
.B2(n_907),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_937),
.Y(n_1195)
);

OAI21xp33_ASAP7_75t_L g1196 ( 
.A1(n_1058),
.A2(n_790),
.B(n_615),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_940),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1058),
.A2(n_922),
.B(n_790),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1058),
.A2(n_790),
.B(n_907),
.C(n_909),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_964),
.A2(n_949),
.B(n_625),
.Y(n_1200)
);

AO21x1_ASAP7_75t_SL g1201 ( 
.A1(n_1113),
.A2(n_1123),
.B(n_1104),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1195),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1093),
.A2(n_1196),
.B1(n_1172),
.B2(n_1159),
.Y(n_1203)
);

AO21x1_ASAP7_75t_SL g1204 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1145),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1126),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1182),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1110),
.B(n_1116),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1069),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1093),
.A2(n_1196),
.B1(n_1115),
.B2(n_1192),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1075),
.B(n_1082),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1194),
.A2(n_1128),
.B1(n_1191),
.B2(n_1106),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1095),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1142),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1103),
.B(n_1120),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1100),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1100),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1099),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1191),
.A2(n_1081),
.B1(n_1076),
.B2(n_1186),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1173),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1178),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1120),
.B(n_1189),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1103),
.B(n_1098),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1071),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1171),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1177),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1170),
.A2(n_1176),
.B1(n_1180),
.B2(n_1072),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1199),
.A2(n_1168),
.B(n_1181),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1084),
.Y(n_1228)
);

BUFx8_ASAP7_75t_L g1229 ( 
.A(n_1187),
.Y(n_1229)
);

NAND2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1189),
.B(n_1076),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1197),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1107),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1155),
.A2(n_1200),
.B(n_1184),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1085),
.B(n_1143),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1166),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1189),
.B(n_1129),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1087),
.B(n_1088),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1090),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1079),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1083),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1132),
.Y(n_1241)
);

CKINVDCx6p67_ASAP7_75t_R g1242 ( 
.A(n_1165),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1077),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1089),
.B(n_1198),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1105),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1174),
.A2(n_1183),
.B1(n_1162),
.B2(n_1117),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1101),
.A2(n_1097),
.B1(n_1164),
.B2(n_1169),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1130),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1096),
.Y(n_1249)
);

AO21x1_ASAP7_75t_L g1250 ( 
.A1(n_1160),
.A2(n_1179),
.B(n_1125),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1073),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1193),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1131),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1094),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1136),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1129),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1074),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1119),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1091),
.B(n_1185),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1101),
.A2(n_1138),
.B1(n_1117),
.B2(n_1112),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1190),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1119),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1119),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1118),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1084),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1080),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1080),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1148),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1102),
.A2(n_1133),
.B1(n_1188),
.B2(n_1175),
.Y(n_1269)
);

AO21x1_ASAP7_75t_SL g1270 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_1156),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1161),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1161),
.A2(n_1167),
.B1(n_1163),
.B2(n_1175),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1153),
.B(n_1149),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1152),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

BUFx2_ASAP7_75t_R g1276 ( 
.A(n_1134),
.Y(n_1276)
);

BUFx2_ASAP7_75t_R g1277 ( 
.A(n_1114),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1135),
.A2(n_1151),
.B(n_1078),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1121),
.B(n_1084),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1163),
.A2(n_1188),
.B1(n_1167),
.B2(n_1141),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1109),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1137),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1139),
.Y(n_1283)
);

AO21x2_ASAP7_75t_L g1284 ( 
.A1(n_1146),
.A2(n_1157),
.B(n_1158),
.Y(n_1284)
);

AOI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1150),
.A2(n_1140),
.B(n_1154),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1150),
.A2(n_1144),
.B(n_1124),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1108),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1070),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1092),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1092),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1092),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1137),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1086),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1093),
.B(n_922),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1173),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1182),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1170),
.A2(n_922),
.B1(n_674),
.B2(n_790),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1075),
.A2(n_790),
.B1(n_909),
.B2(n_922),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1166),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1170),
.A2(n_922),
.B1(n_674),
.B2(n_790),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1195),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1173),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1111),
.A2(n_1016),
.B(n_934),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1173),
.Y(n_1304)
);

INVx6_ASAP7_75t_L g1305 ( 
.A(n_1122),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1126),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1075),
.B(n_790),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1207),
.B(n_1259),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1236),
.B(n_1258),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1294),
.A2(n_1297),
.B1(n_1300),
.B2(n_1209),
.Y(n_1310)
);

AO21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1227),
.A2(n_1232),
.B(n_1213),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1235),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1299),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1268),
.B(n_1213),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1238),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1205),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1239),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1233),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1226),
.B(n_1210),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1221),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1240),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1237),
.B(n_1244),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1306),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1207),
.B(n_1259),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1261),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1251),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1256),
.B(n_1201),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1219),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1298),
.A2(n_1203),
.B(n_1307),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1211),
.A2(n_1218),
.B(n_1247),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1256),
.B(n_1201),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1275),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1253),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1232),
.B(n_1215),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1248),
.B(n_1254),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1219),
.Y(n_1337)
);

INVxp33_ASAP7_75t_L g1338 ( 
.A(n_1257),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1236),
.B(n_1258),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1262),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1275),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1303),
.A2(n_1285),
.B(n_1286),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1234),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1234),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1262),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1263),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1250),
.A2(n_1278),
.B(n_1221),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1274),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1278),
.A2(n_1250),
.B(n_1284),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1274),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1216),
.B(n_1204),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1273),
.A2(n_1230),
.B(n_1281),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1246),
.B(n_1278),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1221),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1282),
.B(n_1279),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1204),
.B(n_1231),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1295),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1222),
.B(n_1214),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1208),
.A2(n_1217),
.B(n_1220),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1222),
.B(n_1214),
.Y(n_1360)
);

OAI21xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1279),
.A2(n_1212),
.B(n_1296),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1255),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1230),
.A2(n_1281),
.B(n_1269),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1206),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1295),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1230),
.A2(n_1260),
.B(n_1252),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1245),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1241),
.B(n_1214),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1228),
.A2(n_1265),
.B(n_1270),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1265),
.A2(n_1270),
.B(n_1288),
.Y(n_1370)
);

NAND2xp33_ASAP7_75t_R g1371 ( 
.A(n_1293),
.B(n_1222),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1240),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1302),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1302),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1202),
.Y(n_1375)
);

NOR2x1_ASAP7_75t_L g1376 ( 
.A(n_1329),
.B(n_1281),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1335),
.B(n_1280),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1308),
.B(n_1264),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1308),
.B(n_1324),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1324),
.B(n_1264),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1349),
.B(n_1264),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1349),
.B(n_1290),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1370),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1351),
.B(n_1290),
.Y(n_1384)
);

CKINVDCx14_ASAP7_75t_R g1385 ( 
.A(n_1372),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1349),
.B(n_1291),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1370),
.B(n_1291),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1370),
.B(n_1289),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1316),
.Y(n_1389)
);

NAND2x1_ASAP7_75t_L g1390 ( 
.A(n_1309),
.B(n_1305),
.Y(n_1390)
);

OR2x6_ASAP7_75t_L g1391 ( 
.A(n_1309),
.B(n_1339),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1332),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1369),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1353),
.B(n_1304),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1369),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1310),
.A2(n_1271),
.B1(n_1266),
.B2(n_1267),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1322),
.B(n_1304),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1347),
.A2(n_1283),
.B(n_1272),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1353),
.B(n_1292),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1359),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1311),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1369),
.Y(n_1402)
);

INVxp67_ASAP7_75t_SL g1403 ( 
.A(n_1394),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1376),
.B(n_1330),
.C(n_1319),
.Y(n_1404)
);

OAI211xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1376),
.A2(n_1334),
.B(n_1315),
.C(n_1317),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1376),
.B(n_1366),
.C(n_1396),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1397),
.B(n_1333),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1397),
.B(n_1325),
.Y(n_1408)
);

AND2x2_ASAP7_75t_SL g1409 ( 
.A(n_1383),
.B(n_1369),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1379),
.B(n_1326),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1396),
.A2(n_1277),
.B1(n_1368),
.B2(n_1365),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1385),
.A2(n_1328),
.B1(n_1337),
.B2(n_1357),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1394),
.B(n_1362),
.C(n_1336),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1385),
.A2(n_1331),
.B1(n_1327),
.B2(n_1371),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1394),
.B(n_1313),
.C(n_1312),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1377),
.A2(n_1361),
.B1(n_1399),
.B2(n_1327),
.C(n_1331),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1401),
.A2(n_1355),
.B(n_1360),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1379),
.B(n_1348),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1379),
.B(n_1351),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1379),
.B(n_1348),
.Y(n_1420)
);

AND2x2_ASAP7_75t_SL g1421 ( 
.A(n_1383),
.B(n_1320),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1401),
.A2(n_1355),
.B(n_1360),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1378),
.B(n_1350),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1398),
.A2(n_1358),
.B1(n_1309),
.B2(n_1339),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1388),
.B(n_1356),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1382),
.B(n_1350),
.C(n_1361),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1388),
.B(n_1356),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1378),
.B(n_1343),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1390),
.A2(n_1363),
.B(n_1352),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1377),
.B(n_1320),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1388),
.B(n_1311),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1388),
.B(n_1309),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1378),
.B(n_1344),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1387),
.B(n_1339),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1382),
.B(n_1346),
.C(n_1345),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1398),
.A2(n_1358),
.B1(n_1339),
.B2(n_1354),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1400),
.A2(n_1342),
.B(n_1318),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1387),
.B(n_1380),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1392),
.B(n_1341),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1399),
.B(n_1314),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_R g1442 ( 
.A(n_1384),
.B(n_1321),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1392),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1389),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1382),
.B(n_1346),
.C(n_1345),
.Y(n_1445)
);

OAI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1390),
.A2(n_1374),
.B1(n_1373),
.B2(n_1375),
.C(n_1355),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1387),
.B(n_1340),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1381),
.A2(n_1338),
.B1(n_1364),
.B2(n_1367),
.C(n_1323),
.Y(n_1448)
);

NOR3xp33_ASAP7_75t_L g1449 ( 
.A(n_1390),
.B(n_1363),
.C(n_1287),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1444),
.B(n_1382),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1444),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1439),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1426),
.B(n_1393),
.Y(n_1453)
);

INVxp33_ASAP7_75t_L g1454 ( 
.A(n_1412),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1404),
.B(n_1364),
.C(n_1367),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1441),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1426),
.B(n_1428),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1443),
.B(n_1386),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1409),
.B(n_1419),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1433),
.B(n_1393),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1441),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1447),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1407),
.B(n_1386),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1409),
.B(n_1393),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1408),
.B(n_1242),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1403),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1413),
.B(n_1386),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1409),
.B(n_1419),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1438),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1436),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1445),
.Y(n_1471)
);

AND2x4_ASAP7_75t_SL g1472 ( 
.A(n_1449),
.B(n_1391),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1421),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1435),
.B(n_1395),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1432),
.B(n_1421),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1422),
.B(n_1399),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1410),
.B(n_1383),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1429),
.B(n_1395),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1438),
.Y(n_1479)
);

AND2x4_ASAP7_75t_SL g1480 ( 
.A(n_1414),
.B(n_1391),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1418),
.B(n_1391),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1420),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1434),
.B(n_1402),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1425),
.B(n_1391),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1437),
.B(n_1402),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1454),
.A2(n_1406),
.B(n_1415),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1482),
.B(n_1415),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1470),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1465),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1459),
.B(n_1468),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1459),
.B(n_1468),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1461),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1474),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1482),
.B(n_1413),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1463),
.B(n_1424),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1473),
.B(n_1402),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1451),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1455),
.B(n_1430),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1451),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1470),
.B(n_1405),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1471),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1461),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1456),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1463),
.B(n_1431),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1456),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1455),
.B(n_1471),
.C(n_1448),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1474),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1469),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1466),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1467),
.B(n_1440),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1452),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1467),
.B(n_1384),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1452),
.Y(n_1515)
);

NOR2x1p5_ASAP7_75t_SL g1516 ( 
.A(n_1469),
.B(n_1400),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1450),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1469),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1457),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1457),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1457),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1477),
.B(n_1427),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1462),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1462),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1500),
.B(n_1481),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1508),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1492),
.B(n_1473),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1490),
.B(n_1459),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1497),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1490),
.B(n_1480),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1499),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1511),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1503),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1491),
.B(n_1468),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1505),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1513),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_1489),
.Y(n_1537)
);

NOR2x1p5_ASAP7_75t_SL g1538 ( 
.A(n_1508),
.B(n_1479),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1500),
.Y(n_1539)
);

OR2x2_ASAP7_75t_SL g1540 ( 
.A(n_1506),
.B(n_1442),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1515),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1486),
.A2(n_1414),
.B(n_1485),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1523),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1522),
.B(n_1450),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1491),
.B(n_1475),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1458),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1518),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1488),
.B(n_1501),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1524),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1502),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1510),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1518),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1510),
.B(n_1481),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1487),
.B(n_1478),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1493),
.B(n_1475),
.Y(n_1555)
);

NOR2x1_ASAP7_75t_L g1556 ( 
.A(n_1489),
.B(n_1224),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1494),
.B(n_1478),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1504),
.B(n_1483),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1498),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1509),
.B(n_1458),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1519),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1520),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_L g1564 ( 
.A(n_1498),
.B(n_1416),
.C(n_1411),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1493),
.B(n_1475),
.Y(n_1565)
);

INVxp67_ASAP7_75t_SL g1566 ( 
.A(n_1496),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1521),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1529),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1537),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1551),
.B(n_1514),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1545),
.B(n_1507),
.Y(n_1571)
);

NOR2x1_ASAP7_75t_L g1572 ( 
.A(n_1556),
.B(n_1498),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1545),
.B(n_1507),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1539),
.B(n_1229),
.Y(n_1574)
);

NAND3x1_ASAP7_75t_L g1575 ( 
.A(n_1542),
.B(n_1464),
.C(n_1229),
.Y(n_1575)
);

AOI21xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1564),
.A2(n_1498),
.B(n_1496),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1528),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1525),
.B(n_1495),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1529),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1480),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1559),
.A2(n_1480),
.B1(n_1472),
.B2(n_1484),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1540),
.Y(n_1582)
);

NOR2x1_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1224),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1536),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1517),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1550),
.B(n_1554),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1534),
.B(n_1464),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1546),
.B(n_1517),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1555),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1558),
.B(n_1453),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1536),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1530),
.B(n_1464),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1527),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1541),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1530),
.B(n_1472),
.Y(n_1596)
);

AND2x2_ASAP7_75t_SL g1597 ( 
.A(n_1540),
.B(n_1472),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1546),
.B(n_1544),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1527),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1527),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1541),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1555),
.B(n_1460),
.Y(n_1602)
);

AO21x2_ASAP7_75t_L g1603 ( 
.A1(n_1526),
.A2(n_1479),
.B(n_1485),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1582),
.A2(n_1532),
.B1(n_1566),
.B2(n_1567),
.C(n_1533),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1582),
.A2(n_1530),
.B1(n_1565),
.B2(n_1484),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1572),
.A2(n_1535),
.B(n_1533),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1572),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1568),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1568),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1569),
.B(n_1565),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1569),
.B(n_1531),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1569),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

AND3x1_ASAP7_75t_L g1614 ( 
.A(n_1583),
.B(n_1485),
.C(n_1535),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1579),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1576),
.A2(n_1544),
.B(n_1567),
.C(n_1562),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1583),
.A2(n_1538),
.B(n_1293),
.C(n_1516),
.Y(n_1617)
);

AOI21xp33_ASAP7_75t_L g1618 ( 
.A1(n_1597),
.A2(n_1543),
.B(n_1562),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1584),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1597),
.B(n_1563),
.Y(n_1621)
);

AOI21xp33_ASAP7_75t_L g1622 ( 
.A1(n_1600),
.A2(n_1543),
.B(n_1563),
.Y(n_1622)
);

OAI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1586),
.A2(n_1560),
.B(n_1538),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1575),
.A2(n_1549),
.B1(n_1417),
.B2(n_1423),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1584),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

NOR2xp67_ASAP7_75t_L g1628 ( 
.A(n_1594),
.B(n_1561),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1571),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1610),
.B(n_1596),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1628),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1612),
.B(n_1578),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1610),
.B(n_1596),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1619),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1629),
.B(n_1596),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1608),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1608),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1607),
.B(n_1577),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1629),
.B(n_1621),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1626),
.B(n_1598),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1619),
.B(n_1577),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1611),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1609),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1621),
.B(n_1614),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1606),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1618),
.B(n_1574),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1604),
.B(n_1616),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1627),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1648),
.A2(n_1617),
.B(n_1622),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1646),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1645),
.B(n_1617),
.C(n_1623),
.Y(n_1652)
);

AOI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1631),
.A2(n_1644),
.B(n_1647),
.C(n_1642),
.Y(n_1653)
);

AOI211xp5_ASAP7_75t_L g1654 ( 
.A1(n_1644),
.A2(n_1625),
.B(n_1620),
.C(n_1615),
.Y(n_1654)
);

AO21x1_ASAP7_75t_L g1655 ( 
.A1(n_1636),
.A2(n_1627),
.B(n_1613),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1642),
.A2(n_1599),
.B1(n_1605),
.B2(n_1592),
.C(n_1601),
.Y(n_1656)
);

AOI322xp5_ASAP7_75t_L g1657 ( 
.A1(n_1634),
.A2(n_1585),
.A3(n_1588),
.B1(n_1570),
.B2(n_1599),
.C1(n_1624),
.C2(n_1571),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1639),
.B(n_1573),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1639),
.B(n_1573),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_SL g1660 ( 
.A1(n_1634),
.A2(n_1243),
.B(n_1202),
.C(n_1301),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1632),
.A2(n_1598),
.B(n_1595),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1651),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1653),
.B(n_1638),
.C(n_1641),
.Y(n_1663)
);

NAND4xp75_ASAP7_75t_L g1664 ( 
.A(n_1655),
.B(n_1635),
.C(n_1630),
.D(n_1633),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1652),
.A2(n_1640),
.B(n_1633),
.Y(n_1665)
);

OAI322xp33_ASAP7_75t_L g1666 ( 
.A1(n_1650),
.A2(n_1649),
.A3(n_1643),
.B1(n_1637),
.B2(n_1636),
.C1(n_1646),
.C2(n_1640),
.Y(n_1666)
);

NAND2x1p5_ASAP7_75t_SL g1667 ( 
.A(n_1660),
.B(n_1630),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1658),
.B(n_1635),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1659),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1654),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1661),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1665),
.B(n_1657),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1662),
.Y(n_1673)
);

NOR3xp33_ASAP7_75t_SL g1674 ( 
.A(n_1666),
.B(n_1656),
.C(n_1643),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_L g1675 ( 
.A(n_1663),
.B(n_1666),
.C(n_1670),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_L g1676 ( 
.A(n_1671),
.B(n_1649),
.C(n_1637),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1675),
.A2(n_1664),
.B1(n_1668),
.B2(n_1669),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1674),
.B(n_1667),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1676),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1673),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1672),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1675),
.A2(n_1575),
.B1(n_1595),
.B2(n_1601),
.Y(n_1682)
);

NAND4xp75_ASAP7_75t_L g1683 ( 
.A(n_1678),
.B(n_1229),
.C(n_1646),
.D(n_1587),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1679),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1677),
.B(n_1646),
.C(n_1287),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1682),
.B(n_1593),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1680),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1686),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1683),
.B(n_1681),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1685),
.A2(n_1593),
.B1(n_1580),
.B2(n_1602),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1688),
.Y(n_1691)
);

XOR2xp5_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1684),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1687),
.B(n_1689),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1692),
.A2(n_1243),
.B1(n_1301),
.B2(n_1242),
.Y(n_1694)
);

NAND3x2_ASAP7_75t_L g1695 ( 
.A(n_1694),
.B(n_1690),
.C(n_1589),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1693),
.B(n_1589),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1603),
.B(n_1593),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_L g1698 ( 
.A(n_1695),
.B(n_1581),
.C(n_1547),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1698),
.A2(n_1697),
.B(n_1276),
.Y(n_1699)
);

AOI322xp5_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1580),
.A3(n_1587),
.B1(n_1602),
.B2(n_1547),
.C1(n_1552),
.C2(n_1526),
.Y(n_1700)
);

OAI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1225),
.B1(n_1223),
.B2(n_1552),
.C(n_1591),
.Y(n_1701)
);

AOI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1223),
.B(n_1225),
.C(n_1580),
.Y(n_1702)
);


endmodule