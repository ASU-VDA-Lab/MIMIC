module real_aes_15427_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g106 ( .A(n_0), .B(n_107), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_1), .A2(n_4), .B1(n_267), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_2), .A2(n_43), .B1(n_148), .B2(n_240), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_3), .A2(n_22), .B1(n_208), .B2(n_240), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_5), .A2(n_15), .B1(n_180), .B2(n_182), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_6), .A2(n_61), .B1(n_144), .B2(n_210), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_7), .A2(n_16), .B1(n_148), .B2(n_153), .Y(n_499) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_9), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_10), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_11), .A2(n_17), .B1(n_143), .B2(n_147), .Y(n_142) );
OR2x2_ASAP7_75t_L g114 ( .A(n_12), .B(n_38), .Y(n_114) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_14), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_18), .A2(n_98), .B1(n_180), .B2(n_267), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_19), .A2(n_39), .B1(n_172), .B2(n_174), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_20), .B(n_181), .Y(n_229) );
OAI21x1_ASAP7_75t_L g159 ( .A1(n_21), .A2(n_58), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_23), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_24), .A2(n_54), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_24), .Y(n_132) );
INVx4_ASAP7_75t_R g524 ( .A(n_25), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_26), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_27), .B(n_151), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_28), .A2(n_47), .B1(n_193), .B2(n_196), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_29), .A2(n_53), .B1(n_180), .B2(n_196), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_30), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_31), .B(n_172), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_32), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_33), .B(n_240), .Y(n_567) );
INVx1_ASAP7_75t_L g606 ( .A(n_34), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_SL g542 ( .A1(n_35), .A2(n_148), .B(n_150), .C(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_36), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_37), .A2(n_55), .B1(n_148), .B2(n_196), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_40), .A2(n_86), .B1(n_148), .B2(n_207), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_41), .A2(n_79), .B1(n_815), .B2(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_41), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_42), .A2(n_46), .B1(n_148), .B2(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_44), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_45), .A2(n_60), .B1(n_180), .B2(n_194), .Y(n_269) );
INVx1_ASAP7_75t_L g564 ( .A(n_48), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_49), .B(n_148), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_50), .Y(n_583) );
INVx2_ASAP7_75t_L g483 ( .A(n_51), .Y(n_483) );
INVx1_ASAP7_75t_L g112 ( .A(n_52), .Y(n_112) );
BUFx3_ASAP7_75t_L g824 ( .A(n_52), .Y(n_824) );
INVx1_ASAP7_75t_L g133 ( .A(n_54), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_56), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_57), .A2(n_87), .B1(n_148), .B2(n_196), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_59), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_62), .A2(n_74), .B1(n_193), .B2(n_194), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_63), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_64), .A2(n_76), .B1(n_148), .B2(n_153), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_65), .A2(n_97), .B1(n_147), .B2(n_180), .Y(n_216) );
INVx1_ASAP7_75t_L g160 ( .A(n_66), .Y(n_160) );
AND2x4_ASAP7_75t_L g162 ( .A(n_67), .B(n_163), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_68), .A2(n_89), .B1(n_193), .B2(n_196), .Y(n_602) );
AO22x1_ASAP7_75t_L g511 ( .A1(n_69), .A2(n_75), .B1(n_174), .B2(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g163 ( .A(n_70), .Y(n_163) );
AND2x2_ASAP7_75t_L g545 ( .A(n_71), .B(n_235), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_72), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_73), .B(n_210), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_77), .B(n_240), .Y(n_584) );
INVx2_ASAP7_75t_L g151 ( .A(n_78), .Y(n_151) );
INVx1_ASAP7_75t_L g816 ( .A(n_79), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_80), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_81), .B(n_235), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_82), .A2(n_96), .B1(n_196), .B2(n_210), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_83), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_84), .B(n_158), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_85), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_88), .B(n_235), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_90), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_91), .B(n_235), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_92), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
NAND2xp33_ASAP7_75t_L g232 ( .A(n_93), .B(n_181), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_94), .A2(n_155), .B(n_210), .C(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g526 ( .A(n_95), .B(n_527), .Y(n_526) );
NAND2xp33_ASAP7_75t_L g588 ( .A(n_99), .B(n_173), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_115), .B(n_833), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx2_ASAP7_75t_SL g842 ( .A(n_106), .Y(n_842) );
INVx5_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx8_ASAP7_75t_R g121 ( .A(n_109), .Y(n_121) );
INVx3_ASAP7_75t_L g843 ( .A(n_109), .Y(n_843) );
AND2x6_ASAP7_75t_SL g109 ( .A(n_110), .B(n_113), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_112), .Y(n_127) );
AND3x2_ASAP7_75t_L g126 ( .A(n_113), .B(n_127), .C(n_128), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_113), .B(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2x1_ASAP7_75t_L g832 ( .A(n_114), .B(n_824), .Y(n_832) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_479), .B(n_484), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_117), .A2(n_132), .B1(n_834), .B2(n_844), .Y(n_833) );
NOR2x1_ASAP7_75t_L g117 ( .A(n_118), .B(n_123), .Y(n_117) );
NOR2x1_ASAP7_75t_SL g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_130), .Y(n_123) );
BUFx2_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g812 ( .A(n_129), .Y(n_812) );
XNOR2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_134), .Y(n_130) );
NAND4xp25_ASAP7_75t_L g134 ( .A(n_135), .B(n_354), .C(n_408), .D(n_447), .Y(n_134) );
NAND4xp75_ASAP7_75t_L g813 ( .A(n_135), .B(n_354), .C(n_408), .D(n_447), .Y(n_813) );
NOR2x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_312), .Y(n_135) );
NAND3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_255), .C(n_294), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_202), .B1(n_245), .B2(n_250), .Y(n_137) );
INVx1_ASAP7_75t_L g418 ( .A(n_138), .Y(n_418) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_167), .Y(n_138) );
INVx1_ASAP7_75t_L g281 ( .A(n_139), .Y(n_281) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx4_ASAP7_75t_SL g247 ( .A(n_140), .Y(n_247) );
AND2x2_ASAP7_75t_L g299 ( .A(n_140), .B(n_188), .Y(n_299) );
AND2x2_ASAP7_75t_L g338 ( .A(n_140), .B(n_169), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_140), .B(n_275), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_140), .B(n_474), .Y(n_473) );
AO31x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_156), .A3(n_161), .B(n_164), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_149), .B1(n_152), .B2(n_154), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_145), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_146), .Y(n_148) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_146), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_146), .Y(n_183) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
INVx2_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_146), .Y(n_240) );
INVx1_ASAP7_75t_L g268 ( .A(n_146), .Y(n_268) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g153 ( .A(n_148), .Y(n_153) );
INVx1_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_149), .A2(n_171), .B1(n_176), .B2(n_179), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_149), .A2(n_176), .B1(n_192), .B2(n_195), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_149), .A2(n_206), .B1(n_209), .B2(n_211), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_149), .A2(n_154), .B1(n_216), .B2(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_149), .A2(n_231), .B(n_232), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_149), .A2(n_176), .B1(n_239), .B2(n_241), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_149), .A2(n_176), .B1(n_266), .B2(n_269), .Y(n_265) );
OAI22x1_ASAP7_75t_L g498 ( .A1(n_149), .A2(n_211), .B1(n_499), .B2(n_500), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_149), .A2(n_507), .B1(n_550), .B2(n_551), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_149), .A2(n_211), .B1(n_602), .B2(n_603), .Y(n_601) );
INVx6_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
O2A1O1Ixp5_ASAP7_75t_L g227 ( .A1(n_150), .A2(n_153), .B(n_228), .C(n_229), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_150), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_150), .A2(n_588), .B(n_589), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_150), .A2(n_506), .B(n_511), .C(n_514), .Y(n_627) );
BUFx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g155 ( .A(n_151), .Y(n_155) );
INVx2_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
INVx1_ASAP7_75t_L g541 ( .A(n_151), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g582 ( .A1(n_153), .A2(n_583), .B(n_584), .C(n_585), .Y(n_582) );
INVx1_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_156), .A2(n_215), .A3(n_218), .B(n_220), .Y(n_214) );
AOI21x1_ASAP7_75t_L g533 ( .A1(n_156), .A2(n_534), .B(n_545), .Y(n_533) );
AO31x2_ASAP7_75t_L g600 ( .A1(n_156), .A2(n_197), .A3(n_601), .B(n_605), .Y(n_600) );
BUFx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_157), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g527 ( .A(n_157), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_157), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_157), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
INVx2_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
OAI21xp33_ASAP7_75t_L g514 ( .A1(n_158), .A2(n_509), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
AO31x2_ASAP7_75t_L g169 ( .A1(n_161), .A2(n_170), .A3(n_184), .B(n_186), .Y(n_169) );
INVx2_ASAP7_75t_L g219 ( .A(n_161), .Y(n_219) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_161), .A2(n_238), .A3(n_242), .B(n_243), .Y(n_237) );
AO31x2_ASAP7_75t_L g497 ( .A1(n_161), .A2(n_201), .A3(n_498), .B(n_501), .Y(n_497) );
BUFx10_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
INVx1_ASAP7_75t_L g515 ( .A(n_162), .Y(n_515) );
BUFx10_ASAP7_75t_L g552 ( .A(n_162), .Y(n_552) );
NOR2xp33_ASAP7_75t_SL g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx2_ASAP7_75t_L g190 ( .A(n_165), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_165), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g322 ( .A(n_168), .B(n_297), .Y(n_322) );
OR2x2_ASAP7_75t_L g364 ( .A(n_168), .B(n_344), .Y(n_364) );
OR2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_188), .Y(n_168) );
INVx2_ASAP7_75t_L g249 ( .A(n_169), .Y(n_249) );
INVx1_ASAP7_75t_L g275 ( .A(n_169), .Y(n_275) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_169), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_169), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g429 ( .A(n_169), .Y(n_429) );
AND2x2_ASAP7_75t_L g434 ( .A(n_169), .B(n_263), .Y(n_434) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g193 ( .A(n_173), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g523 ( .A1(n_173), .A2(n_183), .B1(n_524), .B2(n_525), .Y(n_523) );
OAI21xp33_ASAP7_75t_SL g560 ( .A1(n_174), .A2(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g507 ( .A(n_177), .Y(n_507) );
BUFx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g586 ( .A(n_178), .Y(n_586) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_181), .Y(n_512) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_184), .A2(n_197), .A3(n_205), .B(n_212), .Y(n_204) );
BUFx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_185), .B(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_185), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_SL g225 ( .A(n_185), .Y(n_225) );
INVx4_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_185), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g568 ( .A(n_185), .B(n_552), .Y(n_568) );
AND2x4_ASAP7_75t_L g248 ( .A(n_188), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g272 ( .A(n_188), .Y(n_272) );
INVx2_ASAP7_75t_L g321 ( .A(n_188), .Y(n_321) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_188), .Y(n_337) );
INVx1_ASAP7_75t_L g474 ( .A(n_188), .Y(n_474) );
AO31x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_191), .A3(n_197), .B(n_199), .Y(n_188) );
AO31x2_ASAP7_75t_L g264 ( .A1(n_189), .A2(n_218), .A3(n_265), .B(n_270), .Y(n_264) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_189), .A2(n_518), .B(n_526), .Y(n_517) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_196), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g604 ( .A(n_196), .Y(n_604) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_SL g233 ( .A(n_198), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_201), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_222), .Y(n_202) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_203), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_203), .B(n_305), .Y(n_309) );
AND2x2_ASAP7_75t_L g366 ( .A(n_203), .B(n_353), .Y(n_366) );
AND2x4_ASAP7_75t_SL g475 ( .A(n_203), .B(n_277), .Y(n_475) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
BUFx2_ASAP7_75t_L g256 ( .A(n_204), .Y(n_256) );
OR2x2_ASAP7_75t_L g293 ( .A(n_204), .B(n_279), .Y(n_293) );
AND2x4_ASAP7_75t_L g306 ( .A(n_204), .B(n_254), .Y(n_306) );
INVx2_ASAP7_75t_L g334 ( .A(n_204), .Y(n_334) );
OR2x2_ASAP7_75t_L g360 ( .A(n_204), .B(n_237), .Y(n_360) );
INVx1_ASAP7_75t_L g413 ( .A(n_204), .Y(n_413) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_208), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_211), .B(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g254 ( .A(n_214), .Y(n_254) );
BUFx2_ASAP7_75t_L g332 ( .A(n_214), .Y(n_332) );
AND2x2_ASAP7_75t_L g420 ( .A(n_214), .B(n_334), .Y(n_420) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_219), .A2(n_519), .B(n_522), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_222), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
AND2x4_ASAP7_75t_L g333 ( .A(n_223), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g407 ( .A(n_223), .B(n_254), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_223), .B(n_256), .Y(n_425) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
BUFx2_ASAP7_75t_L g358 ( .A(n_224), .Y(n_358) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_234), .Y(n_224) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_225), .A2(n_226), .B(n_234), .Y(n_260) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_230), .B(n_233), .Y(n_226) );
INVx2_ASAP7_75t_L g242 ( .A(n_235), .Y(n_242) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_235), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_236), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_237), .Y(n_292) );
INVx1_ASAP7_75t_L g328 ( .A(n_237), .Y(n_328) );
AND2x2_ASAP7_75t_L g353 ( .A(n_237), .B(n_260), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_240), .B(n_537), .Y(n_536) );
AO31x2_ASAP7_75t_L g548 ( .A1(n_242), .A2(n_549), .A3(n_552), .B(n_553), .Y(n_548) );
AND2x2_ASAP7_75t_L g445 ( .A(n_245), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g478 ( .A(n_245), .B(n_343), .Y(n_478) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
INVx1_ASAP7_75t_L g441 ( .A(n_246), .Y(n_441) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g273 ( .A(n_247), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g308 ( .A(n_247), .B(n_263), .Y(n_308) );
INVx1_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
INVx2_ASAP7_75t_L g350 ( .A(n_247), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_247), .B(n_272), .Y(n_363) );
OR2x2_ASAP7_75t_L g372 ( .A(n_247), .B(n_326), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_247), .B(n_320), .Y(n_382) );
AND2x2_ASAP7_75t_L g451 ( .A(n_247), .B(n_429), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_248), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g307 ( .A(n_248), .B(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_248), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_248), .B(n_284), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_248), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g463 ( .A(n_248), .B(n_349), .Y(n_463) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_251), .A2(n_317), .B1(n_401), .B2(n_402), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_252), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g457 ( .A(n_253), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g477 ( .A(n_253), .B(n_353), .Y(n_477) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g289 ( .A(n_254), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_254), .B(n_278), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_254), .B(n_416), .Y(n_415) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_254), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B1(n_283), .B2(n_287), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_256), .B(n_258), .Y(n_345) );
NAND2x1_ASAP7_75t_L g406 ( .A(n_256), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g460 ( .A(n_256), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B1(n_276), .B2(n_280), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_259), .Y(n_416) );
INVx1_ASAP7_75t_L g458 ( .A(n_259), .Y(n_458) );
INVx1_ASAP7_75t_L g279 ( .A(n_260), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_273), .Y(n_261) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_262), .A2(n_347), .B(n_351), .C(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g384 ( .A(n_262), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_262), .B(n_338), .Y(n_422) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_272), .Y(n_262) );
INVx3_ASAP7_75t_L g344 ( .A(n_263), .Y(n_344) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g282 ( .A(n_264), .B(n_272), .Y(n_282) );
INVx2_ASAP7_75t_L g286 ( .A(n_264), .Y(n_286) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_268), .B(n_539), .Y(n_538) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_273), .B(n_343), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_273), .B(n_336), .Y(n_375) );
INVx1_ASAP7_75t_L g404 ( .A(n_273), .Y(n_404) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_276), .A2(n_462), .B(n_465), .Y(n_461) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_277), .A2(n_296), .B(n_300), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_277), .B(n_431), .Y(n_467) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx3_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
AND2x4_ASAP7_75t_L g444 ( .A(n_282), .B(n_311), .Y(n_444) );
AND2x2_ASAP7_75t_L g450 ( .A(n_282), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g381 ( .A(n_284), .Y(n_381) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g301 ( .A(n_285), .B(n_292), .Y(n_301) );
AND2x2_ASAP7_75t_L g427 ( .A(n_285), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g298 ( .A(n_286), .Y(n_298) );
OR2x2_ASAP7_75t_L g348 ( .A(n_286), .B(n_321), .Y(n_348) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2x1p5_ASAP7_75t_L g359 ( .A(n_289), .B(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_289), .B(n_293), .Y(n_446) );
INVx1_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
NOR2x1_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp67_ASAP7_75t_SL g376 ( .A(n_293), .B(n_377), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_302), .B1(n_303), .B2(n_307), .C1(n_309), .C2(n_310), .Y(n_294) );
AOI21xp33_ASAP7_75t_L g339 ( .A1(n_296), .A2(n_340), .B(n_345), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_297), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g464 ( .A(n_297), .Y(n_464) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_298), .Y(n_470) );
AND2x4_ASAP7_75t_L g310 ( .A(n_299), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_299), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g454 ( .A(n_299), .Y(n_454) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
AND2x2_ASAP7_75t_L g395 ( .A(n_304), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g388 ( .A(n_305), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g327 ( .A(n_306), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_329), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_323), .B2(n_327), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_322), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx2_ASAP7_75t_L g377 ( .A(n_328), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_328), .B(n_333), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_328), .B(n_431), .Y(n_430) );
AOI211x1_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_335), .B(n_339), .C(n_346), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_330), .A2(n_444), .B(n_445), .Y(n_443) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g396 ( .A(n_332), .B(n_333), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_333), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g389 ( .A(n_333), .Y(n_389) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g453 ( .A(n_336), .B(n_434), .Y(n_453) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g351 ( .A(n_338), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_338), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g371 ( .A(n_344), .B(n_363), .Y(n_371) );
OR2x2_ASAP7_75t_L g472 ( .A(n_344), .B(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_348), .Y(n_405) );
INVx2_ASAP7_75t_L g442 ( .A(n_348), .Y(n_442) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND5xp2_ASAP7_75t_L g448 ( .A(n_351), .B(n_401), .C(n_449), .D(n_452), .E(n_454), .Y(n_448) );
AND2x2_ASAP7_75t_L g419 ( .A(n_353), .B(n_420), .Y(n_419) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_392), .Y(n_354) );
NAND2xp67_ASAP7_75t_SL g355 ( .A(n_356), .B(n_373), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_361), .B1(n_366), .B2(n_367), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g361 ( .A(n_362), .B(n_364), .C(n_365), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g398 ( .A(n_365), .Y(n_398) );
NAND3xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_371), .C(n_372), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g391 ( .A(n_370), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_SL g403 ( .A1(n_371), .A2(n_404), .B(n_405), .C(n_406), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B1(n_378), .B2(n_379), .C(n_383), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_380), .B(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_388), .B2(n_390), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_384), .A2(n_410), .B(n_436), .C(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g399 ( .A(n_385), .Y(n_399) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g424 ( .A(n_387), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_397), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g402 ( .A(n_396), .Y(n_402) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_400), .C(n_403), .Y(n_397) );
AND3x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_435), .C(n_443), .Y(n_408) );
AOI221x1_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_417), .B1(n_419), .B2(n_421), .C(n_423), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_430), .B2(n_433), .Y(n_423) );
INVx1_ASAP7_75t_L g437 ( .A(n_428), .Y(n_437) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AOI211x1_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_455), .B(n_461), .C(n_476), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_468), .B1(n_471), .B2(n_475), .Y(n_465) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_482), .B(n_841), .Y(n_840) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g821 ( .A(n_483), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_483), .B(n_830), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_483), .B(n_843), .Y(n_847) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_819), .B(n_825), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_814), .B1(n_817), .B2(n_818), .Y(n_485) );
INVx2_ASAP7_75t_L g817 ( .A(n_486), .Y(n_817) );
AO22x2_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_809), .B1(n_810), .B2(n_813), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
NOR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_723), .Y(n_488) );
NAND4xp75_ASAP7_75t_L g489 ( .A(n_490), .B(n_628), .C(n_670), .D(n_694), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI211xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_528), .B(n_569), .C(n_607), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g714 ( .A(n_494), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g808 ( .A(n_494), .B(n_745), .Y(n_808) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g623 ( .A(n_496), .B(n_579), .Y(n_623) );
AND2x2_ASAP7_75t_L g664 ( .A(n_496), .B(n_625), .Y(n_664) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g575 ( .A(n_497), .B(n_517), .Y(n_575) );
OR2x2_ASAP7_75t_L g593 ( .A(n_497), .B(n_517), .Y(n_593) );
INVx2_ASAP7_75t_L g615 ( .A(n_497), .Y(n_615) );
AND2x2_ASAP7_75t_L g645 ( .A(n_497), .B(n_579), .Y(n_645) );
AND2x2_ASAP7_75t_L g674 ( .A(n_497), .B(n_516), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_497), .B(n_626), .Y(n_710) );
AND2x2_ASAP7_75t_L g687 ( .A(n_503), .B(n_616), .Y(n_687) );
INVx2_ASAP7_75t_L g782 ( .A(n_503), .Y(n_782) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_516), .Y(n_503) );
INVx2_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
AND2x4_ASAP7_75t_L g613 ( .A(n_504), .B(n_517), .Y(n_613) );
AOI21x1_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_510), .B(n_513), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI21x1_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_507), .A2(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_515), .A2(n_535), .B(n_542), .Y(n_534) );
AND2x2_ASAP7_75t_L g772 ( .A(n_516), .B(n_574), .Y(n_772) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g636 ( .A(n_517), .Y(n_636) );
AND2x2_ASAP7_75t_L g693 ( .A(n_517), .B(n_579), .Y(n_693) );
AND2x2_ASAP7_75t_L g708 ( .A(n_517), .B(n_616), .Y(n_708) );
AND2x2_ASAP7_75t_L g730 ( .A(n_517), .B(n_574), .Y(n_730) );
OAI211xp5_ASAP7_75t_SL g777 ( .A1(n_528), .A2(n_778), .B(n_780), .C(n_787), .Y(n_777) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_555), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g764 ( .A(n_531), .B(n_700), .Y(n_764) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_546), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_532), .B(n_557), .Y(n_663) );
INVxp67_ASAP7_75t_L g677 ( .A(n_532), .Y(n_677) );
AND2x2_ASAP7_75t_L g697 ( .A(n_532), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_532), .B(n_610), .Y(n_704) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g597 ( .A(n_533), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_538), .B(n_540), .Y(n_535) );
BUFx4f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_541), .B(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g638 ( .A(n_546), .B(n_620), .Y(n_638) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g686 ( .A(n_547), .B(n_597), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_547), .B(n_600), .Y(n_692) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g596 ( .A(n_548), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g661 ( .A(n_548), .B(n_600), .Y(n_661) );
BUFx2_ASAP7_75t_L g668 ( .A(n_548), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_548), .B(n_600), .Y(n_748) );
INVx1_ASAP7_75t_L g591 ( .A(n_552), .Y(n_591) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g678 ( .A(n_556), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g807 ( .A(n_556), .B(n_596), .Y(n_807) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g610 ( .A(n_557), .Y(n_610) );
AND2x2_ASAP7_75t_L g621 ( .A(n_557), .B(n_600), .Y(n_621) );
AND2x2_ASAP7_75t_L g667 ( .A(n_557), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g700 ( .A(n_557), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_557), .B(n_611), .Y(n_717) );
AND2x2_ASAP7_75t_L g756 ( .A(n_557), .B(n_757), .Y(n_756) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_565), .B(n_568), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_576), .B(n_594), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_571), .A2(n_735), .B1(n_736), .B2(n_738), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
AND2x2_ASAP7_75t_L g732 ( .A(n_572), .B(n_623), .Y(n_732) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g647 ( .A(n_573), .Y(n_647) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g796 ( .A(n_574), .B(n_616), .Y(n_796) );
AND2x2_ASAP7_75t_L g760 ( .A(n_575), .B(n_655), .Y(n_760) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_592), .Y(n_576) );
OR2x2_ASAP7_75t_L g657 ( .A(n_577), .B(n_634), .Y(n_657) );
OR2x2_ASAP7_75t_L g769 ( .A(n_577), .B(n_593), .Y(n_769) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g632 ( .A(n_578), .Y(n_632) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
BUFx3_ASAP7_75t_L g698 ( .A(n_579), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_587), .B(n_590), .Y(n_581) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g766 ( .A(n_593), .B(n_625), .Y(n_766) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
AND2x2_ASAP7_75t_L g608 ( .A(n_596), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g649 ( .A(n_596), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g786 ( .A(n_596), .Y(n_786) );
INVx1_ASAP7_75t_L g805 ( .A(n_596), .Y(n_805) );
INVx2_ASAP7_75t_L g620 ( .A(n_597), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_597), .B(n_600), .Y(n_669) );
INVx1_ASAP7_75t_L g733 ( .A(n_598), .Y(n_733) );
BUFx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g794 ( .A(n_599), .Y(n_794) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g611 ( .A(n_600), .Y(n_611) );
INVx1_ASAP7_75t_L g701 ( .A(n_600), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_612), .B1(n_617), .B2(n_622), .Y(n_607) );
AND2x4_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_L g650 ( .A(n_610), .Y(n_650) );
AND2x2_ASAP7_75t_L g652 ( .A(n_610), .B(n_637), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_610), .B(n_620), .Y(n_712) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx3_ASAP7_75t_L g643 ( .A(n_613), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_613), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g737 ( .A(n_613), .B(n_721), .Y(n_737) );
INVx1_ASAP7_75t_L g641 ( .A(n_614), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_614), .A2(n_652), .B1(n_653), .B2(n_658), .C1(n_664), .C2(n_665), .Y(n_651) );
OAI21xp33_ASAP7_75t_SL g681 ( .A1(n_614), .A2(n_682), .B(n_683), .Y(n_681) );
AND2x2_ASAP7_75t_L g705 ( .A(n_614), .B(n_624), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_614), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OR2x2_ASAP7_75t_L g634 ( .A(n_615), .B(n_626), .Y(n_634) );
INVx1_ASAP7_75t_L g722 ( .A(n_615), .Y(n_722) );
BUFx2_ASAP7_75t_L g656 ( .A(n_616), .Y(n_656) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_619), .B(n_660), .Y(n_689) );
OR2x2_ASAP7_75t_L g801 ( .A(n_619), .B(n_661), .Y(n_801) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g684 ( .A(n_621), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g799 ( .A(n_621), .Y(n_799) );
OAI31xp33_ASAP7_75t_L g780 ( .A1(n_622), .A2(n_781), .A3(n_783), .B(n_784), .Y(n_780) );
AND2x4_ASAP7_75t_SL g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_623), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_651), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_637), .B(n_639), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x6_ASAP7_75t_L g750 ( .A(n_632), .B(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g682 ( .A(n_635), .Y(n_682) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g773 ( .A(n_636), .B(n_710), .Y(n_773) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_638), .A2(n_727), .B1(n_729), .B2(n_731), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g787 ( .A1(n_638), .A2(n_699), .B(n_761), .C(n_788), .Y(n_787) );
AOI21xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_644), .B(n_648), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND4xp25_ASAP7_75t_L g740 ( .A(n_643), .B(n_741), .C(n_742), .D(n_744), .Y(n_740) );
NAND2x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_645), .B(n_647), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_645), .B(n_730), .Y(n_753) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g719 ( .A(n_650), .B(n_679), .Y(n_719) );
NAND2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_657), .A2(n_801), .B1(n_802), .B2(n_804), .Y(n_800) );
AOI221x1_ASAP7_75t_L g739 ( .A1(n_658), .A2(n_740), .B1(n_746), .B2(n_749), .C(n_752), .Y(n_739) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g679 ( .A(n_661), .Y(n_679) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g691 ( .A(n_663), .B(n_692), .Y(n_691) );
NAND2x1p5_ASAP7_75t_L g754 ( .A(n_664), .B(n_745), .Y(n_754) );
O2A1O1Ixp5_ASAP7_75t_L g767 ( .A1(n_665), .A2(n_749), .B(n_768), .C(n_770), .Y(n_767) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx2_ASAP7_75t_L g716 ( .A(n_668), .Y(n_716) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_680), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_672), .A2(n_690), .B1(n_760), .B2(n_761), .C(n_763), .Y(n_759) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g696 ( .A(n_674), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_674), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g795 ( .A(n_674), .B(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
NAND2x1_ASAP7_75t_L g774 ( .A(n_677), .B(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g798 ( .A(n_677), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g738 ( .A(n_678), .Y(n_738) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B1(n_687), .B2(n_688), .C1(n_690), .C2(n_693), .Y(n_680) );
INVx1_ASAP7_75t_L g765 ( .A(n_684), .Y(n_765) );
INVx1_ASAP7_75t_L g728 ( .A(n_685), .Y(n_728) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g762 ( .A(n_686), .Y(n_762) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g703 ( .A(n_692), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g757 ( .A(n_692), .Y(n_757) );
AND2x2_ASAP7_75t_L g720 ( .A(n_693), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_713), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_699), .B1(n_702), .B2(n_705), .C1(n_706), .C2(n_711), .Y(n_695) );
INVx3_ASAP7_75t_L g745 ( .A(n_698), .Y(n_745) );
BUFx2_ASAP7_75t_L g803 ( .A(n_698), .Y(n_803) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g775 ( .A(n_700), .Y(n_775) );
OR2x2_ASAP7_75t_L g785 ( .A(n_700), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx2_ASAP7_75t_SL g743 ( .A(n_708), .Y(n_743) );
AND2x2_ASAP7_75t_L g788 ( .A(n_709), .B(n_745), .Y(n_788) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_710), .Y(n_741) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g747 ( .A(n_712), .B(n_748), .Y(n_747) );
NOR2x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
OR2x2_ASAP7_75t_L g804 ( .A(n_717), .B(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx1_ASAP7_75t_L g735 ( .A(n_719), .Y(n_735) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g742 ( .A(n_722), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g792 ( .A(n_722), .Y(n_792) );
NAND4xp75_ASAP7_75t_L g723 ( .A(n_724), .B(n_758), .C(n_776), .D(n_789), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_739), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_733), .B(n_734), .Y(n_725) );
INVxp33_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_728), .B(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g751 ( .A(n_730), .Y(n_751) );
AND2x2_ASAP7_75t_L g791 ( .A(n_730), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g761 ( .A(n_733), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g779 ( .A(n_744), .Y(n_779) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp33_ASAP7_75t_SL g770 ( .A1(n_747), .A2(n_771), .B1(n_773), .B2(n_774), .Y(n_770) );
INVx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI21xp33_ASAP7_75t_SL g752 ( .A1(n_753), .A2(n_754), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g783 ( .A(n_754), .Y(n_783) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_767), .Y(n_758) );
AOI21xp5_ASAP7_75t_SL g763 ( .A1(n_764), .A2(n_765), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx3_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_806), .Y(n_789) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_793), .B1(n_795), .B2(n_797), .C(n_800), .Y(n_790) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx12f_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g831 ( .A(n_812), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g818 ( .A(n_814), .Y(n_818) );
BUFx12f_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
AND2x6_ASAP7_75t_SL g820 ( .A(n_821), .B(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
INVx5_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
BUFx10_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
INVx8_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
OR2x6_ASAP7_75t_L g838 ( .A(n_839), .B(n_843), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OR2x4_ASAP7_75t_L g846 ( .A(n_841), .B(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
CKINVDCx16_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
BUFx10_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
endmodule