module real_jpeg_27033_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_300;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_299;
wire n_173;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_244;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx5_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_1),
.A2(n_40),
.B1(n_47),
.B2(n_50),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_3),
.A2(n_76),
.B1(n_77),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_3),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_128),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_128),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_3),
.A2(n_47),
.B1(n_50),
.B2(n_128),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_4),
.A2(n_76),
.B1(n_77),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_4),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_156),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_156),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_4),
.A2(n_47),
.B1(n_50),
.B2(n_156),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_57),
.B1(n_76),
.B2(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_7),
.A2(n_47),
.B1(n_50),
.B2(n_57),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_8),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_8),
.A2(n_76),
.B1(n_77),
.B2(n_150),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_150),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_8),
.A2(n_47),
.B1(n_50),
.B2(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_9),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_9),
.B(n_72),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_29),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_29),
.B(n_195),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_154),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_9),
.A2(n_47),
.B(n_51),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_9),
.B(n_122),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_9),
.A2(n_89),
.B1(n_95),
.B2(n_243),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_38),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_172)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_49),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_44),
.B1(n_47),
.B2(n_50),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_12),
.A2(n_44),
.B1(n_76),
.B2(n_77),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_19),
.B(n_105),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_86),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_58),
.B2(n_59),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_69),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_25),
.A2(n_33),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_25),
.A2(n_33),
.B1(n_149),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_25),
.A2(n_33),
.B1(n_181),
.B2(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_27),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g196 ( 
.A(n_27),
.B(n_35),
.Y(n_196)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_29),
.A2(n_30),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_29),
.B(n_73),
.Y(n_170)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_30),
.A2(n_81),
.B1(n_153),
.B2(n_170),
.Y(n_169)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_30),
.A2(n_34),
.A3(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_33),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_35),
.A2(n_49),
.B(n_154),
.C(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_37),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_42),
.A2(n_54),
.B(n_203),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_45),
.B(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_54),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_46),
.A2(n_54),
.B1(n_100),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_46),
.A2(n_52),
.B(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_46),
.A2(n_54),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_46),
.A2(n_54),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_46),
.A2(n_54),
.B1(n_202),
.B2(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_46),
.B(n_154),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_50),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_54),
.A2(n_63),
.B(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_70),
.B1(n_84),
.B2(n_85),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_66),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_66),
.A2(n_68),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B(n_79),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_71),
.A2(n_126),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_71),
.A2(n_126),
.B1(n_127),
.B2(n_162),
.Y(n_279)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_73),
.B(n_77),
.C(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_72),
.B(n_103),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_72),
.A2(n_80),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_77),
.Y(n_81)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g153 ( 
.A(n_77),
.B(n_154),
.CON(n_153),
.SN(n_153)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_98),
.B(n_102),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_102),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_88),
.A2(n_99),
.B1(n_109),
.B2(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B(n_96),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_89),
.A2(n_93),
.B1(n_141),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_89),
.A2(n_118),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_89),
.A2(n_235),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_90),
.A2(n_97),
.B(n_143),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_90),
.A2(n_94),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_97),
.Y(n_118)
);

INVx11_ASAP7_75t_L g244 ( 
.A(n_94),
.Y(n_244)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_117),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_95),
.A2(n_115),
.B(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_95),
.B(n_154),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_99),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_111),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_106),
.B(n_110),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_111),
.A2(n_112),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_121),
.C(n_124),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_114),
.B(n_119),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_121),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_299),
.B(n_304),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_286),
.B(n_298),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_185),
.B(n_267),
.C(n_285),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_173),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_136),
.B(n_173),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_157),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_138),
.B(n_144),
.C(n_157),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_139),
.B(n_140),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_152),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_168),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_159),
.B(n_164),
.C(n_168),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_167),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_171),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_179),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_174),
.A2(n_175),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_184),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_266),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_259),
.B(n_265),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_213),
.B(n_258),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_204),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_189),
.B(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_197),
.C(n_200),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_190),
.A2(n_191),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_193),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_205),
.B(n_211),
.C(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_252),
.B(n_257),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_231),
.B(n_251),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_223),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_216),
.B(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_221),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_239),
.B(n_250),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_237),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_245),
.B(n_249),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_283),
.B2(n_284),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.C(n_284),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_278),
.C(n_281),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_295),
.C(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);


endmodule