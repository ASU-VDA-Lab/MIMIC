module real_aes_7776_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g244 ( .A1(n_0), .A2(n_245), .B(n_246), .C(n_250), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_1), .B(n_186), .Y(n_251) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_2), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g468 ( .A(n_2), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_3), .B(n_158), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_4), .A2(n_144), .B(n_149), .C(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_5), .A2(n_139), .B(n_554), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_6), .A2(n_139), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_7), .B(n_186), .Y(n_560) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_8), .A2(n_174), .B(n_190), .Y(n_189) );
AND2x6_ASAP7_75t_L g144 ( .A(n_9), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_10), .A2(n_144), .B(n_149), .C(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g498 ( .A(n_11), .Y(n_498) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_12), .B(n_41), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_13), .B(n_249), .Y(n_518) );
INVx1_ASAP7_75t_L g168 ( .A(n_14), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_15), .B(n_158), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_16), .A2(n_159), .B(n_506), .C(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_17), .B(n_186), .Y(n_509) );
AOI22xp5_ASAP7_75t_SL g473 ( .A1(n_18), .A2(n_466), .B1(n_474), .B2(n_755), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_19), .A2(n_47), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_19), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_19), .B(n_223), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_20), .A2(n_149), .B(n_200), .C(n_219), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_21), .A2(n_198), .B(n_248), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_22), .B(n_249), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_23), .B(n_249), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_24), .Y(n_545) );
INVx1_ASAP7_75t_L g537 ( .A(n_25), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_26), .A2(n_149), .B(n_193), .C(n_200), .Y(n_192) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_27), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_28), .Y(n_514) );
INVx1_ASAP7_75t_L g594 ( .A(n_29), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_30), .A2(n_139), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g142 ( .A(n_31), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_32), .A2(n_147), .B(n_162), .C(n_208), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_33), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_34), .A2(n_248), .B(n_557), .C(n_559), .Y(n_556) );
INVxp67_ASAP7_75t_L g595 ( .A(n_35), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_36), .A2(n_46), .B1(n_130), .B2(n_131), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_36), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_37), .B(n_195), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_38), .A2(n_149), .B(n_200), .C(n_536), .Y(n_535) );
CKINVDCx14_ASAP7_75t_R g555 ( .A(n_39), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_40), .A2(n_45), .B1(n_481), .B2(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_40), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_41), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_42), .A2(n_250), .B(n_496), .C(n_497), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_43), .B(n_217), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_44), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_45), .Y(n_481) );
INVx1_ASAP7_75t_L g131 ( .A(n_46), .Y(n_131) );
INVx1_ASAP7_75t_L g127 ( .A(n_47), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_48), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_49), .B(n_139), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_50), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_51), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_52), .A2(n_147), .B(n_152), .C(n_162), .Y(n_146) );
INVx1_ASAP7_75t_L g247 ( .A(n_53), .Y(n_247) );
INVx1_ASAP7_75t_L g153 ( .A(n_54), .Y(n_153) );
INVx1_ASAP7_75t_L g526 ( .A(n_55), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_56), .B(n_139), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_57), .Y(n_226) );
CKINVDCx14_ASAP7_75t_R g494 ( .A(n_58), .Y(n_494) );
INVx1_ASAP7_75t_L g145 ( .A(n_59), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_60), .B(n_139), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_61), .B(n_186), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_62), .A2(n_180), .B(n_182), .C(n_184), .Y(n_179) );
INVx1_ASAP7_75t_L g167 ( .A(n_63), .Y(n_167) );
INVx1_ASAP7_75t_SL g558 ( .A(n_64), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_65), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_66), .B(n_158), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_67), .B(n_186), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_68), .B(n_159), .Y(n_261) );
INVx1_ASAP7_75t_L g548 ( .A(n_69), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_70), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_71), .B(n_155), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_72), .A2(n_149), .B(n_162), .C(n_232), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_73), .Y(n_178) );
INVx1_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_75), .A2(n_139), .B(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_76), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_77), .A2(n_139), .B(n_503), .Y(n_502) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_78), .A2(n_476), .B1(n_477), .B2(n_483), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_78), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_79), .A2(n_217), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g504 ( .A(n_80), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_81), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_82), .B(n_154), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_83), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_83), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_84), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_85), .A2(n_139), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g507 ( .A(n_86), .Y(n_507) );
INVx2_ASAP7_75t_L g165 ( .A(n_87), .Y(n_165) );
INVx1_ASAP7_75t_L g517 ( .A(n_88), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_89), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_90), .A2(n_105), .B1(n_117), .B2(n_760), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_91), .B(n_249), .Y(n_262) );
INVx2_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
OR2x2_ASAP7_75t_L g465 ( .A(n_92), .B(n_466), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_93), .A2(n_149), .B(n_162), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_94), .B(n_139), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_95), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g209 ( .A(n_96), .Y(n_209) );
INVxp67_ASAP7_75t_L g183 ( .A(n_97), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_98), .B(n_174), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_99), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g233 ( .A(n_100), .Y(n_233) );
INVx1_ASAP7_75t_L g257 ( .A(n_101), .Y(n_257) );
INVx2_ASAP7_75t_L g529 ( .A(n_102), .Y(n_529) );
AND2x2_ASAP7_75t_L g169 ( .A(n_103), .B(n_164), .Y(n_169) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g760 ( .A(n_107), .Y(n_760) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g485 ( .A(n_113), .Y(n_485) );
INVx1_ASAP7_75t_L g754 ( .A(n_113), .Y(n_754) );
NOR2x2_ASAP7_75t_L g757 ( .A(n_113), .B(n_466), .Y(n_757) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_472), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g759 ( .A(n_121), .Y(n_759) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_462), .B(n_470), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_128), .Y(n_124) );
XOR2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_132), .A2(n_485), .B1(n_486), .B2(n_753), .Y(n_484) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR5x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_335), .C(n_413), .D(n_437), .E(n_454), .Y(n_133) );
OAI211xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_201), .B(n_252), .C(n_312), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_170), .Y(n_135) );
AND2x2_ASAP7_75t_L g266 ( .A(n_136), .B(n_172), .Y(n_266) );
INVx5_ASAP7_75t_SL g294 ( .A(n_136), .Y(n_294) );
AND2x2_ASAP7_75t_L g330 ( .A(n_136), .B(n_315), .Y(n_330) );
OR2x2_ASAP7_75t_L g369 ( .A(n_136), .B(n_171), .Y(n_369) );
OR2x2_ASAP7_75t_L g400 ( .A(n_136), .B(n_291), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_136), .B(n_304), .Y(n_436) );
AND2x2_ASAP7_75t_L g448 ( .A(n_136), .B(n_291), .Y(n_448) );
OR2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_169), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_146), .B(n_164), .Y(n_137) );
BUFx2_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_140), .B(n_144), .Y(n_258) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
INVx1_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
INVx1_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_143), .Y(n_159) );
INVx1_ASAP7_75t_L g195 ( .A(n_143), .Y(n_195) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_143), .Y(n_249) );
INVx4_ASAP7_75t_SL g163 ( .A(n_144), .Y(n_163) );
BUFx3_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_148), .A2(n_163), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_148), .A2(n_163), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_148), .A2(n_163), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_148), .A2(n_163), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_148), .A2(n_163), .B(n_526), .C(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_148), .A2(n_163), .B(n_555), .C(n_556), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_SL g590 ( .A1(n_148), .A2(n_163), .B(n_591), .C(n_592), .Y(n_590) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx3_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_150), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .C(n_160), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_154), .A2(n_160), .B(n_209), .C(n_210), .Y(n_208) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_154), .A2(n_517), .B(n_518), .C(n_519), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_154), .A2(n_519), .B(n_548), .C(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_158), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g245 ( .A(n_158), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_158), .A2(n_222), .B(n_537), .C(n_538), .Y(n_536) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_158), .A2(n_181), .B1(n_594), .B2(n_595), .Y(n_593) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_159), .B(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g250 ( .A(n_161), .Y(n_250) );
INVx1_ASAP7_75t_L g508 ( .A(n_161), .Y(n_508) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_164), .A2(n_206), .B(n_207), .Y(n_205) );
INVx2_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_164), .Y(n_227) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_164), .A2(n_492), .B(n_499), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_164), .A2(n_258), .B(n_534), .C(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_165), .B(n_166), .Y(n_164) );
AND2x2_ASAP7_75t_L g175 ( .A(n_165), .B(n_166), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AND2x2_ASAP7_75t_L g447 ( .A(n_170), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
OR2x2_ASAP7_75t_L g310 ( .A(n_171), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_188), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_172), .B(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_172), .Y(n_303) );
INVx3_ASAP7_75t_L g318 ( .A(n_172), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_172), .B(n_188), .Y(n_342) );
OR2x2_ASAP7_75t_L g351 ( .A(n_172), .B(n_294), .Y(n_351) );
AND2x2_ASAP7_75t_L g355 ( .A(n_172), .B(n_315), .Y(n_355) );
AND2x2_ASAP7_75t_L g361 ( .A(n_172), .B(n_362), .Y(n_361) );
INVxp67_ASAP7_75t_L g398 ( .A(n_172), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_172), .B(n_255), .Y(n_412) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_185), .Y(n_172) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_173), .A2(n_502), .B(n_509), .Y(n_501) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_173), .A2(n_524), .B(n_530), .Y(n_523) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_173), .A2(n_553), .B(n_560), .Y(n_552) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g187 ( .A(n_174), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_174), .A2(n_191), .B(n_192), .Y(n_190) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g265 ( .A(n_175), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_180), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_181), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_181), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g222 ( .A(n_184), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_184), .B(n_593), .Y(n_592) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_186), .A2(n_241), .B(n_251), .Y(n_240) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_187), .B(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_187), .A2(n_230), .B(n_238), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_187), .B(n_239), .Y(n_238) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_187), .A2(n_256), .B(n_263), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_187), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_187), .B(n_540), .Y(n_539) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_187), .A2(n_544), .B(n_550), .Y(n_543) );
OR2x2_ASAP7_75t_L g304 ( .A(n_188), .B(n_255), .Y(n_304) );
AND2x2_ASAP7_75t_L g315 ( .A(n_188), .B(n_291), .Y(n_315) );
AND2x2_ASAP7_75t_L g327 ( .A(n_188), .B(n_318), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_188), .B(n_255), .Y(n_350) );
INVx1_ASAP7_75t_SL g362 ( .A(n_188), .Y(n_362) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g254 ( .A(n_189), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_189), .B(n_294), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B(n_197), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_197), .A2(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
AND2x2_ASAP7_75t_L g275 ( .A(n_203), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_203), .B(n_228), .Y(n_279) );
AND2x2_ASAP7_75t_L g282 ( .A(n_203), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_203), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g307 ( .A(n_203), .B(n_298), .Y(n_307) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_203), .Y(n_326) );
AND2x2_ASAP7_75t_L g347 ( .A(n_203), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g357 ( .A(n_203), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g403 ( .A(n_203), .B(n_286), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_203), .B(n_309), .Y(n_430) );
INVx5_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g300 ( .A(n_204), .Y(n_300) );
AND2x2_ASAP7_75t_L g366 ( .A(n_204), .B(n_298), .Y(n_366) );
AND2x2_ASAP7_75t_L g450 ( .A(n_204), .B(n_318), .Y(n_450) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_211), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_213), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_213), .Y(n_439) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_228), .Y(n_213) );
AND2x2_ASAP7_75t_L g269 ( .A(n_214), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g278 ( .A(n_214), .B(n_276), .Y(n_278) );
INVx5_ASAP7_75t_L g286 ( .A(n_214), .Y(n_286) );
AND2x2_ASAP7_75t_L g309 ( .A(n_214), .B(n_240), .Y(n_309) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_214), .Y(n_346) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
AOI21xp5_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_218), .B(n_223), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_224), .B(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_227), .A2(n_513), .B(n_520), .Y(n_512) );
INVx1_ASAP7_75t_L g387 ( .A(n_228), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_228), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g420 ( .A(n_228), .B(n_286), .Y(n_420) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_228), .A2(n_343), .B(n_450), .C(n_451), .Y(n_449) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_240), .Y(n_228) );
BUFx2_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
INVx2_ASAP7_75t_L g274 ( .A(n_229), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g559 ( .A(n_236), .Y(n_559) );
INVx2_ASAP7_75t_L g276 ( .A(n_240), .Y(n_276) );
AND2x2_ASAP7_75t_L g283 ( .A(n_240), .B(n_274), .Y(n_283) );
AND2x2_ASAP7_75t_L g374 ( .A(n_240), .B(n_286), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_248), .B(n_558), .Y(n_557) );
INVx4_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g496 ( .A(n_249), .Y(n_496) );
INVx2_ASAP7_75t_L g519 ( .A(n_250), .Y(n_519) );
AOI211x1_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_267), .B(n_280), .C(n_305), .Y(n_252) );
INVx1_ASAP7_75t_L g371 ( .A(n_253), .Y(n_371) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_266), .Y(n_253) );
INVx5_ASAP7_75t_SL g291 ( .A(n_255), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_255), .B(n_361), .Y(n_360) );
AOI311xp33_ASAP7_75t_L g379 ( .A1(n_255), .A2(n_380), .A3(n_382), .B(n_383), .C(n_389), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_255), .A2(n_327), .B(n_415), .C(n_418), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_259), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_258), .A2(n_514), .B(n_515), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_258), .A2(n_545), .B(n_546), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g587 ( .A(n_265), .Y(n_587) );
INVxp67_ASAP7_75t_L g334 ( .A(n_266), .Y(n_334) );
NAND4xp25_ASAP7_75t_SL g267 ( .A(n_268), .B(n_271), .C(n_277), .D(n_279), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_268), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g325 ( .A(n_269), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_272), .B(n_278), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_272), .B(n_285), .Y(n_405) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_273), .B(n_286), .Y(n_423) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g298 ( .A(n_274), .Y(n_298) );
INVxp67_ASAP7_75t_L g333 ( .A(n_275), .Y(n_333) );
AND2x4_ASAP7_75t_L g285 ( .A(n_276), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g359 ( .A(n_276), .B(n_298), .Y(n_359) );
INVx1_ASAP7_75t_L g386 ( .A(n_276), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_276), .B(n_373), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_277), .B(n_347), .Y(n_367) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_278), .B(n_300), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_278), .B(n_347), .Y(n_446) );
INVx1_ASAP7_75t_L g457 ( .A(n_279), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B(n_287), .C(n_295), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g299 ( .A(n_283), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g337 ( .A(n_283), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
AND2x2_ASAP7_75t_L g296 ( .A(n_285), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_285), .B(n_347), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_285), .B(n_366), .Y(n_390) );
OR2x2_ASAP7_75t_L g306 ( .A(n_286), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_286), .B(n_298), .Y(n_353) );
AND2x2_ASAP7_75t_L g410 ( .A(n_286), .B(n_366), .Y(n_410) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_286), .Y(n_417) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_288), .A2(n_300), .B1(n_422), .B2(n_424), .C(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g311 ( .A(n_291), .B(n_294), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_291), .B(n_361), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_291), .B(n_318), .Y(n_426) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g411 ( .A(n_293), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g425 ( .A(n_293), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_294), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_315), .Y(n_322) );
AND2x2_ASAP7_75t_L g392 ( .A(n_294), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_294), .B(n_341), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_294), .B(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_299), .B(n_301), .Y(n_295) );
INVx2_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
OR2x2_ASAP7_75t_L g352 ( .A(n_300), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g455 ( .A(n_300), .B(n_423), .Y(n_455) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AOI21xp33_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_308), .B(n_310), .Y(n_305) );
INVx1_ASAP7_75t_L g459 ( .A(n_306), .Y(n_459) );
INVx2_ASAP7_75t_SL g373 ( .A(n_307), .Y(n_373) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_310), .A2(n_391), .B(n_455), .C(n_456), .Y(n_454) );
OAI322xp33_ASAP7_75t_SL g323 ( .A1(n_311), .A2(n_324), .A3(n_327), .B1(n_328), .B2(n_329), .C1(n_331), .C2(n_334), .Y(n_323) );
INVx2_ASAP7_75t_L g343 ( .A(n_311), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .B1(n_320), .B2(n_322), .C(n_323), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp33_ASAP7_75t_SL g389 ( .A1(n_314), .A2(n_390), .B1(n_391), .B2(n_394), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_315), .B(n_318), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_315), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g388 ( .A(n_317), .B(n_350), .Y(n_388) );
INVx1_ASAP7_75t_L g378 ( .A(n_318), .Y(n_378) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_322), .A2(n_432), .B(n_434), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_324), .A2(n_357), .B(n_360), .Y(n_356) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2xp67_ASAP7_75t_SL g385 ( .A(n_326), .B(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_326), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g442 ( .A(n_327), .Y(n_442) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND4xp25_ASAP7_75t_L g335 ( .A(n_336), .B(n_363), .C(n_379), .D(n_395), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B(n_344), .C(n_356), .Y(n_336) );
INVx1_ASAP7_75t_L g428 ( .A(n_337), .Y(n_428) );
AND2x2_ASAP7_75t_L g376 ( .A(n_338), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_343), .B(n_378), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B1(n_352), .B2(n_354), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_346), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g408 ( .A1(n_347), .A2(n_386), .B(n_409), .C(n_411), .Y(n_408) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g393 ( .A(n_350), .Y(n_393) );
INVx1_ASAP7_75t_L g453 ( .A(n_351), .Y(n_453) );
NAND2xp33_ASAP7_75t_SL g443 ( .A(n_352), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B(n_368), .C(n_370), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_375), .B2(n_377), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_373), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_378), .B(n_399), .Y(n_461) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI21xp33_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_387), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_401), .B1(n_404), .B2(n_406), .C(n_408), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_411), .A2(n_428), .B1(n_429), .B2(n_430), .Y(n_427) );
NAND3xp33_ASAP7_75t_SL g413 ( .A(n_414), .B(n_421), .C(n_431), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_440), .C(n_449), .Y(n_437) );
INVx1_ASAP7_75t_L g458 ( .A(n_438), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B1(n_445), .B2(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_456) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g471 ( .A(n_465), .Y(n_471) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_470), .B(n_473), .C(n_758), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_683), .Y(n_486) );
NAND5xp2_ASAP7_75t_L g487 ( .A(n_488), .B(n_598), .C(n_630), .D(n_647), .E(n_670), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_531), .B1(n_561), .B2(n_565), .C(n_569), .Y(n_488) );
INVx1_ASAP7_75t_L g710 ( .A(n_489), .Y(n_710) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_510), .Y(n_489) );
AND3x2_ASAP7_75t_L g685 ( .A(n_490), .B(n_512), .C(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_500), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_491), .B(n_567), .Y(n_566) );
BUFx3_ASAP7_75t_L g576 ( .A(n_491), .Y(n_576) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_522), .Y(n_580) );
INVx2_ASAP7_75t_L g607 ( .A(n_491), .Y(n_607) );
OR2x2_ASAP7_75t_L g618 ( .A(n_491), .B(n_523), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_491), .B(n_511), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_491), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g697 ( .A(n_491), .B(n_523), .Y(n_697) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_500), .Y(n_579) );
AND2x2_ASAP7_75t_L g638 ( .A(n_500), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_500), .B(n_511), .Y(n_657) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_511), .Y(n_568) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_501), .Y(n_575) );
AND2x2_ASAP7_75t_L g624 ( .A(n_501), .B(n_523), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_501), .B(n_510), .C(n_607), .Y(n_649) );
AND2x2_ASAP7_75t_L g714 ( .A(n_501), .B(n_512), .Y(n_714) );
AND2x2_ASAP7_75t_L g748 ( .A(n_501), .B(n_511), .Y(n_748) );
INVxp67_ASAP7_75t_L g577 ( .A(n_510), .Y(n_577) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_511), .B(n_607), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_511), .B(n_638), .Y(n_646) );
AND2x2_ASAP7_75t_L g696 ( .A(n_511), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g724 ( .A(n_511), .Y(n_724) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g631 ( .A(n_512), .B(n_624), .Y(n_631) );
BUFx3_ASAP7_75t_L g663 ( .A(n_512), .Y(n_663) );
INVx2_ASAP7_75t_L g639 ( .A(n_522), .Y(n_639) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_523), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_531), .A2(n_699), .B1(n_701), .B2(n_702), .Y(n_698) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
AND2x2_ASAP7_75t_L g561 ( .A(n_532), .B(n_562), .Y(n_561) );
INVx3_ASAP7_75t_SL g572 ( .A(n_532), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_532), .B(n_602), .Y(n_634) );
OR2x2_ASAP7_75t_L g653 ( .A(n_532), .B(n_542), .Y(n_653) );
AND2x2_ASAP7_75t_L g658 ( .A(n_532), .B(n_610), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_532), .B(n_603), .Y(n_661) );
AND2x2_ASAP7_75t_L g673 ( .A(n_532), .B(n_552), .Y(n_673) );
AND2x2_ASAP7_75t_L g689 ( .A(n_532), .B(n_543), .Y(n_689) );
AND2x4_ASAP7_75t_L g692 ( .A(n_532), .B(n_563), .Y(n_692) );
OR2x2_ASAP7_75t_L g709 ( .A(n_532), .B(n_645), .Y(n_709) );
OR2x2_ASAP7_75t_L g740 ( .A(n_532), .B(n_585), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_532), .B(n_668), .Y(n_742) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_539), .Y(n_532) );
AND2x2_ASAP7_75t_L g616 ( .A(n_541), .B(n_583), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_541), .B(n_603), .Y(n_735) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_552), .Y(n_541) );
AND2x2_ASAP7_75t_L g571 ( .A(n_542), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g602 ( .A(n_542), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g610 ( .A(n_542), .B(n_585), .Y(n_610) );
AND2x2_ASAP7_75t_L g628 ( .A(n_542), .B(n_563), .Y(n_628) );
OR2x2_ASAP7_75t_L g645 ( .A(n_542), .B(n_603), .Y(n_645) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g564 ( .A(n_543), .Y(n_564) );
AND2x2_ASAP7_75t_L g668 ( .A(n_543), .B(n_552), .Y(n_668) );
INVx2_ASAP7_75t_L g563 ( .A(n_552), .Y(n_563) );
INVx1_ASAP7_75t_L g680 ( .A(n_552), .Y(n_680) );
AND2x2_ASAP7_75t_L g730 ( .A(n_552), .B(n_572), .Y(n_730) );
AND2x2_ASAP7_75t_L g582 ( .A(n_562), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g614 ( .A(n_562), .B(n_572), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_562), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g601 ( .A(n_563), .B(n_572), .Y(n_601) );
OR2x2_ASAP7_75t_L g717 ( .A(n_564), .B(n_691), .Y(n_717) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_567), .B(n_697), .Y(n_703) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OAI32xp33_ASAP7_75t_L g659 ( .A1(n_568), .A2(n_660), .A3(n_662), .B1(n_664), .B2(n_665), .Y(n_659) );
OR2x2_ASAP7_75t_L g676 ( .A(n_568), .B(n_618), .Y(n_676) );
OAI21xp33_ASAP7_75t_SL g701 ( .A1(n_568), .A2(n_578), .B(n_606), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B1(n_578), .B2(n_581), .Y(n_569) );
INVxp33_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_571), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_572), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g627 ( .A(n_572), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g727 ( .A(n_572), .B(n_668), .Y(n_727) );
OR2x2_ASAP7_75t_L g751 ( .A(n_572), .B(n_645), .Y(n_751) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_573), .A2(n_633), .B(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g611 ( .A(n_575), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_575), .B(n_580), .Y(n_629) );
AND2x2_ASAP7_75t_L g651 ( .A(n_576), .B(n_624), .Y(n_651) );
INVx1_ASAP7_75t_L g664 ( .A(n_576), .Y(n_664) );
OR2x2_ASAP7_75t_L g669 ( .A(n_576), .B(n_603), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_579), .B(n_618), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_580), .A2(n_600), .B1(n_605), .B2(n_609), .Y(n_599) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_583), .A2(n_642), .B1(n_649), .B2(n_650), .Y(n_648) );
AND2x2_ASAP7_75t_L g726 ( .A(n_583), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_585), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g745 ( .A(n_585), .B(n_628), .Y(n_745) );
AO21x2_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B(n_596), .Y(n_585) );
INVx1_ASAP7_75t_L g604 ( .A(n_586), .Y(n_604) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OA21x2_ASAP7_75t_L g603 ( .A1(n_589), .A2(n_597), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_611), .B1(n_612), .B2(n_617), .C(n_619), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_601), .B(n_603), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_601), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g620 ( .A(n_602), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_602), .A2(n_708), .B(n_709), .C(n_710), .Y(n_707) );
AND2x2_ASAP7_75t_L g712 ( .A(n_602), .B(n_692), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_SL g750 ( .A1(n_602), .A2(n_691), .B(n_751), .C(n_752), .Y(n_750) );
BUFx3_ASAP7_75t_L g642 ( .A(n_603), .Y(n_642) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_606), .B(n_663), .Y(n_706) );
AOI211xp5_ASAP7_75t_L g725 ( .A1(n_606), .A2(n_726), .B(n_728), .C(n_734), .Y(n_725) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVxp67_ASAP7_75t_L g686 ( .A(n_608), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_610), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_614), .A2(n_631), .B(n_632), .C(n_640), .Y(n_630) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g715 ( .A(n_618), .Y(n_715) );
OR2x2_ASAP7_75t_L g732 ( .A(n_618), .B(n_662), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_626), .B2(n_629), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_621), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
OR2x2_ASAP7_75t_L g719 ( .A(n_623), .B(n_663), .Y(n_719) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g674 ( .A(n_624), .B(n_664), .Y(n_674) );
INVx1_ASAP7_75t_L g682 ( .A(n_625), .Y(n_682) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_628), .B(n_642), .Y(n_690) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_638), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g747 ( .A(n_639), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_646), .Y(n_640) );
INVx1_ASAP7_75t_L g677 ( .A(n_641), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_642), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_642), .B(n_673), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_642), .B(n_668), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_642), .B(n_689), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_642), .A2(n_652), .B(n_692), .C(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AOI221xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_652), .B1(n_654), .B2(n_658), .C(n_659), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_656), .B(n_664), .Y(n_738) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g749 ( .A1(n_658), .A2(n_673), .B(n_675), .C(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_661), .B(n_668), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_662), .B(n_715), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g662 ( .A(n_663), .Y(n_662) );
INVxp33_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
AOI21xp33_ASAP7_75t_SL g678 ( .A1(n_667), .A2(n_679), .B(n_681), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_667), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_668), .B(n_722), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B1(n_675), .B2(n_677), .C(n_678), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_674), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g708 ( .A(n_680), .Y(n_708) );
NAND5xp2_ASAP7_75t_L g683 ( .A(n_684), .B(n_711), .C(n_725), .D(n_736), .E(n_749), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_694), .C(n_707), .Y(n_684) );
INVx2_ASAP7_75t_SL g731 ( .A(n_685), .Y(n_731) );
NAND4xp25_ASAP7_75t_SL g687 ( .A(n_688), .B(n_690), .C(n_691), .D(n_693), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_693), .A2(n_695), .B(n_698), .C(n_704), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_696), .A2(n_737), .B1(n_739), .B2(n_741), .C(n_743), .Y(n_736) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_713), .B1(n_716), .B2(n_718), .C(n_720), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_719), .A2(n_742), .B1(n_744), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule