module fake_jpeg_566_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_55;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx4f_ASAP7_75t_SL g8 ( 
.A(n_6),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_7),
.B(n_5),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_17),
.C(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_16),
.B1(n_15),
.B2(n_12),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_4),
.Y(n_24)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_11),
.B(n_10),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_17),
.B1(n_13),
.B2(n_14),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.C(n_25),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_11),
.B(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

AO32x1_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_20),
.A3(n_18),
.B1(n_23),
.B2(n_19),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_48),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_42),
.B(n_33),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.C(n_45),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_32),
.B(n_29),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.A3(n_47),
.B1(n_43),
.B2(n_20),
.C1(n_11),
.C2(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_47),
.Y(n_54)
);

OAI221xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_11),
.B1(n_21),
.B2(n_27),
.C(n_41),
.Y(n_56)
);


endmodule