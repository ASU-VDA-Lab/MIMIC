module real_jpeg_16977_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_366;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_0),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_1),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_1),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_2),
.Y(n_156)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_3),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_3),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_3),
.B(n_136),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_41),
.Y(n_240)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_5),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_5),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_5),
.B(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_5),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_5),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_5),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_5),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_6),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_6),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_6),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_7),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_7),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_11),
.B1(n_39),
.B2(n_44),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_8),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_8),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_8),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_8),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_8),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_8),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_8),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_9),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_9),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_9),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_9),
.B(n_115),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_9),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_9),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_9),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_62),
.Y(n_61)
);

AND2x4_ASAP7_75t_SL g92 ( 
.A(n_10),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_10),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_10),
.B(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_10),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_11),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_11),
.B(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_11),
.Y(n_231)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_12),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_14),
.Y(n_149)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_14),
.Y(n_290)
);

NAND2x1_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_15),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_15),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_15),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_15),
.B(n_298),
.Y(n_297)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_16),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_210),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_208),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_166),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_20),
.B(n_166),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.C(n_138),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_21),
.A2(n_22),
.B1(n_101),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_66),
.Y(n_22)
);

INVxp33_ASAP7_75t_SL g168 ( 
.A(n_23),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.C(n_50),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_24),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_28),
.C(n_32),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_37),
.A2(n_38),
.B1(n_50),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_38),
.A2(n_227),
.B(n_230),
.Y(n_226)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_50),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_61),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_51),
.A2(n_52),
.B1(n_61),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_51),
.A2(n_52),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_54),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_56),
.B(n_143),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_80),
.B1(n_99),
.B2(n_100),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_68),
.B(n_70),
.C(n_76),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_70),
.A2(n_71),
.B1(n_241),
.B2(n_242),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_71),
.B(n_236),
.C(n_241),
.Y(n_235)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_80),
.B(n_168),
.C(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_91),
.C(n_94),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_81),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.C(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_82),
.A2(n_89),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_82),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_82),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_85),
.B(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_90),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_97),
.Y(n_229)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_101),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_125),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_113),
.C(n_125),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.C(n_110),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_104),
.A2(n_110),
.B1(n_111),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_108),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_110),
.B(n_261),
.C(n_262),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_110),
.A2(n_111),
.B1(n_261),
.B2(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_114),
.B(n_118),
.C(n_121),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_118),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_118),
.A2(n_124),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_119),
.Y(n_292)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_119),
.Y(n_320)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_123),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_131),
.C(n_135),
.Y(n_183)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_139),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_160),
.C(n_163),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_140),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_151),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_142),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_145),
.B(n_151),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_146),
.B(n_150),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_149),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_152),
.A2(n_155),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_152),
.Y(n_257)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_155),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_155),
.A2(n_258),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_155),
.B(n_322),
.C(n_326),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_156),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_157),
.B(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_160),
.B(n_163),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_184),
.B1(n_206),
.B2(n_207),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_188),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_268),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_248),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_214),
.B(n_218),
.Y(n_367)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_244),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_235),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_226),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_224),
.B(n_277),
.C(n_280),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_236),
.B(n_354),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_SL g310 ( 
.A(n_237),
.B(n_240),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_237),
.A2(n_317),
.B1(n_318),
.B2(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_251),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.C(n_266),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_252),
.B(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_254),
.B(n_266),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_264),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_255),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_260),
.B(n_265),
.Y(n_359)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

XOR2x1_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.C(n_367),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_362),
.B(n_366),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_348),
.B(n_361),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_313),
.B(n_347),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_301),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_274),
.B(n_301),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.C(n_293),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_275),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_284),
.A2(n_285),
.B1(n_293),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_286),
.B(n_291),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

AO22x1_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.Y(n_293)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_294),
.Y(n_299)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_297),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_337),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_303),
.B(n_304),
.C(n_307),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_310),
.C(n_311),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_341),
.B(n_346),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_329),
.B(n_340),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_321),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_336),
.B(n_339),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_334),
.Y(n_339)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_345),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_360),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_SL g361 ( 
.A(n_349),
.B(n_360),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_357),
.B2(n_358),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_355),
.B2(n_356),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_356),
.C(n_357),
.Y(n_365)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_365),
.Y(n_366)
);


endmodule