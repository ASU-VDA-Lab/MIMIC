module fake_jpeg_14709_n_351 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_351);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_44),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_48),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_19),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_29),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_36),
.B1(n_31),
.B2(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_36),
.B1(n_33),
.B2(n_46),
.Y(n_99)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_47),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_31),
.B1(n_33),
.B2(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_66),
.B1(n_46),
.B2(n_43),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_41),
.B(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_32),
.C(n_35),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_44),
.C(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_31),
.B1(n_33),
.B2(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_76),
.B(n_88),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_17),
.B(n_37),
.C(n_27),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_85),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_26),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_91),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_55),
.B(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_100),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_106),
.C(n_51),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_101),
.B1(n_108),
.B2(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_32),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_35),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_25),
.B1(n_37),
.B2(n_17),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_18),
.B(n_37),
.C(n_23),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_70),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_25),
.B1(n_18),
.B2(n_38),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_17),
.B1(n_27),
.B2(n_25),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_65),
.B(n_27),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_65),
.B(n_23),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_21),
.B(n_34),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_117),
.A2(n_125),
.B(n_139),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_88),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_136),
.C(n_141),
.Y(n_163)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_142),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_89),
.B1(n_77),
.B2(n_97),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_28),
.B(n_35),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_21),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_38),
.B1(n_75),
.B2(n_54),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_140),
.B1(n_83),
.B2(n_93),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_70),
.B1(n_34),
.B2(n_30),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_35),
.B(n_1),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_96),
.B1(n_106),
.B2(n_94),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_51),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_35),
.C(n_34),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_0),
.B(n_1),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_89),
.C(n_102),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_146),
.B(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_157),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_153),
.B1(n_143),
.B2(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_102),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_165),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_97),
.B1(n_110),
.B2(n_77),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_128),
.B1(n_134),
.B2(n_129),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_160),
.B(n_171),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_92),
.B1(n_81),
.B2(n_93),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_166),
.B1(n_172),
.B2(n_128),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_83),
.B(n_105),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_103),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_107),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_105),
.B1(n_104),
.B2(n_87),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_169),
.Y(n_203)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_115),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_103),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_122),
.A2(n_34),
.B1(n_30),
.B2(n_24),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_173),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_86),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_84),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_118),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_140),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_189),
.C(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_196),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_141),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_121),
.C(n_142),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_200),
.C(n_204),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_211),
.B1(n_147),
.B2(n_167),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_201),
.B1(n_209),
.B2(n_147),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_177),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_160),
.C(n_154),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_117),
.A3(n_124),
.B1(n_30),
.B2(n_24),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_30),
.Y(n_202)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_24),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_24),
.B(n_21),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_208),
.B(n_175),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_4),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_9),
.C(n_14),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_172),
.C(n_149),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_2),
.B(n_3),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_152),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_215),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_217),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_182),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_220),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_180),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_187),
.B1(n_191),
.B2(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_184),
.B(n_158),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_232),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_235),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_233),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_159),
.B(n_173),
.Y(n_229)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_164),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_179),
.B(n_156),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_240),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_199),
.B(n_147),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_183),
.A2(n_169),
.B1(n_168),
.B2(n_161),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_195),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_178),
.C(n_189),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_247),
.C(n_254),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_233),
.A2(n_199),
.B1(n_186),
.B2(n_208),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_252),
.B1(n_255),
.B2(n_227),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_192),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_200),
.C(n_204),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_217),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_190),
.C(n_179),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_210),
.B1(n_185),
.B2(n_193),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_207),
.C(n_205),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_260),
.C(n_215),
.Y(n_274)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_203),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_198),
.C(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_236),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_268),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_242),
.C(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_222),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_282),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_255),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_250),
.B(n_240),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_231),
.B1(n_226),
.B2(n_221),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_279),
.A2(n_286),
.B1(n_206),
.B2(n_7),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_244),
.B1(n_248),
.B2(n_228),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_280),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_247),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_216),
.B1(n_237),
.B2(n_214),
.Y(n_296)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_245),
.B1(n_260),
.B2(n_231),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_274),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_299),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_277),
.B1(n_280),
.B2(n_11),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_271),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_267),
.A2(n_253),
.B(n_265),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_252),
.C(n_234),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_234),
.C(n_232),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_206),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_5),
.C(n_8),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_302),
.B(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_312),
.C(n_302),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_269),
.B(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_272),
.B1(n_283),
.B2(n_270),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_279),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_319),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_16),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_299),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_12),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_291),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_290),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_320),
.B(n_321),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_298),
.C(n_287),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_303),
.B1(n_295),
.B2(n_297),
.Y(n_322)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_328),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_307),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_329),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_13),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_310),
.C(n_315),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_322),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_305),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_335),
.Y(n_340)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_325),
.B(n_309),
.CI(n_318),
.CON(n_335),
.SN(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_324),
.A2(n_309),
.B(n_16),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_16),
.B(n_332),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_324),
.C(n_328),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_343),
.C(n_337),
.Y(n_346)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_341),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_323),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_342),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_339),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_347),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_345),
.C(n_340),
.Y(n_349)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_344),
.B(n_338),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_335),
.Y(n_351)
);


endmodule