module fake_jpeg_19268_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_43),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_17),
.B1(n_26),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_52),
.B1(n_54),
.B2(n_61),
.Y(n_71)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_17),
.B1(n_26),
.B2(n_32),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_17),
.B1(n_26),
.B2(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_19),
.B1(n_31),
.B2(n_20),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_24),
.B1(n_44),
.B2(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_34),
.B1(n_30),
.B2(n_19),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_31),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_34),
.B1(n_30),
.B2(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_77),
.B1(n_84),
.B2(n_87),
.Y(n_134)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_36),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_74),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_18),
.B1(n_23),
.B2(n_16),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_75),
.A2(n_103),
.B1(n_48),
.B2(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_44),
.B1(n_42),
.B2(n_37),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_44),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_86),
.C(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_43),
.B(n_18),
.C(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_35),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_35),
.B1(n_30),
.B2(n_34),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_97),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_43),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_28),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_105),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_46),
.A2(n_28),
.B(n_25),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_34),
.B1(n_30),
.B2(n_33),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_0),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_0),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_25),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_16),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_135),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_54),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_127),
.B(n_128),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_65),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

AO21x1_ASAP7_75t_SL g132 ( 
.A1(n_68),
.A2(n_64),
.B(n_33),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_107),
.B1(n_86),
.B2(n_78),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_69),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_104),
.B1(n_102),
.B2(n_98),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_33),
.B1(n_23),
.B2(n_16),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_124),
.B1(n_109),
.B2(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_137),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_88),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_145),
.B(n_149),
.Y(n_190)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_85),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_82),
.C(n_99),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_151),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_71),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_153),
.B1(n_167),
.B2(n_73),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_87),
.B1(n_79),
.B2(n_84),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_170),
.B1(n_115),
.B2(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_160),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_107),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_3),
.B(n_5),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_108),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_72),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_96),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_166),
.A3(n_106),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_96),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_95),
.B1(n_97),
.B2(n_86),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_95),
.C(n_105),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_1),
.C(n_2),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_127),
.B(n_122),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_140),
.B1(n_168),
.B2(n_146),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_143),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_185),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_134),
.B(n_110),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_7),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_176),
.A2(n_186),
.B(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_122),
.B1(n_114),
.B2(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_122),
.B1(n_136),
.B2(n_105),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_130),
.B1(n_103),
.B2(n_119),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_119),
.B1(n_117),
.B2(n_94),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_23),
.B(n_117),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_222)
);

FAx1_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_73),
.CI(n_94),
.CON(n_188),
.SN(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_100),
.B(n_90),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_189),
.A2(n_198),
.B(n_199),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_5),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_144),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_193),
.B1(n_147),
.B2(n_142),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_146),
.B1(n_149),
.B2(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_139),
.C(n_161),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_3),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_3),
.B(n_4),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_7),
.CI(n_9),
.CON(n_216),
.SN(n_216)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_150),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_212),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_206),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_140),
.B(n_145),
.C(n_160),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_211),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_208),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_171),
.B(n_148),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_210),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_154),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_155),
.B1(n_141),
.B2(n_6),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_141),
.B1(n_6),
.B2(n_8),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_223),
.B(n_200),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_222),
.B1(n_224),
.B2(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_12),
.C(n_14),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.C(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_15),
.C(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_183),
.B1(n_201),
.B2(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_238),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_186),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_248),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_202),
.B1(n_171),
.B2(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_206),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_173),
.C(n_189),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_207),
.C(n_209),
.Y(n_256)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_180),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_209),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_215),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_260),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_270),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_205),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_268),
.B(n_232),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_247),
.A2(n_229),
.B(n_188),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_241),
.B(n_198),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_211),
.C(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_250),
.C(n_248),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_227),
.B1(n_188),
.B2(n_222),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_213),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_278),
.B(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_231),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_247),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_240),
.B(n_242),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_283),
.C(n_273),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_233),
.B(n_251),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_261),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_238),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_253),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_243),
.C(n_225),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_262),
.C(n_264),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_289),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_279),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_255),
.B(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_257),
.C(n_261),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_179),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_259),
.B(n_249),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_297),
.B(n_249),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_179),
.C(n_184),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_281),
.C(n_282),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_299),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_271),
.B1(n_277),
.B2(n_274),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_280),
.C(n_274),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_284),
.Y(n_310)
);

OAI22x1_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_290),
.B1(n_216),
.B2(n_191),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_185),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_312),
.B(n_184),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_307),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_304),
.C(n_309),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_302),
.C(n_298),
.Y(n_319)
);

AOI321xp33_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_313),
.A3(n_310),
.B1(n_303),
.B2(n_199),
.C(n_194),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_198),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_15),
.Y(n_322)
);


endmodule