module fake_jpeg_10592_n_67 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_12),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_12),
.B(n_8),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_26),
.B1(n_11),
.B2(n_13),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_30),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_11),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_29),
.B(n_31),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_14),
.C(n_17),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_33),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_28),
.B(n_27),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_9),
.Y(n_43)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.C(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_24),
.B1(n_10),
.B2(n_22),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_19),
.B(n_2),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_14),
.C(n_9),
.Y(n_54)
);

NOR4xp25_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_38),
.C(n_5),
.D(n_24),
.Y(n_52)
);

AOI221xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_9),
.B1(n_5),
.B2(n_4),
.C(n_2),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_55),
.B(n_56),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

AOI21x1_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_51),
.B(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_54),
.B1(n_2),
.B2(n_4),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_59),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_64),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_1),
.Y(n_67)
);


endmodule