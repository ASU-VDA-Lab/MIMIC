module fake_jpeg_10863_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_44),
.B(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_9),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_9),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_51),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_15),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_67),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_37),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_108)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_37),
.B(n_19),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_104),
.B(n_1),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_40),
.B1(n_31),
.B2(n_19),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_97),
.B1(n_74),
.B2(n_82),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_37),
.B1(n_22),
.B2(n_31),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_92),
.B1(n_103),
.B2(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_91),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_40),
.B1(n_31),
.B2(n_19),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_105),
.B1(n_109),
.B2(n_15),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_39),
.B1(n_38),
.B2(n_22),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_100),
.B1(n_95),
.B2(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_25),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_43),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_30),
.C(n_32),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_6),
.C(n_10),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_35),
.B1(n_36),
.B2(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_35),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_83),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_36),
.B1(n_27),
.B2(n_39),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_63),
.A2(n_38),
.B(n_27),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_7),
.B1(n_14),
.B2(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_7),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_11),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_6),
.B1(n_13),
.B2(n_3),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_65),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_83),
.B(n_95),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_118),
.A2(n_134),
.B1(n_128),
.B2(n_120),
.Y(n_174)
);

BUFx24_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_119),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_127),
.Y(n_166)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_97),
.B1(n_80),
.B2(n_87),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_135),
.B1(n_142),
.B2(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_75),
.B(n_10),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_75),
.B(n_10),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_145),
.B(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_11),
.B1(n_15),
.B2(n_88),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_114),
.B1(n_138),
.B2(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_82),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_71),
.A2(n_81),
.B1(n_72),
.B2(n_73),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_139),
.Y(n_171)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_143),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_71),
.A2(n_81),
.B1(n_72),
.B2(n_101),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_93),
.C(n_98),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_98),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_106),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_149),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_137),
.B(n_161),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_115),
.B1(n_121),
.B2(n_147),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_173),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_113),
.B1(n_148),
.B2(n_118),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_145),
.B1(n_150),
.B2(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_125),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_165),
.B1(n_173),
.B2(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_120),
.B1(n_131),
.B2(n_117),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_146),
.B1(n_140),
.B2(n_119),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_166),
.B(n_175),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_192),
.B(n_177),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_186),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_183),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_171),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_119),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_168),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_122),
.C(n_137),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_161),
.B1(n_172),
.B2(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_153),
.B1(n_154),
.B2(n_176),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_160),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_174),
.B(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_212),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_215),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_187),
.B1(n_194),
.B2(n_190),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_214),
.B(n_218),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_177),
.B(n_169),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_184),
.B(n_190),
.Y(n_233)
);

NAND2x1p5_ASAP7_75t_R g212 ( 
.A(n_192),
.B(n_154),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_187),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_156),
.B(n_162),
.C(n_179),
.D(n_188),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_156),
.B1(n_179),
.B2(n_186),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_189),
.B1(n_181),
.B2(n_195),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_183),
.C(n_185),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_223),
.C(n_227),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_183),
.C(n_185),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_225),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_199),
.B(n_184),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_183),
.C(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_219),
.B1(n_210),
.B2(n_214),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_206),
.C(n_198),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_187),
.C(n_188),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_241),
.B1(n_226),
.B2(n_239),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_217),
.A3(n_201),
.B1(n_208),
.B2(n_213),
.C1(n_218),
.C2(n_212),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_241),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_231),
.A2(n_219),
.B1(n_191),
.B2(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_191),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_240),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_205),
.B1(n_207),
.B2(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_237),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_221),
.B(n_227),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_246),
.C(n_236),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_234),
.B(n_207),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_251),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_237),
.A2(n_193),
.B1(n_226),
.B2(n_179),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_255),
.A2(n_236),
.B1(n_245),
.B2(n_242),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_243),
.Y(n_256)
);

AOI31xp67_ASAP7_75t_SL g257 ( 
.A1(n_252),
.A2(n_248),
.A3(n_246),
.B(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_259),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_243),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_260),
.A2(n_253),
.B(n_251),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_261),
.B(n_258),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_262),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_264),
.Y(n_265)
);


endmodule