module real_aes_7886_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1106;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_994;
wire n_528;
wire n_578;
wire n_495;
wire n_892;
wire n_1072;
wire n_1078;
wire n_938;
wire n_384;
wire n_744;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_976;
wire n_872;
wire n_636;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_656;
wire n_532;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_455;
wire n_973;
wire n_725;
wire n_671;
wire n_960;
wire n_1084;
wire n_1081;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_1105;
wire n_902;
wire n_471;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_968;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_1114;
wire n_566;
wire n_719;
wire n_967;
wire n_837;
wire n_871;
wire n_1045;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_1040;
wire n_1097;
wire n_652;
wire n_500;
wire n_601;
wire n_703;
wire n_661;
wire n_463;
wire n_1102;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_1076;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_1119;
wire n_868;
wire n_877;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_0), .A2(n_163), .B1(n_567), .B2(n_709), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_1), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_2), .B(n_552), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_3), .B(n_637), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_4), .Y(n_662) );
OA22x2_ASAP7_75t_L g761 ( .A1(n_5), .A2(n_762), .B1(n_763), .B2(n_789), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_5), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g890 ( .A1(n_6), .A2(n_152), .B1(n_514), .B2(n_727), .C(n_891), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_7), .A2(n_399), .B1(n_495), .B2(n_496), .Y(n_398) );
INVx1_ASAP7_75t_L g496 ( .A(n_7), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g1023 ( .A1(n_8), .A2(n_282), .B1(n_521), .B2(n_594), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_9), .A2(n_344), .B1(n_605), .B2(n_616), .Y(n_907) );
AOI22xp5_ASAP7_75t_SL g565 ( .A1(n_10), .A2(n_379), .B1(n_566), .B2(n_567), .Y(n_565) );
AO22x2_ASAP7_75t_L g408 ( .A1(n_11), .A2(n_215), .B1(n_409), .B2(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g1071 ( .A(n_11), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_12), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_13), .A2(n_292), .B1(n_486), .B2(n_733), .Y(n_739) );
AOI22xp5_ASAP7_75t_SL g558 ( .A1(n_14), .A2(n_241), .B1(n_527), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_15), .A2(n_19), .B1(n_521), .B2(n_634), .Y(n_912) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_16), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_17), .A2(n_381), .B1(n_620), .B2(n_884), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g1031 ( .A(n_18), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_20), .A2(n_261), .B1(n_428), .B2(n_748), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g926 ( .A1(n_21), .A2(n_331), .B1(n_664), .B2(n_927), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_22), .A2(n_164), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_23), .A2(n_334), .B1(n_679), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_24), .A2(n_101), .B1(n_448), .B2(n_452), .Y(n_447) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_25), .A2(n_104), .B1(n_409), .B2(n_413), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_26), .Y(n_930) );
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_27), .A2(n_257), .B1(n_426), .B2(n_642), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_28), .A2(n_192), .B1(n_773), .B2(n_774), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_29), .A2(n_94), .B1(n_587), .B2(n_631), .Y(n_824) );
INVx1_ASAP7_75t_L g1119 ( .A(n_30), .Y(n_1119) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_31), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_32), .A2(n_316), .B1(n_448), .B2(n_610), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_33), .A2(n_220), .B1(n_503), .B2(n_504), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_34), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_35), .Y(n_1047) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_36), .A2(n_268), .B1(n_422), .B2(n_562), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_37), .B(n_593), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_38), .A2(n_266), .B1(n_535), .B2(n_593), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_39), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_40), .A2(n_326), .B1(n_525), .B2(n_1127), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g1087 ( .A(n_41), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_42), .Y(n_1043) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_43), .A2(n_187), .B1(n_546), .B2(n_593), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_44), .A2(n_359), .B1(n_642), .B2(n_833), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_45), .B(n_914), .Y(n_1002) );
AOI222xp33_ASAP7_75t_L g894 ( .A1(n_46), .A2(n_207), .B1(n_305), .B2(n_546), .C1(n_630), .C2(n_895), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_47), .A2(n_311), .B1(n_566), .B2(n_909), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_48), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_49), .A2(n_323), .B1(n_614), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_50), .A2(n_209), .B1(n_884), .B2(n_1082), .Y(n_1081) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_51), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_52), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_53), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_54), .A2(n_180), .B1(n_432), .B2(n_773), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1090 ( .A(n_55), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_56), .A2(n_363), .B1(n_428), .B2(n_613), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g747 ( .A1(n_57), .A2(n_289), .B1(n_508), .B2(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_SL g655 ( .A1(n_58), .A2(n_656), .B1(n_681), .B2(n_682), .Y(n_655) );
CKINVDCx16_ASAP7_75t_R g682 ( .A(n_58), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_59), .A2(n_200), .B1(n_569), .B2(n_619), .Y(n_984) );
INVx1_ASAP7_75t_L g572 ( .A(n_60), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g532 ( .A1(n_61), .A2(n_198), .B1(n_234), .B2(n_533), .C1(n_534), .C2(n_536), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_62), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_63), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_64), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_65), .A2(n_201), .B1(n_522), .B2(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_66), .A2(n_294), .B1(n_774), .B2(n_1130), .Y(n_1129) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_67), .A2(n_265), .B1(n_571), .B2(n_644), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_68), .A2(n_275), .B1(n_525), .B2(n_569), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_69), .A2(n_93), .B1(n_571), .B2(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_70), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_71), .A2(n_252), .B1(n_468), .B2(n_519), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_72), .A2(n_146), .B1(n_559), .B2(n_567), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_73), .Y(n_419) );
AOI22xp5_ASAP7_75t_SL g560 ( .A1(n_74), .A2(n_249), .B1(n_561), .B2(n_563), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_75), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_76), .A2(n_245), .B1(n_606), .B2(n_644), .Y(n_814) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_77), .A2(n_121), .B1(n_529), .B2(n_563), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_78), .A2(n_274), .B1(n_508), .B2(n_767), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_79), .A2(n_212), .B1(n_448), .B2(n_776), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_80), .A2(n_109), .B1(n_525), .B2(n_527), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g1022 ( .A(n_81), .Y(n_1022) );
AO22x2_ASAP7_75t_L g418 ( .A1(n_82), .A2(n_256), .B1(n_409), .B2(n_410), .Y(n_418) );
INVx1_ASAP7_75t_L g1068 ( .A(n_82), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_83), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_84), .A2(n_254), .B1(n_531), .B2(n_608), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_85), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_86), .A2(n_89), .B1(n_426), .B2(n_774), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_87), .A2(n_306), .B1(n_767), .B2(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_88), .A2(n_378), .B1(n_529), .B2(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_90), .Y(n_424) );
AOI22xp5_ASAP7_75t_SL g568 ( .A1(n_91), .A2(n_205), .B1(n_569), .B2(n_571), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_92), .A2(n_290), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI211xp5_ASAP7_75t_L g834 ( .A1(n_95), .A2(n_559), .B(n_835), .C(n_840), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_96), .A2(n_279), .B1(n_733), .B2(n_787), .Y(n_826) );
AOI222xp33_ASAP7_75t_L g732 ( .A1(n_97), .A2(n_226), .B1(n_237), .B2(n_533), .C1(n_536), .C2(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g1054 ( .A(n_98), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_99), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_100), .A2(n_188), .B1(n_486), .B2(n_521), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_102), .A2(n_194), .B1(n_637), .B2(n_638), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_103), .A2(n_169), .B1(n_467), .B2(n_519), .Y(n_954) );
INVx1_ASAP7_75t_L g1072 ( .A(n_104), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_105), .A2(n_248), .B1(n_530), .B2(n_620), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_106), .B(n_1092), .Y(n_1091) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_107), .Y(n_584) );
XOR2xp5_ASAP7_75t_L g719 ( .A(n_108), .B(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_110), .A2(n_328), .B1(n_519), .B2(n_521), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_111), .A2(n_190), .B1(n_672), .B2(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_112), .B(n_515), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_113), .A2(n_324), .B1(n_508), .B2(n_642), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_114), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_115), .A2(n_181), .B1(n_426), .B2(n_432), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_116), .A2(n_302), .B1(n_726), .B2(n_727), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g703 ( .A1(n_117), .A2(n_203), .B1(n_704), .B2(n_705), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_118), .A2(n_358), .B1(n_426), .B2(n_619), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_119), .A2(n_236), .B1(n_569), .B2(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_120), .A2(n_133), .B1(n_486), .B2(n_535), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_122), .A2(n_318), .B1(n_563), .B2(n_833), .Y(n_939) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_123), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_124), .A2(n_329), .B1(n_452), .B2(n_529), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_125), .A2(n_238), .B1(n_519), .B2(n_588), .Y(n_744) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_126), .A2(n_244), .B1(n_733), .B2(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_127), .A2(n_366), .B1(n_830), .B2(n_869), .Y(n_868) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_128), .A2(n_341), .B1(n_486), .B2(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_129), .A2(n_199), .B1(n_608), .B2(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_130), .A2(n_183), .B1(n_515), .B2(n_638), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_131), .A2(n_360), .B1(n_616), .B2(n_619), .Y(n_615) );
XNOR2x2_ASAP7_75t_L g901 ( .A(n_132), .B(n_902), .Y(n_901) );
OA22x2_ASAP7_75t_L g919 ( .A1(n_134), .A2(n_920), .B1(n_921), .B2(n_940), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_134), .Y(n_920) );
INVx1_ASAP7_75t_L g755 ( .A(n_135), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_136), .B(n_552), .Y(n_1026) );
AND2x6_ASAP7_75t_L g387 ( .A(n_137), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_137), .Y(n_1065) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_138), .A2(n_368), .B1(n_566), .B2(n_884), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_139), .A2(n_179), .B1(n_421), .B2(n_672), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_140), .B(n_1051), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_141), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_142), .B(n_514), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_143), .A2(n_346), .B1(n_644), .B2(n_722), .Y(n_1012) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_144), .B(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_145), .A2(n_264), .B1(n_629), .B2(n_630), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_147), .Y(n_510) );
AO22x1_ASAP7_75t_L g873 ( .A1(n_148), .A2(n_874), .B1(n_896), .B2(n_897), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_148), .Y(n_896) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_149), .A2(n_170), .B1(n_421), .B2(n_957), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_150), .Y(n_806) );
AOI222xp33_ASAP7_75t_L g913 ( .A1(n_151), .A2(n_202), .B1(n_335), .B2(n_485), .C1(n_629), .C2(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_153), .A2(n_229), .B1(n_515), .B2(n_701), .Y(n_827) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_154), .A2(n_246), .B1(n_409), .B2(n_413), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g1069 ( .A(n_154), .B(n_1070), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_155), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_156), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_157), .A2(n_168), .B1(n_448), .B2(n_889), .Y(n_1124) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_158), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g1029 ( .A1(n_159), .A2(n_283), .B1(n_404), .B2(n_618), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_160), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_161), .A2(n_173), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g829 ( .A1(n_162), .A2(n_263), .B1(n_722), .B2(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g1089 ( .A(n_165), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_166), .A2(n_197), .B1(n_421), .B2(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_167), .A2(n_175), .B1(n_555), .B2(n_664), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_171), .A2(n_258), .B1(n_428), .B2(n_529), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_172), .A2(n_182), .B1(n_637), .B2(n_638), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_174), .A2(n_314), .B1(n_608), .B2(n_610), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_176), .A2(n_304), .B1(n_619), .B2(n_773), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g875 ( .A1(n_177), .A2(n_196), .B1(n_678), .B2(n_774), .C(n_876), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_178), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_184), .Y(n_850) );
INVx1_ASAP7_75t_L g1106 ( .A(n_185), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_185), .A2(n_1106), .B1(n_1108), .B2(n_1131), .Y(n_1107) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_186), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_189), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_191), .B(n_550), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_193), .A2(n_247), .B1(n_428), .B2(n_613), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_195), .A2(n_291), .B1(n_452), .B2(n_865), .Y(n_864) );
XNOR2xp5_ASAP7_75t_L g819 ( .A(n_204), .B(n_820), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_206), .A2(n_235), .B1(n_527), .B2(n_1008), .Y(n_1007) );
AOI22xp33_ASAP7_75t_SL g1009 ( .A1(n_208), .A2(n_228), .B1(n_563), .B2(n_752), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_210), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_211), .A2(n_231), .B1(n_674), .B2(n_884), .C(n_885), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_213), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_214), .A2(n_338), .B1(n_865), .B2(n_889), .Y(n_1083) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_216), .B(n_514), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_217), .A2(n_317), .B1(n_433), .B2(n_504), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_218), .A2(n_351), .B1(n_486), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_219), .A2(n_260), .B1(n_679), .B2(n_754), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g981 ( .A1(n_221), .A2(n_296), .B1(n_452), .B2(n_982), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_222), .B(n_610), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_223), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_224), .A2(n_357), .B1(n_674), .B2(n_675), .Y(n_673) );
OA22x2_ASAP7_75t_L g992 ( .A1(n_225), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_225), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_227), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_230), .A2(n_250), .B1(n_506), .B2(n_508), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_232), .A2(n_321), .B1(n_504), .B2(n_774), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_233), .Y(n_1042) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_239), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_240), .Y(n_544) );
INVx2_ASAP7_75t_L g391 ( .A(n_242), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_243), .A2(n_288), .B1(n_508), .B2(n_754), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_251), .A2(n_278), .B1(n_556), .B2(n_634), .Y(n_1053) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_253), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_255), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_259), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g977 ( .A(n_262), .Y(n_977) );
OA22x2_ASAP7_75t_L g621 ( .A1(n_267), .A2(n_622), .B1(n_623), .B2(n_648), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_267), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g612 ( .A1(n_269), .A2(n_286), .B1(n_613), .B2(n_614), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_270), .Y(n_457) );
AOI22x1_ASAP7_75t_L g844 ( .A1(n_271), .A2(n_845), .B1(n_871), .B2(n_872), .Y(n_844) );
INVx1_ASAP7_75t_L g871 ( .A(n_271), .Y(n_871) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_272), .A2(n_383), .B(n_392), .C(n_1073), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_273), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_276), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_277), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g409 ( .A(n_280), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_280), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_281), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_284), .B(n_637), .Y(n_1052) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_285), .A2(n_322), .B1(n_421), .B2(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_287), .A2(n_367), .B1(n_672), .B2(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_293), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g1086 ( .A(n_295), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_297), .A2(n_692), .B1(n_693), .B2(n_716), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_297), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_298), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_299), .A2(n_319), .B1(n_404), .B2(n_773), .Y(n_1123) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_300), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g1094 ( .A(n_301), .Y(n_1094) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_303), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g1116 ( .A(n_307), .Y(n_1116) );
INVx1_ASAP7_75t_L g390 ( .A(n_308), .Y(n_390) );
INVx1_ASAP7_75t_L g1120 ( .A(n_309), .Y(n_1120) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_310), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g970 ( .A(n_312), .Y(n_970) );
INVx1_ASAP7_75t_L g388 ( .A(n_313), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_315), .Y(n_797) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_320), .A2(n_365), .B1(n_678), .B2(n_679), .Y(n_677) );
XOR2x2_ASAP7_75t_L g960 ( .A(n_325), .B(n_961), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g937 ( .A1(n_327), .A2(n_333), .B1(n_571), .B2(n_938), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_330), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_332), .B(n_726), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_336), .A2(n_1075), .B1(n_1096), .B2(n_1097), .Y(n_1074) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_336), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_337), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_339), .A2(n_373), .B1(n_521), .B2(n_594), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_340), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_342), .B(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_343), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_345), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_347), .A2(n_354), .B1(n_485), .B2(n_535), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_348), .A2(n_361), .B1(n_571), .B2(n_909), .Y(n_908) );
XNOR2x1_ASAP7_75t_L g793 ( .A(n_349), .B(n_794), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_350), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_352), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_353), .A2(n_376), .B1(n_529), .B2(n_610), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_355), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_356), .B(n_552), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_362), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_364), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_369), .B(n_631), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_370), .B(n_535), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_371), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_372), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_374), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g1111 ( .A(n_375), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_377), .B(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_380), .Y(n_1114) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_384), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_388), .Y(n_1064) );
OAI21xp5_ASAP7_75t_L g1104 ( .A1(n_389), .A2(n_1063), .B(n_1105), .Y(n_1104) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_816), .B1(n_1058), .B2(n_1059), .C(n_1060), .Y(n_392) );
INVx1_ASAP7_75t_L g1058 ( .A(n_393), .Y(n_1058) );
XOR2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_651), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B1(n_574), .B2(n_575), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_497), .B1(n_498), .B2(n_573), .Y(n_397) );
INVx2_ASAP7_75t_L g573 ( .A(n_398), .Y(n_573) );
INVx1_ASAP7_75t_L g495 ( .A(n_399), .Y(n_495) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_400), .B(n_455), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_437), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_419), .B1(n_420), .B2(n_424), .C(n_425), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g503 ( .A(n_403), .Y(n_503) );
INVx5_ASAP7_75t_SL g613 ( .A(n_403), .Y(n_613) );
INVx4_ASAP7_75t_L g909 ( .A(n_403), .Y(n_909) );
INVx2_ASAP7_75t_SL g957 ( .A(n_403), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_403), .A2(n_526), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
INVx11_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx11_ASAP7_75t_L g570 ( .A(n_404), .Y(n_570) );
AND2x6_ASAP7_75t_L g404 ( .A(n_405), .B(n_414), .Y(n_404) );
AND2x4_ASAP7_75t_L g517 ( .A(n_405), .B(n_440), .Y(n_517) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_412), .Y(n_406) );
AND2x2_ASAP7_75t_L g423 ( .A(n_407), .B(n_412), .Y(n_423) );
AND2x2_ASAP7_75t_L g430 ( .A(n_407), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g471 ( .A(n_408), .B(n_416), .Y(n_471) );
AND2x2_ASAP7_75t_L g475 ( .A(n_408), .B(n_412), .Y(n_475) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_411), .Y(n_413) );
INVx2_ASAP7_75t_L g431 ( .A(n_412), .Y(n_431) );
INVx1_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
AND2x4_ASAP7_75t_L g422 ( .A(n_414), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g429 ( .A(n_414), .B(n_430), .Y(n_429) );
AND2x6_ASAP7_75t_L g474 ( .A(n_414), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
AND2x2_ASAP7_75t_L g440 ( .A(n_415), .B(n_418), .Y(n_440) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g435 ( .A(n_416), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_416), .B(n_418), .Y(n_445) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g436 ( .A(n_418), .Y(n_436) );
INVx1_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx6_ASAP7_75t_L g526 ( .A(n_422), .Y(n_526) );
BUFx3_ASAP7_75t_L g606 ( .A(n_422), .Y(n_606) );
BUFx3_ASAP7_75t_L g722 ( .A(n_422), .Y(n_722) );
AND2x2_ASAP7_75t_L g451 ( .A(n_423), .B(n_435), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g464 ( .A(n_423), .B(n_440), .Y(n_464) );
AND2x6_ASAP7_75t_L g552 ( .A(n_423), .B(n_440), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g838 ( .A(n_423), .B(n_435), .Y(n_838) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_427), .A2(n_1042), .B1(n_1043), .B2(n_1044), .Y(n_1041) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g605 ( .A(n_428), .Y(n_605) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_428), .Y(n_714) );
BUFx3_ASAP7_75t_L g773 ( .A(n_428), .Y(n_773) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g507 ( .A(n_429), .Y(n_507) );
BUFx2_ASAP7_75t_SL g559 ( .A(n_429), .Y(n_559) );
BUFx2_ASAP7_75t_SL g678 ( .A(n_429), .Y(n_678) );
AND2x2_ASAP7_75t_L g434 ( .A(n_430), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g439 ( .A(n_430), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g443 ( .A(n_430), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_430), .B(n_435), .Y(n_882) );
AND2x2_ASAP7_75t_L g469 ( .A(n_431), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g480 ( .A(n_431), .Y(n_480) );
BUFx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g508 ( .A(n_434), .Y(n_508) );
BUFx3_ASAP7_75t_L g566 ( .A(n_434), .Y(n_566) );
BUFx3_ASAP7_75t_L g618 ( .A(n_434), .Y(n_618) );
INVx1_ASAP7_75t_L g494 ( .A(n_436), .Y(n_494) );
OAI221xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_441), .B1(n_442), .B2(n_446), .C(n_447), .Y(n_437) );
INVx2_ASAP7_75t_L g1082 ( .A(n_438), .Y(n_1082) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g527 ( .A(n_439), .Y(n_527) );
BUFx3_ASAP7_75t_L g620 ( .A(n_439), .Y(n_620) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_439), .Y(n_679) );
BUFx3_ASAP7_75t_L g833 ( .A(n_439), .Y(n_833) );
INVx1_ASAP7_75t_L g461 ( .A(n_440), .Y(n_461) );
INVx1_ASAP7_75t_L g767 ( .A(n_442), .Y(n_767) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g504 ( .A(n_443), .Y(n_504) );
BUFx2_ASAP7_75t_L g567 ( .A(n_443), .Y(n_567) );
BUFx2_ASAP7_75t_SL g614 ( .A(n_443), .Y(n_614) );
BUFx2_ASAP7_75t_SL g642 ( .A(n_443), .Y(n_642) );
BUFx3_ASAP7_75t_L g748 ( .A(n_443), .Y(n_748) );
BUFx3_ASAP7_75t_L g884 ( .A(n_443), .Y(n_884) );
AND2x2_ASAP7_75t_L g754 ( .A(n_444), .B(n_480), .Y(n_754) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x6_ASAP7_75t_L g453 ( .A(n_445), .B(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g529 ( .A(n_450), .Y(n_529) );
INVx4_ASAP7_75t_L g562 ( .A(n_450), .Y(n_562) );
INVx5_ASAP7_75t_L g752 ( .A(n_450), .Y(n_752) );
INVx1_ASAP7_75t_L g938 ( .A(n_450), .Y(n_938) );
INVx8_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx6_ASAP7_75t_SL g531 ( .A(n_453), .Y(n_531) );
INVx1_ASAP7_75t_SL g610 ( .A(n_453), .Y(n_610) );
INVx1_ASAP7_75t_SL g776 ( .A(n_453), .Y(n_776) );
INVx1_ASAP7_75t_L g520 ( .A(n_454), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .C(n_482), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_462), .B2(n_463), .Y(n_456) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g965 ( .A(n_459), .Y(n_965) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_460), .Y(n_582) );
BUFx3_ASAP7_75t_L g798 ( .A(n_460), .Y(n_798) );
OAI22xp5_ASAP7_75t_SL g581 ( .A1(n_463), .A2(n_582), .B1(n_583), .B2(n_584), .Y(n_581) );
BUFx3_ASAP7_75t_L g800 ( .A(n_463), .Y(n_800) );
INVx2_ASAP7_75t_L g968 ( .A(n_463), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_463), .A2(n_798), .B1(n_998), .B2(n_999), .Y(n_997) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g512 ( .A(n_464), .Y(n_512) );
OAI222xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_472), .B1(n_473), .B2(n_476), .C1(n_477), .C2(n_481), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g781 ( .A(n_467), .Y(n_781) );
BUFx4f_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_468), .Y(n_535) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_468), .Y(n_588) );
BUFx2_ASAP7_75t_L g629 ( .A(n_468), .Y(n_629) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_468), .Y(n_664) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g488 ( .A(n_470), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_471), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g487 ( .A(n_471), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g519 ( .A(n_471), .B(n_520), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_473), .A2(n_738), .B(n_739), .Y(n_737) );
OAI21xp33_ASAP7_75t_SL g801 ( .A1(n_473), .A2(n_802), .B(n_803), .Y(n_801) );
OAI221xp5_ASAP7_75t_L g847 ( .A1(n_473), .A2(n_848), .B1(n_849), .B2(n_850), .C(n_851), .Y(n_847) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_473), .A2(n_970), .B1(n_971), .B2(n_972), .C(n_973), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g1113 ( .A1(n_473), .A2(n_1114), .B1(n_1115), .B2(n_1116), .C(n_1117), .Y(n_1113) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_474), .Y(n_533) );
INVx4_ASAP7_75t_L g543 ( .A(n_474), .Y(n_543) );
INVx2_ASAP7_75t_SL g590 ( .A(n_474), .Y(n_590) );
INVx2_ASAP7_75t_L g626 ( .A(n_474), .Y(n_626) );
BUFx3_ASAP7_75t_L g914 ( .A(n_474), .Y(n_914) );
INVx1_ASAP7_75t_L g492 ( .A(n_475), .Y(n_492) );
AND2x4_ASAP7_75t_L g522 ( .A(n_475), .B(n_494), .Y(n_522) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_SL g667 ( .A(n_478), .Y(n_667) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g597 ( .A(n_479), .Y(n_597) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_479), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_479), .A2(n_491), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_489), .B2(n_490), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx4f_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_487), .Y(n_594) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_487), .Y(n_631) );
INVx1_ASAP7_75t_L g783 ( .A(n_487), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_490), .A2(n_667), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g600 ( .A(n_491), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_491), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_665) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
XNOR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_539), .Y(n_498) );
AO22x1_ASAP7_75t_L g654 ( .A1(n_499), .A2(n_655), .B1(n_683), .B2(n_684), .Y(n_654) );
INVx1_ASAP7_75t_L g684 ( .A(n_499), .Y(n_684) );
XOR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_538), .Y(n_499) );
NAND4xp75_ASAP7_75t_L g500 ( .A(n_501), .B(n_509), .C(n_523), .D(n_532), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g1008 ( .A(n_507), .Y(n_1008) );
OA211x2_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_513), .C(n_518), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_511), .A2(n_582), .B1(n_659), .B2(n_660), .Y(n_658) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g855 ( .A(n_512), .Y(n_855) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx5_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g637 ( .A(n_516), .Y(n_637) );
INVx2_ASAP7_75t_L g726 ( .A(n_516), .Y(n_726) );
INVx2_ASAP7_75t_L g742 ( .A(n_516), .Y(n_742) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
INVx1_ASAP7_75t_L g635 ( .A(n_519), .Y(n_635) );
BUFx2_ASAP7_75t_L g787 ( .A(n_519), .Y(n_787) );
BUFx2_ASAP7_75t_L g927 ( .A(n_519), .Y(n_927) );
INVx1_ASAP7_75t_SL g706 ( .A(n_521), .Y(n_706) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx2_ASAP7_75t_SL g556 ( .A(n_522), .Y(n_556) );
BUFx3_ASAP7_75t_L g733 ( .A(n_522), .Y(n_733) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .Y(n_523) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g571 ( .A(n_526), .Y(n_571) );
INVx2_ASAP7_75t_L g675 ( .A(n_526), .Y(n_675) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g563 ( .A(n_531), .Y(n_563) );
BUFx4f_ASAP7_75t_SL g889 ( .A(n_531), .Y(n_889) );
INVx2_ASAP7_75t_L g696 ( .A(n_533), .Y(n_696) );
INVx2_ASAP7_75t_SL g779 ( .A(n_533), .Y(n_779) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g547 ( .A(n_535), .Y(n_547) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
XOR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_572), .Y(n_539) );
NAND3x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_557), .C(n_564), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_544), .B(n_545), .Y(n_542) );
INVx4_ASAP7_75t_L g895 ( .A(n_543), .Y(n_895) );
BUFx2_ASAP7_75t_L g929 ( .A(n_543), .Y(n_929) );
OAI21xp5_ASAP7_75t_L g948 ( .A1(n_543), .A2(n_949), .B(n_950), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g1021 ( .A1(n_543), .A2(n_1022), .B(n_1023), .Y(n_1021) );
OAI21xp5_ASAP7_75t_SL g1046 ( .A1(n_543), .A2(n_1047), .B(n_1048), .Y(n_1046) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .C(n_554), .Y(n_548) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_SL g638 ( .A(n_551), .Y(n_638) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g701 ( .A(n_552), .Y(n_701) );
BUFx4f_ASAP7_75t_L g727 ( .A(n_552), .Y(n_727) );
BUFx2_ASAP7_75t_L g1051 ( .A(n_552), .Y(n_1051) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g609 ( .A(n_562), .Y(n_609) );
BUFx6f_ASAP7_75t_L g982 ( .A(n_562), .Y(n_982) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
BUFx2_ASAP7_75t_L g830 ( .A(n_566), .Y(n_830) );
INVx1_ASAP7_75t_L g1128 ( .A(n_566), .Y(n_1128) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g644 ( .A(n_570), .Y(n_644) );
INVx3_ASAP7_75t_L g674 ( .A(n_570), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_570), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_621), .B1(n_649), .B2(n_650), .Y(n_576) );
INVx2_ASAP7_75t_L g649 ( .A(n_577), .Y(n_649) );
XNOR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_602), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_585), .C(n_596), .Y(n_580) );
OAI222xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_589), .B1(n_590), .B2(n_591), .C1(n_592), .C2(n_595), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_SL g1115 ( .A(n_587), .Y(n_1115) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI21xp5_ASAP7_75t_SL g661 ( .A1(n_590), .A2(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx4f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI22xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_598), .B1(n_599), .B2(n_601), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_597), .A2(n_807), .B1(n_892), .B2(n_893), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_599), .A2(n_975), .B1(n_976), .B2(n_977), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_599), .A2(n_667), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g807 ( .A(n_600), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_611), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g870 ( .A(n_606), .Y(n_870) );
INVx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_615), .Y(n_611) );
INVx1_ASAP7_75t_L g770 ( .A(n_613), .Y(n_770) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx4f_ASAP7_75t_SL g672 ( .A(n_618), .Y(n_672) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g650 ( .A(n_621), .Y(n_650) );
INVx2_ASAP7_75t_L g648 ( .A(n_623), .Y(n_648) );
NAND2x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_639), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_632), .Y(n_624) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_627), .B(n_628), .Y(n_625) );
INVx2_ASAP7_75t_L g971 ( .A(n_630), .Y(n_971) );
BUFx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_631), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_636), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g704 ( .A(n_635), .Y(n_704) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_645), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AOI22xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_758), .B1(n_759), .B2(n_815), .Y(n_651) );
INVx1_ASAP7_75t_L g815 ( .A(n_652), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_685), .B2(n_686), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g683 ( .A(n_655), .Y(n_683) );
INVx2_ASAP7_75t_L g681 ( .A(n_656), .Y(n_681) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_669), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .C(n_665), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_664), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_667), .A2(n_805), .B1(n_806), .B2(n_807), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_667), .A2(n_807), .B1(n_857), .B2(n_858), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_676), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx2_ASAP7_75t_L g878 ( .A(n_675), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .Y(n_676) );
INVx4_ASAP7_75t_L g710 ( .A(n_679), .Y(n_710) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_717), .B2(n_718), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g716 ( .A(n_693), .Y(n_716) );
NAND3x1_ASAP7_75t_L g693 ( .A(n_694), .B(n_707), .C(n_712), .Y(n_693) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_699), .Y(n_694) );
OAI21xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_697), .B(n_698), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g822 ( .A1(n_696), .A2(n_823), .B(n_824), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .C(n_703), .Y(n_699) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx4_ASAP7_75t_L g774 ( .A(n_710), .Y(n_774) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AO22x2_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_734), .B1(n_756), .B2(n_757), .Y(n_718) );
INVx1_ASAP7_75t_L g756 ( .A(n_719), .Y(n_756) );
NAND5xp2_ASAP7_75t_SL g720 ( .A(n_721), .B(n_723), .C(n_724), .D(n_729), .E(n_732), .Y(n_720) );
AND2x2_ASAP7_75t_SL g724 ( .A(n_725), .B(n_728), .Y(n_724) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx2_ASAP7_75t_L g757 ( .A(n_734), .Y(n_757) );
XOR2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_755), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g735 ( .A(n_736), .B(n_745), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .C(n_744), .Y(n_740) );
NOR2x1_ASAP7_75t_L g745 ( .A(n_746), .B(n_750), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_749), .Y(n_746) );
INVx2_ASAP7_75t_L g863 ( .A(n_748), .Y(n_863) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_748), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .Y(n_750) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_752), .Y(n_865) );
INVx3_ASAP7_75t_L g792 ( .A(n_757), .Y(n_792) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_790), .B2(n_791), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g789 ( .A(n_763), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_777), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_771), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_785), .Y(n_777) );
OAI222xp33_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B1(n_781), .B2(n_782), .C1(n_783), .C2(n_784), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
XNOR2x1_ASAP7_75t_SL g791 ( .A(n_792), .B(n_793), .Y(n_791) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_808), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_801), .C(n_804), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_798), .A2(n_853), .B1(n_854), .B2(n_855), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_798), .A2(n_855), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_798), .A2(n_967), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g1059 ( .A(n_816), .Y(n_1059) );
XOR2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_990), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B1(n_842), .B2(n_989), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND3x1_ASAP7_75t_L g820 ( .A(n_821), .B(n_828), .C(n_834), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_825), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
BUFx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
OAI21xp33_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B(n_839), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_837), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
BUFx2_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g989 ( .A(n_842), .Y(n_989) );
XNOR2x1_ASAP7_75t_L g842 ( .A(n_843), .B(n_900), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_873), .B1(n_898), .B2(n_899), .Y(n_843) );
INVx1_ASAP7_75t_L g898 ( .A(n_844), .Y(n_898) );
INVx2_ASAP7_75t_SL g872 ( .A(n_845), .Y(n_872) );
AND2x4_ASAP7_75t_L g845 ( .A(n_846), .B(n_859), .Y(n_845) );
NOR3xp33_ASAP7_75t_SL g846 ( .A(n_847), .B(n_852), .C(n_856), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_849), .A2(n_929), .B1(n_1089), .B2(n_1090), .C(n_1091), .Y(n_1088) );
NOR2x1_ASAP7_75t_L g859 ( .A(n_860), .B(n_866), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .Y(n_860) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g899 ( .A(n_873), .Y(n_899) );
INVx1_ASAP7_75t_L g897 ( .A(n_874), .Y(n_897) );
AND4x1_ASAP7_75t_L g874 ( .A(n_875), .B(n_883), .C(n_890), .D(n_894), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_876) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1044 ( .A(n_881), .Y(n_1044) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_889), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_915), .B1(n_987), .B2(n_988), .Y(n_900) );
INVx2_ASAP7_75t_L g987 ( .A(n_901), .Y(n_987) );
NAND4xp75_ASAP7_75t_L g902 ( .A(n_903), .B(n_906), .C(n_910), .D(n_913), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .Y(n_903) );
AND2x2_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
AND2x2_ASAP7_75t_SL g910 ( .A(n_911), .B(n_912), .Y(n_910) );
INVx1_ASAP7_75t_L g988 ( .A(n_915), .Y(n_988) );
AOI22xp5_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_917), .B1(n_960), .B2(n_986), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
OAI22xp5_ASAP7_75t_SL g917 ( .A1(n_918), .A2(n_919), .B1(n_941), .B2(n_942), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx2_ASAP7_75t_SL g940 ( .A(n_921), .Y(n_940) );
NAND2x1p5_ASAP7_75t_L g921 ( .A(n_922), .B(n_932), .Y(n_921) );
NOR2xp67_ASAP7_75t_SL g922 ( .A(n_923), .B(n_928), .Y(n_922) );
NAND3xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .C(n_926), .Y(n_923) );
OAI21xp5_ASAP7_75t_SL g928 ( .A1(n_929), .A2(n_930), .B(n_931), .Y(n_928) );
NOR2x1_ASAP7_75t_L g932 ( .A(n_933), .B(n_936), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_939), .Y(n_936) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
XOR2x2_ASAP7_75t_L g942 ( .A(n_943), .B(n_959), .Y(n_942) );
NAND3x1_ASAP7_75t_L g943 ( .A(n_944), .B(n_947), .C(n_955), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
NOR2x1_ASAP7_75t_L g947 ( .A(n_948), .B(n_951), .Y(n_947) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .C(n_954), .Y(n_951) );
AND2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_958), .Y(n_955) );
INVx2_ASAP7_75t_L g986 ( .A(n_960), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_978), .Y(n_961) );
NOR3xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_969), .C(n_974), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_965), .B1(n_966), .B2(n_967), .Y(n_963) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_979), .B(n_983), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_981), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_985), .Y(n_983) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_1013), .B1(n_1056), .B2(n_1057), .Y(n_991) );
INVx2_ASAP7_75t_SL g1056 ( .A(n_992), .Y(n_1056) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
AND3x1_ASAP7_75t_L g995 ( .A(n_996), .B(n_1006), .C(n_1010), .Y(n_995) );
NOR3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_1000), .C(n_1003), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1009), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1013), .Y(n_1057) );
OA22x2_ASAP7_75t_L g1013 ( .A1(n_1014), .A2(n_1015), .B1(n_1032), .B2(n_1055), .Y(n_1013) );
INVx3_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
XOR2x2_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1031), .Y(n_1015) );
NAND3x1_ASAP7_75t_SL g1016 ( .A(n_1017), .B(n_1020), .C(n_1028), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
NOR2x1_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1024), .Y(n_1020) );
NAND3xp33_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1026), .C(n_1027), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1030), .Y(n_1028) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1032), .Y(n_1055) );
XOR2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1054), .Y(n_1032) );
AND2x2_ASAP7_75t_SL g1033 ( .A(n_1034), .B(n_1045), .Y(n_1033) );
NOR3xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1038), .C(n_1041), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1049), .Y(n_1045) );
NAND3xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1052), .C(n_1053), .Y(n_1049) );
INVx1_ASAP7_75t_SL g1060 ( .A(n_1061), .Y(n_1060) );
NOR2x1_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1066), .Y(n_1061) );
OR2x2_ASAP7_75t_SL g1134 ( .A(n_1062), .B(n_1067), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1065), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_1063), .Y(n_1100) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1064), .B(n_1102), .Y(n_1105) );
CKINVDCx16_ASAP7_75t_R g1102 ( .A(n_1065), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g1066 ( .A(n_1067), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1069), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1072), .Y(n_1070) );
OAI322xp33_ASAP7_75t_L g1073 ( .A1(n_1074), .A2(n_1098), .A3(n_1101), .B1(n_1103), .B2(n_1106), .C1(n_1107), .C2(n_1132), .Y(n_1073) );
INVx1_ASAP7_75t_SL g1097 ( .A(n_1075), .Y(n_1097) );
AND2x2_ASAP7_75t_SL g1075 ( .A(n_1076), .B(n_1084), .Y(n_1075) );
NOR2xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1080), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1079), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1083), .Y(n_1080) );
NOR3xp33_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1088), .C(n_1093), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
CKINVDCx16_ASAP7_75t_R g1103 ( .A(n_1104), .Y(n_1103) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1108), .Y(n_1131) );
AND2x2_ASAP7_75t_SL g1108 ( .A(n_1109), .B(n_1121), .Y(n_1108) );
NOR3xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1113), .C(n_1118), .Y(n_1109) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1125), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1124), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1129), .Y(n_1125) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
CKINVDCx20_ASAP7_75t_R g1132 ( .A(n_1133), .Y(n_1132) );
CKINVDCx20_ASAP7_75t_R g1133 ( .A(n_1134), .Y(n_1133) );
endmodule