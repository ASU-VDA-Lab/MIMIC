module real_jpeg_4631_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_0),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_0),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_0),
.B(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_0),
.B(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_2),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_2),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_2),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_2),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_2),
.B(n_66),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_2),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_3),
.B(n_27),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_3),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_3),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_3),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_3),
.B(n_213),
.Y(n_421)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_4),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_4),
.Y(n_273)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_6),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_6),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_6),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_6),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_6),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_7),
.Y(n_203)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_7),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_7),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_7),
.Y(n_393)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_8),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_8),
.Y(n_395)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_11),
.B(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_11),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_11),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_11),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_11),
.B(n_335),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_11),
.A2(n_390),
.B(n_395),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_12),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_13),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_13),
.B(n_94),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_13),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_13),
.B(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_13),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_13),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_13),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_14),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_14),
.B(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_14),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_14),
.B(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_14),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_14),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_15),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_15),
.B(n_27),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_15),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_15),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_15),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_15),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_15),
.B(n_304),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_470),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_219),
.B(n_467),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_174),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_SL g467 ( 
.A1(n_19),
.A2(n_468),
.B(n_469),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_137),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_20),
.B(n_137),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_21),
.B(n_103),
.C(n_119),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_68),
.C(n_81),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_22),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_50),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_23),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_26),
.B(n_35),
.C(n_38),
.Y(n_105)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_29),
.A2(n_35),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_29),
.A2(n_35),
.B1(n_198),
.B2(n_199),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_29),
.B(n_199),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_32),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_33),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_33),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_40),
.C(n_45),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_36),
.A2(n_38),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_36),
.A2(n_38),
.B1(n_343),
.B2(n_347),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_36),
.B(n_343),
.C(n_348),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_38),
.B(n_108),
.C(n_115),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_39),
.B(n_50),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_40),
.A2(n_123),
.B1(n_124),
.B2(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_40),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_40),
.A2(n_45),
.B1(n_129),
.B2(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_44),
.Y(n_150)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_45),
.Y(n_146)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_49),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_49),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_64),
.B2(n_65),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_55),
.Y(n_238)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_56),
.Y(n_316)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_57),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_57),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_58),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_62),
.C(n_65),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_58),
.B(n_188),
.Y(n_414)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_63),
.B(n_187),
.C(n_189),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_64),
.A2(n_65),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_68),
.A2(n_81),
.B1(n_82),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_76),
.C(n_79),
.Y(n_121)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_71),
.B(n_257),
.Y(n_389)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_74),
.B(n_85),
.C(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_74),
.A2(n_79),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_78),
.Y(n_320)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_93),
.C(n_98),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_83),
.A2(n_84),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.C(n_91),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_85),
.A2(n_91),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_85),
.A2(n_157),
.B1(n_163),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_85),
.A2(n_157),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_85),
.B(n_253),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_87),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_87),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_87),
.A2(n_159),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_87),
.B(n_399),
.C(n_402),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_89),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_90),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_91),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_93),
.A2(n_98),
.B1(n_99),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_97),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_98),
.A2(n_99),
.B1(n_166),
.B2(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_162),
.C(n_166),
.Y(n_161)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_119),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_138),
.C(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_103),
.B(n_138),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_105),
.CI(n_106),
.CON(n_103),
.SN(n_103)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_108),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_107),
.A2(n_108),
.B1(n_376),
.B2(n_380),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_107),
.B(n_369),
.C(n_380),
.Y(n_415)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_108),
.B(n_125),
.C(n_129),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_127),
.Y(n_126)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_112),
.Y(n_312)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_117),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_121),
.B(n_122),
.C(n_130),
.Y(n_474)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_125),
.A2(n_126),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_125),
.A2(n_126),
.B1(n_148),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_126),
.B(n_198),
.C(n_204),
.Y(n_197)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_127),
.Y(n_346)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_131),
.B(n_134),
.C(n_135),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_133),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_141),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_161),
.C(n_170),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_155),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_143),
.B(n_147),
.Y(n_438)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_154),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_148),
.Y(n_481)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_SL g335 ( 
.A(n_150),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_154),
.Y(n_195)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_155),
.B(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_170),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_163),
.A2(n_185),
.B1(n_355),
.B2(n_356),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_163),
.B(n_355),
.Y(n_383)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_217),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_175),
.B(n_217),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_176),
.B(n_178),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_180),
.B(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_196),
.C(n_214),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g439 ( 
.A(n_181),
.B(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_194),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_182),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_186),
.B(n_194),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_189),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_196),
.B(n_214),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_206),
.C(n_209),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_197),
.B(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_198),
.A2(n_199),
.B1(n_204),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_203),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_204),
.Y(n_432)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_205),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_206),
.Y(n_424)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_407),
.B1(n_460),
.B2(n_465),
.C(n_466),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_362),
.B(n_406),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_323),
.B(n_361),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_298),
.B(n_322),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_265),
.B(n_297),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_254),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_225),
.B(n_254),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_239),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_226),
.B(n_240),
.C(n_251),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_227),
.B(n_232),
.C(n_236),
.Y(n_308)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_251),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_246),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_242),
.B(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.C(n_261),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_256),
.A2(n_261),
.B1(n_262),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_291),
.B(n_296),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_281),
.B(n_290),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_278),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_274),
.Y(n_292)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_286),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_300),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_307),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_308),
.C(n_309),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_305),
.C(n_306),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_314),
.C(n_321),
.Y(n_357)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_317),
.B2(n_321),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_360),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_360),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_340),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_329),
.C(n_340),
.Y(n_363)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_329)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_336),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_336),
.C(n_337),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_353),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_357),
.C(n_359),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_348),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_353)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_364),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_386),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_366),
.B(n_367),
.C(n_386),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_381),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_382),
.C(n_385),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_375),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_405),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_396),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_396),
.C(n_405),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B(n_394),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_420),
.C(n_421),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_442),
.C(n_446),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_408),
.A2(n_461),
.B(n_464),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_435),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_409),
.B(n_435),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_425),
.C(n_427),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_425),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_418),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_419),
.C(n_422),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.C(n_416),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_417),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_421),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.C(n_433),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_433),
.Y(n_450)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_441),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_439),
.C(n_441),
.Y(n_445)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_445),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_456),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_447),
.A2(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_454),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_454),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_451),
.C(n_452),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_452),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_458),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_490),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_473),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_482),
.B1(n_483),
.B2(n_489),
.Y(n_477)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_478),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_484),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_485),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_487),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);


endmodule