module fake_jpeg_17182_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_46),
.B1(n_43),
.B2(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_81),
.Y(n_100)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_43),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_90),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_44),
.B1(n_54),
.B2(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_92),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_70),
.B1(n_69),
.B2(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_52),
.B1(n_49),
.B2(n_48),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_96),
.B1(n_101),
.B2(n_8),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_51),
.B1(n_55),
.B2(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_17),
.B1(n_36),
.B2(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_0),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_110),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_108),
.A3(n_96),
.B1(n_94),
.B2(n_9),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_85),
.B1(n_92),
.B2(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_105),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_117),
.B1(n_104),
.B2(n_112),
.Y(n_125)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVxp33_ASAP7_75t_SL g121 ( 
.A(n_120),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_125),
.B1(n_119),
.B2(n_112),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_131),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_89),
.B1(n_88),
.B2(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_136),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_118),
.C(n_84),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_118),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_24),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_138),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_141),
.C(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_132),
.B(n_10),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_25),
.C(n_11),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_26),
.C(n_12),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_148),
.A2(n_37),
.B(n_14),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_27),
.B(n_15),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_30),
.B(n_16),
.Y(n_152)
);


endmodule