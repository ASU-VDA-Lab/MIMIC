module fake_netlist_5_363_n_47 (n_8, n_10, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_11, n_6, n_1, n_47);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_11;
input n_6;
input n_1;

output n_47;

wire n_29;
wire n_16;
wire n_43;
wire n_12;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_42;
wire n_22;
wire n_45;
wire n_28;
wire n_24;
wire n_46;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_38;
wire n_32;
wire n_35;
wire n_41;
wire n_17;
wire n_19;
wire n_37;
wire n_26;
wire n_15;
wire n_30;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_20;
wire n_39;

AOI22xp5_ASAP7_75t_L g12 ( 
.A1(n_8),
.A2(n_1),
.B1(n_7),
.B2(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_3),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_4),
.A2(n_9),
.B1(n_11),
.B2(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AND2x4_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_2),
.Y(n_19)
);

AND2x4_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_21),
.C(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_17),
.B(n_14),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_17),
.B(n_20),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_20),
.B1(n_19),
.B2(n_13),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_24),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_29),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_24),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_33),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_37),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_15),
.Y(n_42)
);

XNOR2x1_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_12),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_43),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_22),
.B1(n_19),
.B2(n_34),
.Y(n_47)
);


endmodule