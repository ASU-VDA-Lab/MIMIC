module fake_jpeg_8171_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_22),
.B1(n_27),
.B2(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_16),
.B1(n_25),
.B2(n_37),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_49),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_16),
.B1(n_23),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_23),
.B1(n_21),
.B2(n_32),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_23),
.B1(n_29),
.B2(n_32),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_21),
.B1(n_34),
.B2(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_61),
.B1(n_18),
.B2(n_24),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_18),
.B1(n_34),
.B2(n_31),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_28),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_75),
.B(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_83),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_36),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_77),
.B(n_108),
.C(n_78),
.Y(n_126)
);

NAND2x1_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_46),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_78),
.A2(n_98),
.B(n_90),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_79),
.Y(n_127)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_19),
.B1(n_22),
.B2(n_27),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_19),
.B1(n_22),
.B2(n_27),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_31),
.B1(n_24),
.B2(n_18),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_45),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_95),
.C(n_97),
.Y(n_132)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_24),
.B1(n_53),
.B2(n_64),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_42),
.C(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_42),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_52),
.B(n_31),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_14),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_51),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_42),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_46),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_78),
.C(n_101),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_95),
.B1(n_103),
.B2(n_108),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_137),
.B(n_94),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_76),
.B1(n_104),
.B2(n_83),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_81),
.A2(n_64),
.B1(n_46),
.B2(n_26),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_135),
.A2(n_91),
.B1(n_79),
.B2(n_110),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_44),
.B1(n_35),
.B2(n_33),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_112),
.B1(n_109),
.B2(n_80),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_46),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_136),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_146),
.C(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_144),
.B(n_151),
.Y(n_198)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_145),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_88),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_120),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_106),
.B1(n_75),
.B2(n_88),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_159),
.B1(n_169),
.B2(n_176),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_95),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_152),
.B(n_158),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_153),
.A2(n_154),
.B(n_175),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_111),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_100),
.B1(n_103),
.B2(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_174),
.B1(n_127),
.B2(n_115),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_35),
.B(n_33),
.C(n_20),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_164),
.B(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_100),
.B1(n_20),
.B2(n_35),
.Y(n_159)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_166),
.B1(n_168),
.B2(n_122),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_165),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_41),
.B(n_2),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_172),
.B(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_118),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_41),
.B(n_35),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_41),
.C(n_84),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_170),
.C(n_162),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_116),
.A2(n_33),
.B1(n_26),
.B2(n_96),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_26),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_133),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_33),
.B1(n_92),
.B2(n_84),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_1),
.B(n_2),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_74),
.B1(n_2),
.B2(n_3),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_177),
.A2(n_185),
.B(n_202),
.Y(n_226)
);

XNOR2x2_ASAP7_75t_SL g180 ( 
.A(n_143),
.B(n_128),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_204),
.B(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_182),
.B(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_118),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_194),
.C(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_113),
.B1(n_121),
.B2(n_127),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_191),
.B1(n_197),
.B2(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_113),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_120),
.B1(n_140),
.B2(n_130),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_196),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_144),
.A2(n_130),
.B1(n_117),
.B2(n_138),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_117),
.B1(n_74),
.B2(n_4),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_15),
.C(n_14),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_12),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_1),
.B(n_3),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_157),
.B(n_5),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_1),
.B(n_3),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g236 ( 
.A(n_206),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_155),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_211),
.C(n_214),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_167),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_200),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_227),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_216),
.B(n_228),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_170),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_154),
.B(n_158),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_234),
.C(n_237),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_165),
.B1(n_157),
.B2(n_145),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_225),
.B1(n_229),
.B2(n_232),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_4),
.B(n_5),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_177),
.A2(n_4),
.B(n_6),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_188),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_233),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_178),
.A2(n_160),
.B(n_7),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_184),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_11),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_4),
.C(n_7),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_178),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_259),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_242),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_182),
.B1(n_206),
.B2(n_179),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_258),
.B1(n_225),
.B2(n_191),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_216),
.B(n_198),
.CI(n_190),
.CON(n_245),
.SN(n_245)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_252),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_253),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_204),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_256),
.C(n_260),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_255),
.A2(n_257),
.B1(n_181),
.B2(n_219),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_222),
.C(n_234),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_217),
.A2(n_179),
.B1(n_185),
.B2(n_202),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_186),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_219),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_262),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_277),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_215),
.C(n_231),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_273),
.C(n_278),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_228),
.B(n_229),
.C(n_232),
.D(n_226),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_245),
.B(n_240),
.C(n_243),
.D(n_203),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_217),
.B1(n_187),
.B2(n_215),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_272),
.A2(n_274),
.B1(n_246),
.B2(n_258),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_212),
.C(n_230),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_223),
.B1(n_230),
.B2(n_190),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_260),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_251),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_197),
.C(n_220),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_220),
.C(n_181),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.C(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_209),
.C(n_207),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_246),
.B1(n_257),
.B2(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_289),
.B(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_290),
.C(n_267),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_245),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_271),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_203),
.C(n_8),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_273),
.C(n_279),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_300)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_296),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_268),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_280),
.C(n_267),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_307),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_308),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_285),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_268),
.C(n_276),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_284),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_307),
.C(n_293),
.Y(n_326)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_281),
.B1(n_287),
.B2(n_292),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_291),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_295),
.Y(n_321)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_298),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_326),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_306),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_325),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_313),
.B(n_315),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_330),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_328),
.A2(n_323),
.B(n_324),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_329),
.Y(n_333)
);

OAI221xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_331),
.B1(n_327),
.B2(n_314),
.C(n_320),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_304),
.B1(n_310),
.B2(n_311),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_10),
.B(n_316),
.C(n_310),
.Y(n_337)
);


endmodule