module fake_ariane_1847_n_137 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_54, n_25, n_137);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_54;
input n_25;

output n_137;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_119;
wire n_124;
wire n_90;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_120;
wire n_106;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_100;
wire n_132;
wire n_62;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_82;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_85;
wire n_130;
wire n_94;
wire n_101;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_112;
wire n_129;
wire n_126;
wire n_122;
wire n_135;
wire n_73;
wire n_77;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_81;
wire n_87;
wire n_136;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_63;
wire n_59;
wire n_99;
wire n_127;

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx8_ASAP7_75t_SL g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_18),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_5),
.B(n_6),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

OA21x2_ASAP7_75t_L g70 ( 
.A1(n_35),
.A2(n_40),
.B(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_36),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_31),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_12),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_32),
.B1(n_8),
.B2(n_9),
.Y(n_80)
);

OAI22x1_ASAP7_75t_R g81 ( 
.A1(n_22),
.A2(n_15),
.B1(n_37),
.B2(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_0),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_1),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_1),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_13),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_59),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_14),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_67),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_80),
.B1(n_82),
.B2(n_61),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_60),
.B(n_57),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_62),
.B(n_73),
.C(n_58),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_83),
.Y(n_105)
);

BUFx6f_ASAP7_75t_SL g106 ( 
.A(n_97),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_83),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_78),
.B(n_76),
.C(n_70),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_69),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_90),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_96),
.B(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_111),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_106),
.Y(n_126)
);

OAI211xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_86),
.B(n_121),
.C(n_118),
.Y(n_127)
);

OAI211xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_116),
.B(n_92),
.C(n_124),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_116),
.B1(n_96),
.B2(n_123),
.C(n_106),
.Y(n_130)
);

NOR4xp25_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_66),
.C(n_17),
.D(n_34),
.Y(n_131)
);

NOR4xp75_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_129),
.C(n_66),
.D(n_43),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_132),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_16),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_66),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_134),
.B1(n_46),
.B2(n_50),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_41),
.Y(n_137)
);


endmodule