module fake_jpeg_946_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

OR2x2_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_1),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_10),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_16),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_19),
.B(n_15),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_34),
.B(n_30),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_15),
.B(n_22),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_20),
.B1(n_18),
.B2(n_9),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_30),
.B1(n_23),
.B2(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_36),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_27),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_21),
.C(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_32),
.B1(n_20),
.B2(n_9),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_26),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_42),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_32),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_6),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_40),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_21),
.C(n_6),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_43),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_41),
.B(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_21),
.C(n_3),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

AOI322xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_2),
.A3(n_4),
.B1(n_48),
.B2(n_50),
.C1(n_52),
.C2(n_51),
.Y(n_54)
);


endmodule