module fake_netlist_1_3580_n_537 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_537);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_537;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_60), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_76), .Y(n_78) );
INVxp67_ASAP7_75t_L g79 ( .A(n_23), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_15), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_34), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_64), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_39), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_40), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_47), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_16), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_6), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_26), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_48), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_35), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_46), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_32), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_72), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_33), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_11), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_9), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_62), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_1), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_8), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_51), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_69), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_52), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_68), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_16), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_63), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_10), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_1), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_29), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_38), .Y(n_114) );
INVx6_ASAP7_75t_L g115 ( .A(n_109), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_95), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_109), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_108), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_94), .B(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_89), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_95), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
INVx6_ASAP7_75t_L g124 ( .A(n_79), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_110), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_112), .Y(n_127) );
BUFx10_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_112), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_87), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_80), .B(n_0), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_100), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_96), .B(n_2), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_117), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_117), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_117), .Y(n_139) );
BUFx10_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_124), .B(n_97), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_122), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_122), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_122), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_117), .Y(n_145) );
INVx4_ASAP7_75t_SL g146 ( .A(n_115), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_122), .Y(n_147) );
INVx2_ASAP7_75t_SL g148 ( .A(n_115), .Y(n_148) );
OR2x2_ASAP7_75t_L g149 ( .A(n_129), .B(n_88), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_127), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_123), .B(n_103), .Y(n_151) );
OR2x2_ASAP7_75t_L g152 ( .A(n_127), .B(n_98), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_128), .B(n_120), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_128), .B(n_98), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_122), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_135), .B(n_84), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_130), .Y(n_157) );
NAND2xp33_ASAP7_75t_L g158 ( .A(n_130), .B(n_84), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_123), .B(n_104), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_124), .B(n_105), .Y(n_161) );
AO22x1_ASAP7_75t_L g162 ( .A1(n_150), .A2(n_100), .B1(n_91), .B2(n_78), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
OR2x2_ASAP7_75t_L g164 ( .A(n_150), .B(n_133), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_153), .A2(n_132), .B1(n_136), .B2(n_119), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_154), .B(n_128), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_157), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_154), .B(n_126), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_154), .B(n_124), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_153), .Y(n_174) );
BUFx12f_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_160), .B(n_131), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_160), .B(n_131), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_134), .B1(n_81), .B2(n_82), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_149), .A2(n_111), .B1(n_102), .B2(n_99), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_141), .B(n_124), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_149), .B(n_111), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_137), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_141), .B(n_161), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_152), .B(n_121), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_152), .B(n_125), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_137), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_161), .B(n_106), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_168), .A2(n_158), .B(n_148), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_181), .A2(n_101), .B(n_116), .C(n_121), .Y(n_195) );
CKINVDCx11_ASAP7_75t_R g196 ( .A(n_175), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_181), .A2(n_171), .B(n_172), .C(n_168), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_172), .A2(n_148), .B(n_155), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_178), .B(n_118), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_178), .A2(n_118), .B1(n_125), .B2(n_116), .Y(n_202) );
AND2x4_ASAP7_75t_SL g203 ( .A(n_170), .B(n_140), .Y(n_203) );
NAND2xp33_ASAP7_75t_SL g204 ( .A(n_174), .B(n_135), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_174), .B(n_146), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_163), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_170), .B(n_144), .Y(n_207) );
AO22x1_ASAP7_75t_L g208 ( .A1(n_167), .A2(n_85), .B1(n_86), .B2(n_90), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_85), .B(n_113), .C(n_86), .Y(n_209) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_163), .A2(n_138), .B(n_139), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_175), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_176), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_166), .A2(n_155), .B(n_138), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_170), .B(n_140), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_186), .A2(n_138), .B(n_145), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_115), .B1(n_135), .B2(n_93), .Y(n_218) );
OR2x6_ASAP7_75t_SL g219 ( .A(n_164), .B(n_90), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_169), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_177), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_177), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_170), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_187), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_214), .Y(n_226) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_210), .A2(n_139), .B(n_145), .Y(n_227) );
AOI21xp5_ASAP7_75t_SL g228 ( .A1(n_221), .A2(n_92), .B(n_93), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_222), .B(n_183), .Y(n_229) );
OAI21x1_ASAP7_75t_SL g230 ( .A1(n_198), .A2(n_173), .B(n_107), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
OAI21x1_ASAP7_75t_L g232 ( .A1(n_210), .A2(n_139), .B(n_145), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_203), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_223), .A2(n_164), .B1(n_188), .B2(n_183), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_203), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_199), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_201), .B(n_165), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_220), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_220), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_197), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_209), .A2(n_191), .B(n_182), .C(n_92), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_200), .A2(n_107), .B(n_113), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_196), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_225), .B(n_162), .Y(n_244) );
O2A1O1Ixp5_ASAP7_75t_SL g245 ( .A1(n_218), .A2(n_114), .B(n_159), .C(n_147), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_217), .A2(n_193), .B(n_192), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_224), .B(n_162), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_196), .Y(n_248) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_194), .A2(n_193), .B(n_192), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_204), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_206), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_197), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_237), .A2(n_202), .B1(n_212), .B2(n_213), .Y(n_253) );
AO222x2_ASAP7_75t_L g254 ( .A1(n_248), .A2(n_219), .B1(n_4), .B2(n_5), .C1(n_6), .C2(n_7), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_226), .A2(n_216), .B1(n_209), .B2(n_207), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_226), .A2(n_216), .B1(n_207), .B2(n_195), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_238), .A2(n_215), .B(n_204), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_234), .A2(n_206), .B1(n_205), .B2(n_211), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_229), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_229), .A2(n_206), .B1(n_197), .B2(n_211), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_233), .A2(n_211), .B1(n_197), .B2(n_208), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_247), .A2(n_205), .B1(n_211), .B2(n_179), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_233), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_231), .B(n_205), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_247), .A2(n_179), .B1(n_180), .B2(n_135), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_236), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_244), .A2(n_180), .B1(n_117), .B2(n_144), .C(n_147), .Y(n_268) );
AOI222xp33_ASAP7_75t_L g269 ( .A1(n_244), .A2(n_146), .B1(n_140), .B2(n_7), .C1(n_8), .C2(n_9), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_238), .A2(n_185), .B(n_189), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_236), .B(n_146), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g272 ( .A1(n_235), .A2(n_140), .B1(n_144), .B2(n_147), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_238), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_235), .A2(n_193), .B1(n_192), .B2(n_169), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_273), .B(n_239), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_273), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_266), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_266), .B(n_239), .Y(n_278) );
INVx5_ASAP7_75t_SL g279 ( .A(n_271), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_259), .B(n_267), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_264), .B(n_240), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_263), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
AOI21x1_ASAP7_75t_L g286 ( .A1(n_257), .A2(n_249), .B(n_230), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_269), .B(n_240), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_255), .Y(n_289) );
INVx4_ASAP7_75t_L g290 ( .A(n_271), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_271), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_256), .B(n_230), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_274), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_261), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_269), .B(n_252), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_262), .B(n_252), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_275), .B(n_240), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_277), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_286), .A2(n_249), .B(n_270), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_275), .B(n_252), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_276), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_275), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_278), .B(n_265), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_278), .B(n_253), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_278), .B(n_228), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_283), .B(n_228), .Y(n_310) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_292), .A2(n_258), .B1(n_254), .B2(n_241), .C(n_268), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_276), .B(n_246), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_281), .B(n_289), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_283), .B(n_245), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_283), .B(n_245), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_282), .B(n_242), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_281), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_250), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_282), .Y(n_320) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_292), .A2(n_250), .B1(n_272), .B2(n_251), .C(n_243), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_287), .B(n_251), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_285), .Y(n_325) );
NOR3xp33_ASAP7_75t_L g326 ( .A(n_311), .B(n_285), .C(n_295), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_298), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_298), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_306), .B(n_288), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_317), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_312), .B(n_288), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_299), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_309), .A2(n_295), .B1(n_287), .B2(n_291), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_311), .B(n_295), .C(n_287), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_317), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_324), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_313), .B(n_294), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_324), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_309), .A2(n_291), .B1(n_290), .B2(n_296), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_303), .B(n_294), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_303), .B(n_294), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_305), .B(n_293), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_306), .B(n_291), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_305), .B(n_293), .Y(n_346) );
OAI211xp5_ASAP7_75t_SL g347 ( .A1(n_321), .A2(n_293), .B(n_147), .C(n_159), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_300), .B(n_296), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_318), .B(n_322), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_318), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_322), .B(n_296), .Y(n_351) );
AOI22x1_ASAP7_75t_L g352 ( .A1(n_304), .A2(n_290), .B1(n_279), .B2(n_10), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_304), .B(n_290), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_313), .B(n_279), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_297), .B(n_290), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_308), .B(n_279), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_320), .Y(n_358) );
OAI211xp5_ASAP7_75t_L g359 ( .A1(n_321), .A2(n_3), .B(n_5), .C(n_11), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
OR2x4_ASAP7_75t_L g361 ( .A(n_319), .B(n_279), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_308), .A2(n_144), .B(n_147), .C(n_159), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_297), .B(n_279), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_325), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_302), .B(n_279), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_302), .B(n_242), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_312), .B(n_12), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_349), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_348), .B(n_312), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_339), .B(n_312), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_326), .A2(n_315), .B(n_314), .Y(n_372) );
NOR2xp33_ASAP7_75t_SL g373 ( .A(n_368), .B(n_316), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_348), .B(n_316), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_349), .B(n_323), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_339), .B(n_319), .Y(n_376) );
AND4x1_ASAP7_75t_L g377 ( .A(n_336), .B(n_310), .C(n_323), .D(n_14), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_331), .B(n_310), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_332), .B(n_301), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_332), .B(n_301), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_337), .B(n_351), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_334), .B(n_307), .C(n_314), .D(n_315), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_332), .B(n_301), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_338), .Y(n_384) );
NOR2xp67_ASAP7_75t_SL g385 ( .A(n_359), .B(n_307), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_332), .B(n_301), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_338), .Y(n_387) );
AND2x2_ASAP7_75t_SL g388 ( .A(n_368), .B(n_12), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_351), .B(n_13), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_354), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_365), .B(n_13), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_329), .B(n_14), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_329), .B(n_15), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_365), .B(n_17), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_345), .B(n_17), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_345), .B(n_18), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_327), .Y(n_399) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_359), .B(n_19), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_341), .B(n_159), .C(n_144), .D(n_19), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_356), .B(n_246), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_327), .B(n_232), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_338), .Y(n_404) );
INVx3_ASAP7_75t_SL g405 ( .A(n_358), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_328), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_356), .B(n_232), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_328), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_362), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_330), .B(n_227), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_330), .B(n_227), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_333), .B(n_20), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_342), .B(n_159), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_333), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_352), .B(n_363), .C(n_347), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_335), .B(n_22), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_335), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_361), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_342), .B(n_24), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_343), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_395), .Y(n_422) );
OAI321xp33_ASAP7_75t_L g423 ( .A1(n_401), .A2(n_347), .A3(n_355), .B1(n_353), .B2(n_358), .C(n_357), .Y(n_423) );
OAI33xp33_ASAP7_75t_L g424 ( .A1(n_381), .A2(n_389), .A3(n_391), .B1(n_394), .B2(n_378), .B3(n_369), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_373), .A2(n_361), .B1(n_355), .B2(n_352), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_377), .A2(n_357), .B1(n_343), .B2(n_363), .C(n_344), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_388), .A2(n_361), .B1(n_366), .B2(n_364), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_420), .B(n_346), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_372), .A2(n_344), .B1(n_346), .B2(n_364), .C(n_366), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_374), .B(n_367), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_376), .B(n_367), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_374), .B(n_360), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_376), .B(n_360), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_418), .B(n_360), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_405), .B(n_340), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_390), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_405), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_399), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_375), .B(n_340), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_385), .A2(n_340), .B1(n_190), .B2(n_189), .C(n_185), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
INVx5_ASAP7_75t_L g444 ( .A(n_418), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_388), .A2(n_190), .B1(n_189), .B2(n_185), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_371), .B(n_27), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_392), .B(n_30), .Y(n_447) );
AOI31xp33_ASAP7_75t_L g448 ( .A1(n_394), .A2(n_31), .A3(n_36), .B(n_37), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_415), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_449) );
OAI321xp33_ASAP7_75t_L g450 ( .A1(n_382), .A2(n_44), .A3(n_45), .B1(n_49), .B2(n_50), .C(n_53), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_379), .B(n_54), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g452 ( .A1(n_385), .A2(n_55), .B(n_56), .Y(n_452) );
NAND2x1_ASAP7_75t_SL g453 ( .A(n_400), .B(n_57), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_384), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_408), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_392), .A2(n_58), .B1(n_59), .B2(n_61), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_393), .B(n_66), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_393), .B(n_67), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_397), .A2(n_189), .B1(n_185), .B2(n_190), .C(n_184), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_371), .B(n_70), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_384), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g462 ( .A(n_397), .B(n_71), .C(n_73), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_409), .A2(n_190), .B1(n_189), .B2(n_185), .C(n_184), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_370), .B(n_74), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_370), .B(n_75), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_430), .B(n_386), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_424), .A2(n_428), .B1(n_425), .B2(n_445), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_423), .A2(n_398), .B(n_419), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_421), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_436), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_433), .B(n_380), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_423), .A2(n_398), .B(n_419), .Y(n_474) );
INVxp33_ASAP7_75t_SL g475 ( .A(n_445), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_432), .B(n_402), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_443), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_444), .B(n_379), .Y(n_478) );
AO22x1_ASAP7_75t_L g479 ( .A1(n_439), .A2(n_379), .B1(n_386), .B2(n_383), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_429), .B(n_383), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_455), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_441), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_427), .A2(n_380), .B1(n_417), .B2(n_414), .C(n_402), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_438), .A2(n_407), .B1(n_412), .B2(n_404), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_454), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_462), .A2(n_407), .B1(n_412), .B2(n_410), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_461), .B(n_387), .Y(n_490) );
XOR2xp5_ASAP7_75t_L g491 ( .A(n_464), .B(n_413), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_435), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_453), .B(n_452), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_435), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_482), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_467), .A2(n_448), .B(n_447), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_479), .A2(n_448), .B(n_450), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_478), .A2(n_444), .B(n_451), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_469), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_484), .A2(n_456), .B1(n_457), .B2(n_458), .C(n_442), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_474), .A2(n_449), .B(n_465), .C(n_460), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_492), .Y(n_503) );
NOR2xp67_ASAP7_75t_L g504 ( .A(n_478), .B(n_444), .Y(n_504) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_475), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_470), .Y(n_506) );
INVxp33_ASAP7_75t_SL g507 ( .A(n_491), .Y(n_507) );
XOR2xp5_ASAP7_75t_L g508 ( .A(n_468), .B(n_446), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_487), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_484), .A2(n_459), .B1(n_451), .B2(n_463), .C(n_416), .Y(n_510) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_494), .B(n_413), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_486), .B(n_404), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_466), .A2(n_387), .B1(n_410), .B2(n_403), .C(n_411), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_511), .B(n_473), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_505), .A2(n_489), .B1(n_485), .B2(n_494), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_497), .A2(n_477), .B(n_481), .C(n_472), .Y(n_516) );
AOI222xp33_ASAP7_75t_L g517 ( .A1(n_513), .A2(n_503), .B1(n_507), .B2(n_496), .C1(n_504), .C2(n_506), .Y(n_517) );
AOI221xp5_ASAP7_75t_SL g518 ( .A1(n_497), .A2(n_489), .B1(n_495), .B2(n_493), .C(n_483), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g519 ( .A(n_498), .B(n_480), .C(n_471), .D(n_493), .Y(n_519) );
O2A1O1Ixp5_ASAP7_75t_L g520 ( .A1(n_499), .A2(n_488), .B(n_490), .C(n_476), .Y(n_520) );
AOI211xp5_ASAP7_75t_SL g521 ( .A1(n_502), .A2(n_184), .B(n_146), .C(n_140), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_SL g522 ( .A1(n_512), .A2(n_146), .B(n_185), .C(n_189), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_516), .Y(n_523) );
NAND3xp33_ASAP7_75t_SL g524 ( .A(n_517), .B(n_508), .C(n_501), .Y(n_524) );
NAND4xp75_ASAP7_75t_L g525 ( .A(n_518), .B(n_510), .C(n_500), .D(n_509), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_519), .A2(n_146), .B1(n_190), .B2(n_520), .C(n_515), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_514), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_525), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_524), .Y(n_529) );
NOR3xp33_ASAP7_75t_SL g530 ( .A(n_523), .B(n_521), .C(n_522), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_528), .B(n_527), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_529), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_531), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_533), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_534), .A2(n_528), .B1(n_532), .B2(n_526), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_535), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_536), .A2(n_530), .B1(n_522), .B2(n_190), .Y(n_537) );
endmodule