module fake_netlist_1_10649_n_25 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_25);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx16_ASAP7_75t_R g9 ( .A(n_4), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_8), .B(n_7), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_9), .B(n_0), .Y(n_15) );
OAI21x1_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_0), .B(n_1), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_10), .A2(n_2), .B(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_15), .B(n_13), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_17), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_14), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_20), .B(n_16), .Y(n_22) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_22), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_12), .B1(n_17), .B2(n_5), .Y(n_24) );
AOI22xp33_ASAP7_75t_R g25 ( .A1(n_24), .A2(n_12), .B1(n_2), .B2(n_3), .Y(n_25) );
endmodule