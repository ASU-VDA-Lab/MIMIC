module real_aes_8952_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g263 ( .A1(n_0), .A2(n_264), .B(n_265), .C(n_268), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_1), .B(n_252), .Y(n_269) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_3), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_4), .A2(n_141), .B(n_144), .C(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_5), .A2(n_136), .B(n_568), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_6), .A2(n_136), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_7), .B(n_252), .Y(n_574) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_8), .A2(n_171), .B(n_208), .Y(n_207) );
AND2x6_ASAP7_75t_L g141 ( .A(n_9), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_10), .A2(n_141), .B(n_144), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g512 ( .A(n_11), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_12), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_12), .B(n_40), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_13), .B(n_228), .Y(n_546) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_15), .B(n_180), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_16), .A2(n_181), .B(n_530), .C(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_17), .B(n_252), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_18), .B(n_156), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_19), .A2(n_144), .B(n_147), .C(n_155), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_20), .A2(n_216), .B(n_267), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_21), .B(n_228), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_22), .A2(n_123), .B1(n_124), .B2(n_452), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_22), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_23), .B(n_228), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g559 ( .A(n_24), .Y(n_559) );
INVx1_ASAP7_75t_L g484 ( .A(n_25), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_26), .A2(n_144), .B(n_155), .C(n_211), .Y(n_210) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_28), .Y(n_542) );
INVx1_ASAP7_75t_L g500 ( .A(n_29), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_30), .B(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_31), .A2(n_136), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g139 ( .A(n_32), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_33), .A2(n_184), .B(n_193), .C(n_195), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_34), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_35), .A2(n_267), .B(n_571), .C(n_573), .Y(n_570) );
INVxp67_ASAP7_75t_L g501 ( .A(n_36), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_37), .B(n_213), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_38), .A2(n_144), .B(n_155), .C(n_483), .Y(n_482) );
CKINVDCx14_ASAP7_75t_R g569 ( .A(n_39), .Y(n_569) );
INVx1_ASAP7_75t_L g114 ( .A(n_40), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_41), .A2(n_268), .B(n_510), .C(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_42), .B(n_135), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_43), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_44), .B(n_180), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_45), .B(n_136), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_46), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_47), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_48), .A2(n_184), .B(n_193), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g266 ( .A(n_49), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_50), .A2(n_125), .B1(n_126), .B2(n_451), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_50), .Y(n_125) );
INVx1_ASAP7_75t_L g238 ( .A(n_51), .Y(n_238) );
INVx1_ASAP7_75t_L g518 ( .A(n_52), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_53), .B(n_136), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_54), .Y(n_164) );
CKINVDCx14_ASAP7_75t_R g508 ( .A(n_55), .Y(n_508) );
INVx1_ASAP7_75t_L g142 ( .A(n_56), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_57), .B(n_136), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_58), .B(n_252), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_59), .A2(n_154), .B(n_177), .C(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g161 ( .A(n_60), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_61), .A2(n_100), .B1(n_465), .B2(n_466), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_61), .Y(n_466) );
INVx1_ASAP7_75t_SL g572 ( .A(n_62), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_63), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_64), .B(n_180), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_65), .B(n_252), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_66), .B(n_181), .Y(n_226) );
INVx1_ASAP7_75t_L g562 ( .A(n_67), .Y(n_562) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_68), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_69), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_70), .A2(n_144), .B(n_175), .C(n_184), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_71), .Y(n_247) );
INVx1_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_73), .A2(n_136), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_74), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_75), .A2(n_136), .B(n_527), .Y(n_526) );
AOI222xp33_ASAP7_75t_SL g463 ( .A1(n_76), .A2(n_464), .B1(n_467), .B2(n_747), .C1(n_748), .C2(n_752), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_77), .A2(n_135), .B(n_496), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_78), .Y(n_481) );
INVx1_ASAP7_75t_L g528 ( .A(n_79), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_80), .B(n_152), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_81), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_82), .A2(n_136), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g531 ( .A(n_83), .Y(n_531) );
INVx2_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
INVx1_ASAP7_75t_L g545 ( .A(n_85), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_86), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_87), .B(n_228), .Y(n_227) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_88), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g456 ( .A(n_88), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g470 ( .A(n_88), .B(n_458), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_88), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_89), .A2(n_144), .B(n_184), .C(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_90), .B(n_136), .Y(n_191) );
INVx1_ASAP7_75t_L g196 ( .A(n_91), .Y(n_196) );
INVxp67_ASAP7_75t_L g250 ( .A(n_92), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_93), .A2(n_102), .B1(n_115), .B2(n_756), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_94), .B(n_171), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_95), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g176 ( .A(n_96), .Y(n_176) );
INVx1_ASAP7_75t_L g222 ( .A(n_97), .Y(n_222) );
INVx2_ASAP7_75t_L g521 ( .A(n_98), .Y(n_521) );
AND2x2_ASAP7_75t_L g240 ( .A(n_99), .B(n_158), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_100), .Y(n_465) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx4f_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g756 ( .A(n_105), .Y(n_756) );
AND2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_112), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g458 ( .A(n_108), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_462), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g755 ( .A(n_120), .Y(n_755) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_453), .B(n_460), .Y(n_121) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_126), .A2(n_474), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx2_ASAP7_75t_L g451 ( .A(n_127), .Y(n_451) );
AND3x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_355), .C(n_412), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_300), .C(n_336), .Y(n_128) );
OAI211xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_202), .B(n_254), .C(n_287), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g257 ( .A(n_132), .B(n_258), .Y(n_257) );
INVx5_ASAP7_75t_L g286 ( .A(n_132), .Y(n_286) );
AND2x2_ASAP7_75t_L g359 ( .A(n_132), .B(n_275), .Y(n_359) );
AND2x2_ASAP7_75t_L g397 ( .A(n_132), .B(n_303), .Y(n_397) );
AND2x2_ASAP7_75t_L g417 ( .A(n_132), .B(n_259), .Y(n_417) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_163), .Y(n_132) );
AOI21xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_143), .B(n_156), .Y(n_133) );
BUFx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_137), .B(n_141), .Y(n_223) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
INVx1_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
INVx3_ASAP7_75t_L g181 ( .A(n_140), .Y(n_181) );
INVx1_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_140), .Y(n_228) );
BUFx3_ASAP7_75t_L g155 ( .A(n_141), .Y(n_155) );
INVx4_ASAP7_75t_SL g185 ( .A(n_141), .Y(n_185) );
INVx5_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
BUFx3_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_153), .Y(n_147) );
INVx2_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_152), .A2(n_196), .B(n_197), .C(n_198), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_152), .A2(n_198), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp5_ASAP7_75t_L g544 ( .A1(n_152), .A2(n_545), .B(n_546), .C(n_547), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_152), .A2(n_547), .B(n_562), .C(n_563), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_153), .A2(n_180), .B(n_484), .C(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_154), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_157), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_158), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_158), .A2(n_235), .B(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_158), .A2(n_223), .B(n_481), .C(n_482), .Y(n_480) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_158), .A2(n_506), .B(n_513), .Y(n_505) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g172 ( .A(n_159), .B(n_160), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_165), .A2(n_541), .B(n_548), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_166), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_189), .Y(n_166) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_167), .Y(n_298) );
AND2x2_ASAP7_75t_L g312 ( .A(n_167), .B(n_258), .Y(n_312) );
INVx1_ASAP7_75t_L g335 ( .A(n_167), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_167), .B(n_286), .Y(n_374) );
OR2x2_ASAP7_75t_L g411 ( .A(n_167), .B(n_256), .Y(n_411) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_168), .Y(n_347) );
AND2x2_ASAP7_75t_L g354 ( .A(n_168), .B(n_259), .Y(n_354) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g275 ( .A(n_169), .B(n_259), .Y(n_275) );
BUFx2_ASAP7_75t_L g303 ( .A(n_169), .Y(n_303) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_187), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_170), .B(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_170), .B(n_201), .Y(n_200) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_170), .A2(n_221), .B(n_229), .Y(n_220) );
INVx3_ASAP7_75t_L g252 ( .A(n_170), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_170), .B(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_170), .B(n_549), .Y(n_548) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_170), .A2(n_558), .B(n_564), .Y(n_557) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_171), .A2(n_209), .B(n_210), .Y(n_208) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_186), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_179), .C(n_182), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_178), .A2(n_180), .B1(n_500), .B2(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_178), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_178), .B(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_180), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g264 ( .A(n_180), .Y(n_264) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_181), .B(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g573 ( .A(n_183), .Y(n_573) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_185), .A2(n_194), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g261 ( .A1(n_185), .A2(n_194), .B(n_262), .C(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_185), .A2(n_194), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_185), .A2(n_194), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_185), .A2(n_194), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_185), .A2(n_194), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g568 ( .A1(n_185), .A2(n_194), .B(n_569), .C(n_570), .Y(n_568) );
INVx5_ASAP7_75t_L g256 ( .A(n_189), .Y(n_256) );
BUFx2_ASAP7_75t_L g279 ( .A(n_189), .Y(n_279) );
AND2x2_ASAP7_75t_L g436 ( .A(n_189), .B(n_290), .Y(n_436) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_200), .Y(n_189) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g268 ( .A(n_199), .Y(n_268) );
INVx1_ASAP7_75t_L g532 ( .A(n_199), .Y(n_532) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_241), .Y(n_203) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_204), .A2(n_337), .B1(n_344), .B2(n_345), .C(n_348), .Y(n_336) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_218), .Y(n_204) );
AND2x2_ASAP7_75t_L g242 ( .A(n_205), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_205), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g271 ( .A(n_206), .B(n_219), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_206), .B(n_220), .Y(n_281) );
OR2x2_ASAP7_75t_L g292 ( .A(n_206), .B(n_243), .Y(n_292) );
AND2x2_ASAP7_75t_L g295 ( .A(n_206), .B(n_283), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_206), .B(n_232), .Y(n_311) );
OR2x2_ASAP7_75t_L g327 ( .A(n_206), .B(n_220), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_206), .B(n_243), .Y(n_389) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_207), .B(n_232), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_207), .B(n_220), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_214), .B(n_215), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_215), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g305 ( .A(n_218), .B(n_292), .Y(n_305) );
INVx2_ASAP7_75t_L g331 ( .A(n_218), .Y(n_331) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_232), .Y(n_218) );
AND2x2_ASAP7_75t_L g253 ( .A(n_219), .B(n_233), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_219), .B(n_243), .Y(n_310) );
OR2x2_ASAP7_75t_L g321 ( .A(n_219), .B(n_233), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_219), .B(n_283), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_219), .A2(n_414), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_413) );
INVx5_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_220), .B(n_243), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_223), .A2(n_542), .B(n_543), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_223), .A2(n_559), .B(n_560), .Y(n_558) );
INVx4_ASAP7_75t_L g267 ( .A(n_228), .Y(n_267) );
INVx2_ASAP7_75t_L g510 ( .A(n_228), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g493 ( .A(n_231), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_232), .B(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_232), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g299 ( .A(n_232), .B(n_271), .Y(n_299) );
OR2x2_ASAP7_75t_L g343 ( .A(n_232), .B(n_243), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_232), .B(n_295), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_232), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g408 ( .A(n_232), .B(n_409), .Y(n_408) );
INVx5_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_233), .B(n_242), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_SL g276 ( .A1(n_233), .A2(n_277), .B(n_280), .C(n_284), .Y(n_276) );
OR2x2_ASAP7_75t_L g314 ( .A(n_233), .B(n_310), .Y(n_314) );
OR2x2_ASAP7_75t_L g350 ( .A(n_233), .B(n_292), .Y(n_350) );
OAI311xp33_ASAP7_75t_L g356 ( .A1(n_233), .A2(n_295), .A3(n_357), .B1(n_360), .C1(n_367), .Y(n_356) );
AND2x2_ASAP7_75t_L g407 ( .A(n_233), .B(n_243), .Y(n_407) );
AND2x2_ASAP7_75t_L g415 ( .A(n_233), .B(n_270), .Y(n_415) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_233), .Y(n_433) );
AND2x2_ASAP7_75t_L g450 ( .A(n_233), .B(n_271), .Y(n_450) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_253), .Y(n_241) );
AND2x2_ASAP7_75t_L g278 ( .A(n_242), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g434 ( .A(n_242), .Y(n_434) );
AND2x2_ASAP7_75t_L g270 ( .A(n_243), .B(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g283 ( .A(n_243), .Y(n_283) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
INVxp67_ASAP7_75t_L g365 ( .A(n_243), .Y(n_365) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_251), .Y(n_243) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_244), .A2(n_516), .B(n_522), .Y(n_515) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_244), .A2(n_526), .B(n_533), .Y(n_525) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_244), .A2(n_567), .B(n_574), .Y(n_566) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_252), .A2(n_260), .B(n_269), .Y(n_259) );
AND2x2_ASAP7_75t_L g443 ( .A(n_253), .B(n_291), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_270), .B1(n_272), .B2(n_273), .C(n_276), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_256), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g296 ( .A(n_256), .B(n_286), .Y(n_296) );
AND2x2_ASAP7_75t_L g304 ( .A(n_256), .B(n_258), .Y(n_304) );
OR2x2_ASAP7_75t_L g316 ( .A(n_256), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g334 ( .A(n_256), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g358 ( .A(n_256), .B(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_256), .Y(n_378) );
AND2x2_ASAP7_75t_L g430 ( .A(n_256), .B(n_354), .Y(n_430) );
OAI31xp33_ASAP7_75t_L g438 ( .A1(n_256), .A2(n_307), .A3(n_406), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_257), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g402 ( .A(n_257), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_257), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g290 ( .A(n_258), .B(n_286), .Y(n_290) );
INVx1_ASAP7_75t_L g377 ( .A(n_258), .Y(n_377) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g427 ( .A(n_259), .B(n_286), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_267), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g547 ( .A(n_268), .Y(n_547) );
INVx1_ASAP7_75t_SL g437 ( .A(n_270), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_271), .B(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_272), .A2(n_384), .B1(n_422), .B2(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g285 ( .A(n_275), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g344 ( .A(n_275), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_275), .B(n_296), .Y(n_449) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g419 ( .A(n_278), .B(n_420), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_279), .A2(n_338), .B(n_340), .Y(n_337) );
OR2x2_ASAP7_75t_L g345 ( .A(n_279), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g366 ( .A(n_279), .B(n_354), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_279), .B(n_377), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_279), .B(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_280), .A2(n_394), .B1(n_399), .B2(n_402), .C(n_403), .Y(n_393) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
OR2x2_ASAP7_75t_L g370 ( .A(n_281), .B(n_343), .Y(n_370) );
INVx1_ASAP7_75t_L g409 ( .A(n_281), .Y(n_409) );
INVx2_ASAP7_75t_L g385 ( .A(n_282), .Y(n_385) );
INVx1_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_286), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_286), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g441 ( .A(n_286), .B(n_411), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_291), .B1(n_293), .B2(n_296), .C1(n_297), .C2(n_299), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g297 ( .A(n_290), .B(n_298), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_290), .A2(n_340), .B1(n_368), .B2(n_369), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_290), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OAI21xp33_ASAP7_75t_SL g328 ( .A1(n_299), .A2(n_329), .B(n_332), .Y(n_328) );
OAI211xp5_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_305), .B(n_306), .C(n_328), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_304), .A2(n_307), .B1(n_312), .B2(n_313), .C(n_315), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_304), .B(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g398 ( .A(n_304), .Y(n_398) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
AND2x2_ASAP7_75t_L g400 ( .A(n_309), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g317 ( .A(n_312), .Y(n_317) );
AND2x2_ASAP7_75t_L g323 ( .A(n_312), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_318), .B1(n_322), .B2(n_325), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_319), .B(n_331), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_320), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g420 ( .A(n_324), .Y(n_420) );
AND2x2_ASAP7_75t_L g439 ( .A(n_324), .B(n_354), .Y(n_439) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_331), .B(n_388), .Y(n_447) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_334), .B(n_402), .Y(n_445) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
BUFx2_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_351), .B(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR3xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_371), .C(n_393), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B(n_366), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_375), .B(n_379), .C(n_382), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_372), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2xp67_ASAP7_75t_SL g376 ( .A(n_377), .B(n_378), .Y(n_376) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_SL g401 ( .A(n_381), .Y(n_401) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B(n_390), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AND2x2_ASAP7_75t_L g406 ( .A(n_384), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_408), .B2(n_410), .Y(n_403) );
INVx2_ASAP7_75t_SL g424 ( .A(n_411), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_428), .C(n_440), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_424), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_435), .B2(n_437), .C(n_438), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_429), .A2(n_441), .B(n_442), .C(n_444), .Y(n_440) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_448), .B2(n_450), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_451), .A2(n_468), .B1(n_471), .B2(n_473), .Y(n_467) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g461 ( .A(n_456), .Y(n_461) );
NOR2x2_ASAP7_75t_L g754 ( .A(n_457), .B(n_472), .Y(n_754) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g471 ( .A(n_458), .B(n_472), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_460), .B(n_463), .C(n_755), .Y(n_462) );
INVx1_ASAP7_75t_L g747 ( .A(n_464), .Y(n_747) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g749 ( .A(n_469), .Y(n_749) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g751 ( .A(n_471), .Y(n_751) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
OR5x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_641), .C(n_705), .D(n_721), .E(n_736), .Y(n_474) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_476), .B(n_575), .C(n_602), .D(n_625), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_523), .B(n_534), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx3_ASAP7_75t_SL g554 ( .A(n_479), .Y(n_554) );
AND2x4_ASAP7_75t_L g588 ( .A(n_479), .B(n_577), .Y(n_588) );
OR2x2_ASAP7_75t_L g598 ( .A(n_479), .B(n_556), .Y(n_598) );
OR2x2_ASAP7_75t_L g644 ( .A(n_479), .B(n_491), .Y(n_644) );
AND2x2_ASAP7_75t_L g658 ( .A(n_479), .B(n_555), .Y(n_658) );
AND2x2_ASAP7_75t_L g701 ( .A(n_479), .B(n_591), .Y(n_701) );
AND2x2_ASAP7_75t_L g708 ( .A(n_479), .B(n_566), .Y(n_708) );
AND2x2_ASAP7_75t_L g727 ( .A(n_479), .B(n_617), .Y(n_727) );
AND2x2_ASAP7_75t_L g745 ( .A(n_479), .B(n_587), .Y(n_745) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
INVx1_ASAP7_75t_L g710 ( .A(n_488), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_504), .Y(n_488) );
AND2x2_ASAP7_75t_L g620 ( .A(n_489), .B(n_555), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_489), .B(n_640), .Y(n_639) );
AOI32xp33_ASAP7_75t_L g653 ( .A1(n_489), .A2(n_654), .A3(n_657), .B1(n_659), .B2(n_663), .Y(n_653) );
AND2x2_ASAP7_75t_L g723 ( .A(n_489), .B(n_617), .Y(n_723) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g587 ( .A(n_491), .B(n_556), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_491), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g629 ( .A(n_491), .B(n_576), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_491), .B(n_708), .Y(n_707) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_494), .B(n_502), .Y(n_491) );
INVx1_ASAP7_75t_L g592 ( .A(n_492), .Y(n_592) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OA21x2_ASAP7_75t_L g591 ( .A1(n_495), .A2(n_503), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g594 ( .A(n_504), .B(n_538), .Y(n_594) );
AND2x2_ASAP7_75t_L g670 ( .A(n_504), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g742 ( .A(n_504), .Y(n_742) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
OR2x2_ASAP7_75t_L g537 ( .A(n_505), .B(n_515), .Y(n_537) );
AND2x2_ASAP7_75t_L g551 ( .A(n_505), .B(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_505), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g601 ( .A(n_505), .Y(n_601) );
AND2x2_ASAP7_75t_L g628 ( .A(n_505), .B(n_515), .Y(n_628) );
BUFx3_ASAP7_75t_L g631 ( .A(n_505), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_505), .B(n_606), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_505), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
AND2x2_ASAP7_75t_L g600 ( .A(n_514), .B(n_580), .Y(n_600) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g611 ( .A(n_515), .B(n_525), .Y(n_611) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_515), .Y(n_624) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_524), .B(n_631), .Y(n_681) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_SL g552 ( .A(n_525), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_525), .B(n_600), .C(n_601), .Y(n_599) );
OR2x2_ASAP7_75t_L g607 ( .A(n_525), .B(n_580), .Y(n_607) );
AND2x2_ASAP7_75t_L g627 ( .A(n_525), .B(n_580), .Y(n_627) );
AND2x2_ASAP7_75t_L g671 ( .A(n_525), .B(n_540), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_550), .B(n_553), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g746 ( .A(n_536), .B(n_671), .Y(n_746) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_537), .A2(n_644), .B1(n_686), .B2(n_688), .Y(n_685) );
OR2x2_ASAP7_75t_L g692 ( .A(n_537), .B(n_607), .Y(n_692) );
OR2x2_ASAP7_75t_L g716 ( .A(n_537), .B(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_537), .B(n_636), .Y(n_729) );
AND2x2_ASAP7_75t_L g622 ( .A(n_538), .B(n_623), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_538), .A2(n_695), .B(n_710), .Y(n_709) );
AOI32xp33_ASAP7_75t_L g730 ( .A1(n_538), .A2(n_620), .A3(n_731), .B1(n_733), .B2(n_734), .Y(n_730) );
OR2x2_ASAP7_75t_L g741 ( .A(n_538), .B(n_742), .Y(n_741) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_539), .B(n_623), .Y(n_688) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g580 ( .A(n_540), .Y(n_580) );
AND2x2_ASAP7_75t_L g646 ( .A(n_540), .B(n_611), .Y(n_646) );
AND3x2_ASAP7_75t_L g655 ( .A(n_540), .B(n_551), .C(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g581 ( .A(n_552), .B(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_552), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_552), .B(n_580), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g576 ( .A(n_554), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g616 ( .A(n_554), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g634 ( .A(n_554), .B(n_566), .Y(n_634) );
AND2x2_ASAP7_75t_L g652 ( .A(n_554), .B(n_556), .Y(n_652) );
OR2x2_ASAP7_75t_L g666 ( .A(n_554), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g712 ( .A(n_554), .B(n_640), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_555), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_566), .Y(n_555) );
AND2x2_ASAP7_75t_L g613 ( .A(n_556), .B(n_591), .Y(n_613) );
OR2x2_ASAP7_75t_L g667 ( .A(n_556), .B(n_591), .Y(n_667) );
AND2x2_ASAP7_75t_L g720 ( .A(n_556), .B(n_577), .Y(n_720) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g618 ( .A(n_557), .Y(n_618) );
AND2x2_ASAP7_75t_L g640 ( .A(n_557), .B(n_566), .Y(n_640) );
INVx2_ASAP7_75t_L g577 ( .A(n_566), .Y(n_577) );
INVx1_ASAP7_75t_L g597 ( .A(n_566), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B(n_583), .C(n_595), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_576), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g739 ( .A(n_576), .Y(n_739) );
AND2x2_ASAP7_75t_L g617 ( .A(n_577), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_580), .B(n_581), .Y(n_589) );
INVx1_ASAP7_75t_L g674 ( .A(n_580), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_580), .B(n_601), .Y(n_698) );
AND2x2_ASAP7_75t_L g714 ( .A(n_580), .B(n_628), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_581), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g605 ( .A(n_582), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_589), .B1(n_590), .B2(n_593), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_586), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_587), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g612 ( .A(n_588), .B(n_613), .Y(n_612) );
AOI221xp5_ASAP7_75t_SL g677 ( .A1(n_588), .A2(n_630), .B1(n_678), .B2(n_683), .C(n_685), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_588), .B(n_651), .Y(n_684) );
INVx1_ASAP7_75t_L g744 ( .A(n_590), .Y(n_744) );
BUFx3_ASAP7_75t_L g651 ( .A(n_591), .Y(n_651) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI21xp33_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_598), .B(n_599), .Y(n_595) );
INVx1_ASAP7_75t_L g660 ( .A(n_597), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_597), .B(n_651), .Y(n_704) );
INVx1_ASAP7_75t_L g661 ( .A(n_598), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_598), .B(n_651), .Y(n_662) );
INVxp67_ASAP7_75t_L g682 ( .A(n_600), .Y(n_682) );
AND2x2_ASAP7_75t_L g623 ( .A(n_601), .B(n_624), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_608), .B(n_612), .C(n_614), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_SL g637 ( .A(n_605), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_606), .B(n_637), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_606), .B(n_628), .Y(n_679) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_609), .A2(n_615), .B1(n_619), .B2(n_621), .Y(n_614) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g630 ( .A(n_611), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g675 ( .A(n_611), .B(n_676), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_613), .A2(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_617), .A2(n_626), .B1(n_629), .B2(n_630), .C(n_632), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_617), .B(n_651), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_617), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g733 ( .A(n_623), .Y(n_733) );
INVxp67_ASAP7_75t_L g656 ( .A(n_624), .Y(n_656) );
INVx1_ASAP7_75t_L g663 ( .A(n_626), .Y(n_663) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g702 ( .A(n_627), .B(n_631), .Y(n_702) );
INVx1_ASAP7_75t_L g676 ( .A(n_631), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_631), .B(n_646), .Y(n_706) );
OAI32xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .A3(n_637), .B1(n_638), .B2(n_639), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_SL g645 ( .A(n_640), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_640), .B(n_672), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_640), .B(n_701), .Y(n_732) );
NAND2x1p5_ASAP7_75t_L g740 ( .A(n_640), .B(n_651), .Y(n_740) );
NAND5xp2_ASAP7_75t_L g641 ( .A(n_642), .B(n_664), .C(n_677), .D(n_689), .E(n_690), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_647), .B2(n_649), .C(n_653), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp33_ASAP7_75t_SL g668 ( .A(n_648), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_651), .B(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_652), .A2(n_665), .B1(n_668), .B2(n_672), .Y(n_664) );
INVx2_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_655), .A2(n_660), .B(n_661), .C(n_662), .Y(n_659) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g687 ( .A(n_667), .Y(n_687) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_676), .B(n_725), .Y(n_735) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B1(n_695), .B2(n_699), .C1(n_702), .C2(n_703), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_709), .B2(n_711), .C(n_713), .Y(n_705) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_718), .Y(n_713) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g725 ( .A(n_717), .Y(n_725) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_726), .B2(n_728), .C(n_730), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_740), .B(n_741), .C(n_743), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI21xp33_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_746), .Y(n_743) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx3_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
endmodule