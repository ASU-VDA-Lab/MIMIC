module fake_ibex_464_n_910 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_910);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_910;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx2_ASAP7_75t_SL g171 ( 
.A(n_108),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_49),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_39),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_87),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_65),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_73),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_58),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_95),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_22),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_69),
.Y(n_190)
);

INVx4_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_96),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_27),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_38),
.B(n_25),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_107),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_2),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_25),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_146),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_128),
.Y(n_206)
);

BUFx2_ASAP7_75t_SL g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

INVxp33_ASAP7_75t_SL g209 ( 
.A(n_152),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_76),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_59),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_11),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_82),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_13),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_93),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_13),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_149),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_147),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_117),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_11),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_23),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_68),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_134),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_138),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_30),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_45),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_135),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_55),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_57),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_0),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_126),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_41),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_158),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_144),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_100),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_42),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_124),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_62),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_71),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_83),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_166),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_36),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_78),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_97),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_127),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_81),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_30),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_86),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_141),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_118),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_66),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_75),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_51),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_9),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_12),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_114),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_80),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_6),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_36),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_129),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_29),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_79),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_99),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_32),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_10),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_47),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_26),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_12),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_185),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_201),
.Y(n_282)
);

CKINVDCx11_ASAP7_75t_R g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_1),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_3),
.Y(n_286)
);

CKINVDCx11_ASAP7_75t_R g287 ( 
.A(n_257),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_184),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_184),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_5),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_5),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_246),
.B(n_6),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_205),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_169),
.A2(n_234),
.B(n_227),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_7),
.Y(n_302)
);

AOI22x1_ASAP7_75t_SL g303 ( 
.A1(n_265),
.A2(n_182),
.B1(n_197),
.B2(n_177),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_172),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_186),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_172),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_193),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_169),
.A2(n_91),
.B(n_165),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_195),
.B(n_8),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_172),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_265),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_217),
.Y(n_313)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_205),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_199),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_203),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_172),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_172),
.B(n_15),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_172),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_228),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_223),
.B(n_16),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_228),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_168),
.B(n_17),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_258),
.Y(n_326)
);

CKINVDCx11_ASAP7_75t_R g327 ( 
.A(n_177),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_232),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_237),
.Y(n_330)
);

BUFx8_ASAP7_75t_L g331 ( 
.A(n_234),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_243),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_179),
.B(n_18),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_174),
.B(n_19),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_229),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_176),
.B(n_19),
.Y(n_336)
);

AND2x6_ASAP7_75t_L g337 ( 
.A(n_241),
.B(n_40),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_243),
.Y(n_338)
);

BUFx8_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_233),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g341 ( 
.A(n_170),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g342 ( 
.A(n_279),
.B(n_43),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_238),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_267),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_178),
.B(n_20),
.Y(n_346)
);

CKINVDCx6p67_ASAP7_75t_R g347 ( 
.A(n_253),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_253),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_292),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_285),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_202),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_304),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

AO21x2_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_183),
.B(n_181),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_280),
.B(n_220),
.Y(n_361)
);

BUFx6f_ASAP7_75t_SL g362 ( 
.A(n_282),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_284),
.B(n_226),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_292),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_313),
.A2(n_209),
.B1(n_182),
.B2(n_197),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_288),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_348),
.B(n_187),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_264),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_298),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_L g378 ( 
.A1(n_305),
.A2(n_214),
.B1(n_261),
.B2(n_204),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_288),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_173),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_286),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_209),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_348),
.B(n_190),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_294),
.A2(n_204),
.B1(n_261),
.B2(n_214),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_331),
.B(n_192),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_331),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_SL g392 ( 
.A(n_294),
.B(n_230),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_339),
.B(n_194),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_R g396 ( 
.A(n_305),
.B(n_230),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_L g397 ( 
.A(n_307),
.B(n_200),
.C(n_189),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_329),
.B(n_180),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_329),
.B(n_188),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_337),
.A2(n_255),
.B1(n_271),
.B2(n_275),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_335),
.B(n_212),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_339),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_293),
.B(n_198),
.Y(n_410)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_316),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_324),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_SL g419 ( 
.A1(n_323),
.A2(n_251),
.B(n_196),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_324),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_324),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

NAND2xp33_ASAP7_75t_R g423 ( 
.A(n_326),
.B(n_206),
.Y(n_423)
);

BUFx6f_ASAP7_75t_SL g424 ( 
.A(n_337),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_342),
.B(n_208),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_328),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_323),
.B(n_296),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_337),
.A2(n_278),
.B1(n_171),
.B2(n_207),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_328),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_295),
.Y(n_435)
);

AND2x2_ASAP7_75t_SL g436 ( 
.A(n_308),
.B(n_278),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_330),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_309),
.B(n_325),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_334),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_438),
.B(n_336),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_346),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_351),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_388),
.B(n_303),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_396),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_385),
.A2(n_291),
.B1(n_308),
.B2(n_248),
.Y(n_445)
);

NOR2x2_ASAP7_75t_L g446 ( 
.A(n_378),
.B(n_327),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_371),
.A2(n_312),
.B1(n_281),
.B2(n_287),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_374),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_402),
.B(n_308),
.C(n_219),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_360),
.Y(n_450)
);

OAI221xp5_ASAP7_75t_L g451 ( 
.A1(n_419),
.A2(n_270),
.B1(n_211),
.B2(n_210),
.C(n_213),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_386),
.B(n_215),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_373),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_428),
.B(n_216),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_349),
.B(n_344),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_428),
.B(n_218),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_391),
.B(n_224),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_354),
.A2(n_254),
.B1(n_221),
.B2(n_222),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_406),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_408),
.B(n_225),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_408),
.B(n_239),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_414),
.B(n_242),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_235),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_370),
.B(n_327),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_410),
.B(n_240),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_415),
.B(n_244),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_352),
.B(n_249),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_411),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_392),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_373),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_355),
.A2(n_272),
.B1(n_245),
.B2(n_252),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_396),
.Y(n_476)
);

OAI22xp33_ASAP7_75t_L g477 ( 
.A1(n_357),
.A2(n_312),
.B1(n_262),
.B2(n_260),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_389),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_428),
.B(n_263),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_361),
.B(n_266),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_365),
.B(n_273),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_428),
.B(n_277),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_428),
.B(n_175),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_236),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_376),
.B(n_250),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_432),
.A2(n_297),
.B1(n_295),
.B2(n_320),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_SL g489 ( 
.A(n_424),
.B(n_191),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_368),
.B(n_377),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_356),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

INVx8_ASAP7_75t_L g493 ( 
.A(n_424),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_356),
.B(n_295),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_399),
.B(n_295),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_401),
.B(n_314),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_433),
.A2(n_381),
.B1(n_374),
.B2(n_380),
.Y(n_497)
);

BUFx5_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_379),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_416),
.Y(n_500)
);

AOI21x1_ASAP7_75t_L g501 ( 
.A1(n_380),
.A2(n_320),
.B(n_297),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_381),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_425),
.B(n_330),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_412),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_353),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_460),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_442),
.B(n_397),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_448),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_448),
.A2(n_358),
.B(n_353),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_472),
.A2(n_362),
.B1(n_387),
.B2(n_375),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_497),
.A2(n_359),
.B(n_358),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_439),
.B(n_387),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_491),
.A2(n_366),
.B(n_364),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_440),
.B(n_441),
.Y(n_517)
);

AO22x1_ASAP7_75t_L g518 ( 
.A1(n_476),
.A2(n_283),
.B1(n_287),
.B2(n_423),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_449),
.A2(n_367),
.B(n_369),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_494),
.A2(n_367),
.B(n_369),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_372),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_445),
.A2(n_372),
.B(n_407),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_466),
.B(n_467),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_471),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_447),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_501),
.A2(n_437),
.B(n_382),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_445),
.A2(n_496),
.B(n_495),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_435),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_465),
.B(n_435),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_505),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_477),
.B(n_22),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_24),
.Y(n_532)
);

O2A1O1Ixp33_ASAP7_75t_SL g533 ( 
.A1(n_485),
.A2(n_456),
.B(n_454),
.C(n_479),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_459),
.A2(n_434),
.B1(n_429),
.B2(n_427),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_505),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_468),
.A2(n_407),
.B1(n_427),
.B2(n_421),
.Y(n_536)
);

NOR2x1p5_ASAP7_75t_SL g537 ( 
.A(n_498),
.B(n_384),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_486),
.B(n_350),
.Y(n_538)
);

O2A1O1Ixp33_ASAP7_75t_SL g539 ( 
.A1(n_454),
.A2(n_384),
.B(n_420),
.C(n_418),
.Y(n_539)
);

INVx8_ASAP7_75t_L g540 ( 
.A(n_493),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_489),
.B(n_28),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_450),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_459),
.A2(n_418),
.B1(n_393),
.B2(n_395),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_487),
.Y(n_544)
);

AO32x1_ASAP7_75t_L g545 ( 
.A1(n_488),
.A2(n_417),
.A3(n_413),
.B1(n_409),
.B2(n_405),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_R g546 ( 
.A(n_444),
.B(n_29),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_493),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_453),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_470),
.B(n_31),
.Y(n_549)
);

A2O1A1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_504),
.A2(n_431),
.B(n_403),
.C(n_34),
.Y(n_550)
);

O2A1O1Ixp33_ASAP7_75t_SL g551 ( 
.A1(n_484),
.A2(n_113),
.B(n_167),
.C(n_163),
.Y(n_551)
);

AO32x1_ASAP7_75t_L g552 ( 
.A1(n_461),
.A2(n_403),
.A3(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_464),
.A2(n_112),
.B(n_161),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_453),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_502),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_502),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_443),
.B(n_37),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_458),
.A2(n_38),
.B1(n_44),
.B2(n_46),
.Y(n_558)
);

BUFx5_ASAP7_75t_L g559 ( 
.A(n_473),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_481),
.B(n_48),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_469),
.A2(n_50),
.B(n_52),
.Y(n_561)
);

A2O1A1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_506),
.A2(n_53),
.B(n_54),
.C(n_56),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_502),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_499),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_482),
.B(n_64),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_502),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_452),
.A2(n_67),
.B(n_70),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_474),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_507),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_503),
.A2(n_72),
.B(n_74),
.C(n_77),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_483),
.Y(n_572)
);

NAND2x1p5_ASAP7_75t_L g573 ( 
.A(n_455),
.B(n_457),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_462),
.B(n_162),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_463),
.B(n_85),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_498),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_94),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_503),
.A2(n_101),
.B(n_104),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_492),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_498),
.B(n_106),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_L g581 ( 
.A(n_525),
.B(n_446),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_515),
.A2(n_513),
.B(n_514),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_519),
.A2(n_111),
.B(n_116),
.Y(n_584)
);

INVx8_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_522),
.A2(n_119),
.B(n_122),
.Y(n_586)
);

AO32x2_ASAP7_75t_L g587 ( 
.A1(n_512),
.A2(n_552),
.A3(n_563),
.B1(n_543),
.B2(n_534),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_509),
.B(n_132),
.Y(n_588)
);

BUFx12f_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

BUFx4f_ASAP7_75t_L g590 ( 
.A(n_540),
.Y(n_590)
);

AO32x2_ASAP7_75t_L g591 ( 
.A1(n_552),
.A2(n_136),
.A3(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_591)
);

NAND3x1_ASAP7_75t_L g592 ( 
.A(n_518),
.B(n_142),
.C(n_145),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_542),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_523),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_531),
.B(n_156),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_546),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_520),
.A2(n_511),
.B(n_538),
.Y(n_597)
);

NOR2x1_ASAP7_75t_SL g598 ( 
.A(n_555),
.B(n_556),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_568),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_510),
.B(n_521),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_524),
.B(n_557),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_529),
.A2(n_533),
.B(n_535),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_569),
.Y(n_603)
);

AO31x2_ASAP7_75t_L g604 ( 
.A1(n_550),
.A2(n_577),
.A3(n_570),
.B(n_562),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_569),
.B(n_530),
.Y(n_605)
);

AO31x2_ASAP7_75t_L g606 ( 
.A1(n_567),
.A2(n_561),
.A3(n_553),
.B(n_560),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_566),
.A2(n_558),
.B(n_565),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_579),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_528),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_547),
.B(n_554),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_558),
.A2(n_575),
.B(n_574),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_547),
.B(n_573),
.Y(n_613)
);

NAND2x1_ASAP7_75t_L g614 ( 
.A(n_571),
.B(n_572),
.Y(n_614)
);

OA21x2_ASAP7_75t_L g615 ( 
.A1(n_536),
.A2(n_576),
.B(n_545),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_564),
.B(n_541),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_571),
.Y(n_617)
);

NOR2x1_ASAP7_75t_SL g618 ( 
.A(n_580),
.B(n_559),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_545),
.A2(n_539),
.B(n_551),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_559),
.B(n_537),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_559),
.Y(n_622)
);

OAI21xp33_ASAP7_75t_SL g623 ( 
.A1(n_559),
.A2(n_552),
.B(n_545),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_508),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_517),
.B(n_442),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_516),
.Y(n_626)
);

AO21x1_ASAP7_75t_L g627 ( 
.A1(n_527),
.A2(n_580),
.B(n_578),
.Y(n_627)
);

INVx3_ASAP7_75t_SL g628 ( 
.A(n_540),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_517),
.B(n_460),
.Y(n_629)
);

AOI221xp5_ASAP7_75t_SL g630 ( 
.A1(n_544),
.A2(n_477),
.B1(n_419),
.B2(n_451),
.C(n_472),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_517),
.B(n_442),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_555),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_517),
.B(n_442),
.Y(n_634)
);

BUFx6f_ASAP7_75t_SL g635 ( 
.A(n_518),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_517),
.B(n_442),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_517),
.A2(n_448),
.B(n_383),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_508),
.B(n_460),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_508),
.Y(n_639)
);

OA21x2_ASAP7_75t_L g640 ( 
.A1(n_527),
.A2(n_526),
.B(n_445),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_516),
.Y(n_641)
);

AND3x4_ASAP7_75t_L g642 ( 
.A(n_518),
.B(n_397),
.C(n_446),
.Y(n_642)
);

AO21x2_ASAP7_75t_L g643 ( 
.A1(n_527),
.A2(n_519),
.B(n_522),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_517),
.A2(n_448),
.B(n_383),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_540),
.Y(n_645)
);

CKINVDCx11_ASAP7_75t_R g646 ( 
.A(n_540),
.Y(n_646)
);

AO31x2_ASAP7_75t_L g647 ( 
.A1(n_527),
.A2(n_513),
.A3(n_522),
.B(n_550),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_517),
.A2(n_448),
.B(n_383),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_516),
.Y(n_649)
);

OA22x2_ASAP7_75t_L g650 ( 
.A1(n_508),
.A2(n_388),
.B1(n_371),
.B2(n_447),
.Y(n_650)
);

OAI21xp33_ASAP7_75t_L g651 ( 
.A1(n_517),
.A2(n_460),
.B(n_544),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_516),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_517),
.A2(n_448),
.B(n_383),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_516),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_517),
.B(n_388),
.Y(n_655)
);

CKINVDCx8_ASAP7_75t_R g656 ( 
.A(n_540),
.Y(n_656)
);

BUFx12f_ASAP7_75t_L g657 ( 
.A(n_508),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_532),
.A2(n_549),
.B(n_517),
.C(n_544),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_516),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_508),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_517),
.B(n_442),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_540),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_517),
.A2(n_448),
.B(n_383),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_517),
.B(n_460),
.Y(n_664)
);

OAI21x1_ASAP7_75t_SL g665 ( 
.A1(n_578),
.A2(n_491),
.B(n_558),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_516),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_517),
.B(n_442),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_631),
.Y(n_668)
);

CKINVDCx8_ASAP7_75t_R g669 ( 
.A(n_585),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_612),
.A2(n_583),
.B(n_597),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_620),
.A2(n_602),
.B(n_607),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_629),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_655),
.B(n_664),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_646),
.Y(n_674)
);

CKINVDCx8_ASAP7_75t_R g675 ( 
.A(n_585),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_590),
.Y(n_676)
);

NAND2x1p5_ASAP7_75t_L g677 ( 
.A(n_590),
.B(n_645),
.Y(n_677)
);

BUFx8_ASAP7_75t_L g678 ( 
.A(n_635),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_641),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_634),
.B(n_636),
.Y(n_680)
);

OAI21xp33_ASAP7_75t_SL g681 ( 
.A1(n_595),
.A2(n_621),
.B(n_600),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_661),
.B(n_667),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_588),
.A2(n_643),
.B(n_640),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_660),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_593),
.Y(n_685)
);

INVx6_ASAP7_75t_L g686 ( 
.A(n_645),
.Y(n_686)
);

AO31x2_ASAP7_75t_L g687 ( 
.A1(n_618),
.A2(n_584),
.A3(n_586),
.B(n_598),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_626),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_581),
.B(n_628),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_640),
.A2(n_663),
.B(n_653),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_656),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_637),
.A2(n_644),
.B(n_648),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_639),
.B(n_624),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_589),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_651),
.B(n_632),
.Y(n_695)
);

OAI21x1_ASAP7_75t_SL g696 ( 
.A1(n_618),
.A2(n_598),
.B(n_665),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_649),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_594),
.B(n_601),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_652),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_654),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_659),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_635),
.Y(n_702)
);

NAND2x1p5_ASAP7_75t_L g703 ( 
.A(n_582),
.B(n_662),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_666),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_599),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_609),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_630),
.B(n_610),
.Y(n_707)
);

AOI21xp33_ASAP7_75t_L g708 ( 
.A1(n_623),
.A2(n_650),
.B(n_615),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_622),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_657),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_619),
.A2(n_605),
.B(n_592),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_614),
.A2(n_613),
.B(n_611),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_617),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_647),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_616),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_638),
.B(n_603),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_604),
.B(n_647),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_642),
.B(n_596),
.Y(n_718)
);

INVx5_ASAP7_75t_L g719 ( 
.A(n_633),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_608),
.Y(n_720)
);

NOR2x1_ASAP7_75t_R g721 ( 
.A(n_591),
.B(n_587),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_587),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_591),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_606),
.B(n_625),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_650),
.A2(n_525),
.B1(n_655),
.B2(n_581),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_629),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_629),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_620),
.A2(n_665),
.B(n_627),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_629),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_635),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_629),
.Y(n_731)
);

INVx6_ASAP7_75t_L g732 ( 
.A(n_585),
.Y(n_732)
);

OAI21x1_ASAP7_75t_SL g733 ( 
.A1(n_618),
.A2(n_598),
.B(n_665),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_622),
.B(n_460),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_645),
.B(n_664),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_658),
.A2(n_644),
.B(n_637),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_645),
.B(n_664),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_629),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_625),
.B(n_631),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_695),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_695),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_724),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_696),
.B(n_733),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_685),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_688),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_697),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_693),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_714),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_673),
.B(n_672),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_699),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_700),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_701),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_725),
.A2(n_668),
.B1(n_739),
.B2(n_680),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_704),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_705),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_726),
.B(n_727),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_707),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_684),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_707),
.Y(n_759)
);

AO21x2_ASAP7_75t_L g760 ( 
.A1(n_670),
.A2(n_692),
.B(n_736),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_686),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_706),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_729),
.B(n_731),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_738),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_692),
.A2(n_736),
.B(n_683),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_681),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_735),
.Y(n_767)
);

OAI21x1_ASAP7_75t_SL g768 ( 
.A1(n_711),
.A2(n_668),
.B(n_739),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_737),
.B(n_715),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_681),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_737),
.B(n_698),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_717),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_679),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_719),
.Y(n_774)
);

AO21x2_ASAP7_75t_L g775 ( 
.A1(n_690),
.A2(n_671),
.B(n_708),
.Y(n_775)
);

INVx3_ASAP7_75t_SL g776 ( 
.A(n_732),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_723),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_680),
.B(n_682),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_722),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_709),
.B(n_708),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_721),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_721),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_669),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_728),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_720),
.B(n_719),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_719),
.B(n_712),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_779),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_742),
.B(n_728),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_786),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_753),
.A2(n_718),
.B1(n_678),
.B2(n_689),
.Y(n_790)
);

AOI33xp33_ASAP7_75t_L g791 ( 
.A1(n_744),
.A2(n_710),
.A3(n_713),
.B1(n_676),
.B2(n_678),
.B3(n_730),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_781),
.A2(n_730),
.B1(n_734),
.B2(n_716),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_748),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_781),
.B(n_703),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_766),
.B(n_687),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_757),
.B(n_686),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_770),
.B(n_677),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_757),
.B(n_702),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_770),
.B(n_674),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_772),
.B(n_732),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_749),
.B(n_675),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_782),
.B(n_694),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_782),
.B(n_691),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_780),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_786),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_740),
.B(n_741),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_760),
.B(n_777),
.Y(n_807)
);

BUFx2_ASAP7_75t_SL g808 ( 
.A(n_774),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_743),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_778),
.B(n_747),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_760),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_760),
.B(n_777),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_788),
.B(n_765),
.Y(n_813)
);

AND2x4_ASAP7_75t_SL g814 ( 
.A(n_797),
.B(n_743),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_809),
.B(n_784),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_788),
.B(n_765),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_788),
.B(n_807),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_787),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_807),
.B(n_765),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_804),
.B(n_764),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_793),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_812),
.B(n_775),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_810),
.B(n_762),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_804),
.B(n_759),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_805),
.B(n_759),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_793),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_810),
.B(n_752),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_806),
.B(n_752),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_805),
.B(n_758),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_823),
.B(n_799),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_820),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_817),
.B(n_809),
.Y(n_832)
);

AND2x4_ASAP7_75t_SL g833 ( 
.A(n_815),
.B(n_797),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_820),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_829),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_818),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_819),
.B(n_807),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_829),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_827),
.A2(n_799),
.B1(n_801),
.B2(n_790),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_824),
.B(n_812),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_824),
.B(n_789),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_819),
.B(n_795),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_825),
.B(n_813),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_813),
.B(n_795),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_828),
.B(n_799),
.Y(n_845)
);

AND3x1_ASAP7_75t_L g846 ( 
.A(n_816),
.B(n_791),
.C(n_803),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_833),
.Y(n_847)
);

OAI21xp33_ASAP7_75t_SL g848 ( 
.A1(n_843),
.A2(n_826),
.B(n_821),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_836),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_837),
.B(n_816),
.Y(n_850)
);

NAND4xp25_ASAP7_75t_L g851 ( 
.A(n_839),
.B(n_792),
.C(n_802),
.D(n_798),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_833),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_837),
.B(n_822),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_846),
.B(n_802),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_842),
.B(n_822),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_832),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_835),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_838),
.B(n_803),
.Y(n_858)
);

OAI22xp33_ASAP7_75t_L g859 ( 
.A1(n_854),
.A2(n_841),
.B1(n_840),
.B2(n_843),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_848),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_857),
.B(n_842),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_856),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_853),
.B(n_844),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_851),
.B(n_798),
.C(n_763),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_855),
.B(n_844),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_853),
.B(n_840),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_849),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_SL g868 ( 
.A1(n_847),
.A2(n_841),
.B(n_845),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_849),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_852),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_860),
.A2(n_856),
.B1(n_858),
.B2(n_855),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_859),
.A2(n_814),
.B(n_830),
.Y(n_872)
);

AOI211xp5_ASAP7_75t_L g873 ( 
.A1(n_859),
.A2(n_776),
.B(n_783),
.C(n_834),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_870),
.A2(n_850),
.B1(n_814),
.B2(n_832),
.Y(n_874)
);

OAI21xp33_ASAP7_75t_L g875 ( 
.A1(n_868),
.A2(n_850),
.B(n_831),
.Y(n_875)
);

OAI211xp5_ASAP7_75t_L g876 ( 
.A1(n_873),
.A2(n_870),
.B(n_864),
.C(n_783),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_875),
.B(n_871),
.Y(n_877)
);

OAI21xp33_ASAP7_75t_L g878 ( 
.A1(n_872),
.A2(n_862),
.B(n_861),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_877),
.B(n_863),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_876),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_880),
.B(n_776),
.Y(n_881)
);

NAND4xp25_ASAP7_75t_L g882 ( 
.A(n_879),
.B(n_878),
.C(n_874),
.D(n_769),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_881),
.A2(n_862),
.B1(n_863),
.B2(n_869),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_882),
.B(n_866),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_884),
.B(n_867),
.Y(n_885)
);

AND3x1_ASAP7_75t_L g886 ( 
.A(n_883),
.B(n_761),
.C(n_800),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_885),
.Y(n_887)
);

NAND4xp75_ASAP7_75t_L g888 ( 
.A(n_886),
.B(n_761),
.C(n_776),
.D(n_785),
.Y(n_888)
);

AOI31xp33_ASAP7_75t_L g889 ( 
.A1(n_885),
.A2(n_794),
.A3(n_756),
.B(n_771),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_887),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_888),
.B(n_774),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_889),
.A2(n_800),
.B1(n_865),
.B2(n_794),
.Y(n_892)
);

AO22x2_ASAP7_75t_L g893 ( 
.A1(n_887),
.A2(n_762),
.B1(n_744),
.B2(n_745),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_887),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_894),
.B(n_832),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_890),
.A2(n_796),
.B(n_785),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_891),
.A2(n_800),
.B1(n_808),
.B2(n_811),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_893),
.Y(n_898)
);

AO221x1_ASAP7_75t_L g899 ( 
.A1(n_892),
.A2(n_774),
.B1(n_768),
.B2(n_746),
.C(n_745),
.Y(n_899)
);

OAI21xp33_ASAP7_75t_L g900 ( 
.A1(n_890),
.A2(n_796),
.B(n_767),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_890),
.A2(n_751),
.B(n_746),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_895),
.B(n_750),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_896),
.B(n_750),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_898),
.A2(n_751),
.B(n_755),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_901),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_905),
.A2(n_900),
.B(n_899),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_904),
.B(n_897),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_L g908 ( 
.A1(n_903),
.A2(n_754),
.B1(n_755),
.B2(n_774),
.C(n_773),
.Y(n_908)
);

BUFx24_ASAP7_75t_SL g909 ( 
.A(n_906),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_909),
.A2(n_907),
.B1(n_902),
.B2(n_908),
.Y(n_910)
);


endmodule