module fake_jpeg_2693_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_44),
.B(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx11_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_77),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_78),
.Y(n_89)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_59),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_6),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_39),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_40),
.A3(n_52),
.B1(n_41),
.B2(n_42),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_60),
.B1(n_59),
.B2(n_45),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_57),
.B1(n_45),
.B2(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_40),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_47),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_53),
.B(n_51),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_92),
.B(n_24),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_1),
.C(n_2),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_101),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_17),
.B1(n_36),
.B2(n_35),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_99),
.B1(n_76),
.B2(n_10),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_7),
.CI(n_8),
.CON(n_101),
.SN(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_9),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_25),
.B1(n_34),
.B2(n_33),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_116),
.Y(n_128)
);

NOR4xp25_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_21),
.C(n_30),
.D(n_31),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_12),
.B(n_13),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_13),
.B(n_32),
.C(n_37),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_28),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_114),
.C(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_90),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_23),
.B1(n_14),
.B2(n_16),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_108),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_106),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_112),
.C(n_109),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_140),
.B(n_141),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_132),
.C(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_143),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_131),
.B1(n_126),
.B2(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_140),
.B(n_127),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_123),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_144),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_138),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_134),
.B(n_137),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_120),
.C(n_122),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_122),
.Y(n_153)
);


endmodule