module real_aes_2279_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g522 ( .A(n_0), .B(n_219), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_1), .B(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g153 ( .A(n_3), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_4), .B(n_525), .Y(n_544) );
NAND2xp33_ASAP7_75t_SL g515 ( .A(n_5), .B(n_174), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_6), .B(n_187), .Y(n_210) );
INVx1_ASAP7_75t_L g507 ( .A(n_7), .Y(n_507) );
INVx1_ASAP7_75t_L g244 ( .A(n_8), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_9), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_10), .Y(n_261) );
AND2x2_ASAP7_75t_L g542 ( .A(n_11), .B(n_143), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_12), .A2(n_101), .B1(n_103), .B2(n_112), .Y(n_100) );
INVx2_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_14), .B(n_109), .C(n_111), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_14), .Y(n_121) );
INVx1_ASAP7_75t_L g220 ( .A(n_15), .Y(n_220) );
AOI221x1_ASAP7_75t_L g510 ( .A1(n_16), .A2(n_176), .B1(n_511), .B2(n_513), .C(n_514), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_17), .B(n_525), .Y(n_578) );
NOR2xp33_ASAP7_75t_SL g105 ( .A(n_18), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g125 ( .A(n_18), .Y(n_125) );
INVx1_ASAP7_75t_L g217 ( .A(n_19), .Y(n_217) );
INVx1_ASAP7_75t_SL g165 ( .A(n_20), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_21), .B(n_168), .Y(n_190) );
AOI33xp33_ASAP7_75t_L g235 ( .A1(n_22), .A2(n_50), .A3(n_150), .B1(n_161), .B2(n_236), .B3(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_23), .A2(n_513), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_24), .B(n_219), .Y(n_547) );
AOI221xp5_ASAP7_75t_SL g587 ( .A1(n_25), .A2(n_40), .B1(n_513), .B2(n_525), .C(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g254 ( .A(n_26), .Y(n_254) );
OR2x2_ASAP7_75t_L g145 ( .A(n_27), .B(n_88), .Y(n_145) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_27), .A2(n_88), .B(n_144), .Y(n_178) );
INVxp67_ASAP7_75t_L g509 ( .A(n_28), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_29), .B(n_222), .Y(n_582) );
AND2x2_ASAP7_75t_L g536 ( .A(n_30), .B(n_142), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_31), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_32), .A2(n_513), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_33), .B(n_222), .Y(n_589) );
AND2x2_ASAP7_75t_L g155 ( .A(n_34), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g160 ( .A(n_34), .Y(n_160) );
AND2x2_ASAP7_75t_L g174 ( .A(n_34), .B(n_153), .Y(n_174) );
INVxp67_ASAP7_75t_L g111 ( .A(n_35), .Y(n_111) );
OR2x6_ASAP7_75t_L g123 ( .A(n_35), .B(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_36), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_37), .B(n_148), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_38), .A2(n_177), .B1(n_183), .B2(n_187), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_39), .B(n_192), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_41), .A2(n_80), .B1(n_158), .B2(n_513), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_42), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_43), .B(n_219), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_44), .A2(n_789), .B1(n_791), .B2(n_793), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_45), .B(n_194), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_46), .B(n_168), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_47), .Y(n_186) );
AND2x2_ASAP7_75t_L g526 ( .A(n_48), .B(n_142), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_49), .B(n_142), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_51), .B(n_168), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_52), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_52), .A2(n_62), .B1(n_433), .B2(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g151 ( .A(n_53), .Y(n_151) );
INVx1_ASAP7_75t_L g170 ( .A(n_53), .Y(n_170) );
AND2x2_ASAP7_75t_L g286 ( .A(n_54), .B(n_142), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_55), .A2(n_73), .B1(n_148), .B2(n_158), .C(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_56), .B(n_148), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_57), .B(n_525), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_58), .B(n_177), .Y(n_263) );
AOI21xp5_ASAP7_75t_SL g199 ( .A1(n_59), .A2(n_158), .B(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g563 ( .A(n_60), .B(n_142), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_61), .B(n_222), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_62), .Y(n_808) );
INVx1_ASAP7_75t_L g213 ( .A(n_63), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_64), .B(n_219), .Y(n_561) );
AND2x2_ASAP7_75t_SL g583 ( .A(n_65), .B(n_143), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_66), .A2(n_513), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g284 ( .A(n_67), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_68), .B(n_222), .Y(n_548) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_69), .B(n_194), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_70), .A2(n_158), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g156 ( .A(n_71), .Y(n_156) );
INVx1_ASAP7_75t_L g172 ( .A(n_71), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_72), .B(n_148), .Y(n_238) );
AND2x2_ASAP7_75t_L g175 ( .A(n_74), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g214 ( .A(n_75), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_76), .A2(n_158), .B(n_164), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_77), .A2(n_158), .B(n_189), .C(n_193), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_78), .A2(n_83), .B1(n_148), .B2(n_525), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_79), .B(n_525), .Y(n_562) );
INVx1_ASAP7_75t_L g106 ( .A(n_81), .Y(n_106) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_82), .B(n_176), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_84), .A2(n_158), .B1(n_233), .B2(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_85), .B(n_219), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_86), .B(n_219), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_87), .A2(n_513), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g201 ( .A(n_89), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_90), .B(n_222), .Y(n_560) );
AND2x2_ASAP7_75t_L g239 ( .A(n_91), .B(n_176), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_92), .A2(n_252), .B(n_253), .C(n_255), .Y(n_251) );
INVxp67_ASAP7_75t_L g512 ( .A(n_93), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_94), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_95), .B(n_222), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_96), .A2(n_513), .B(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g116 ( .A(n_97), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_98), .B(n_168), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_99), .Y(n_789) );
BUFx4f_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_106), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_127), .B(n_797), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_115), .B(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_118), .A2(n_799), .B(n_809), .Y(n_798) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_126), .Y(n_118) );
BUFx2_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g809 ( .A(n_120), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x6_ASAP7_75t_SL g497 ( .A(n_121), .B(n_123), .Y(n_497) );
OR2x6_ASAP7_75t_SL g788 ( .A(n_121), .B(n_122), .Y(n_788) );
OR2x2_ASAP7_75t_L g796 ( .A(n_121), .B(n_123), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_789), .B(n_790), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_496), .B1(n_498), .B2(n_786), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_131), .A2(n_496), .B1(n_499), .B2(n_792), .Y(n_791) );
AND3x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_490), .C(n_493), .Y(n_131) );
NAND5xp2_ASAP7_75t_L g132 ( .A(n_133), .B(n_390), .C(n_420), .D(n_434), .E(n_460), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_134), .A2(n_433), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g804 ( .A(n_134), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_339), .Y(n_134) );
NOR3xp33_ASAP7_75t_SL g135 ( .A(n_136), .B(n_287), .C(n_321), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_204), .B(n_226), .C(n_265), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_179), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_139), .B(n_277), .Y(n_342) );
AND2x2_ASAP7_75t_L g429 ( .A(n_139), .B(n_207), .Y(n_429) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g225 ( .A(n_140), .B(n_196), .Y(n_225) );
INVx1_ASAP7_75t_L g267 ( .A(n_140), .Y(n_267) );
INVx2_ASAP7_75t_L g272 ( .A(n_140), .Y(n_272) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_140), .Y(n_300) );
INVx1_ASAP7_75t_L g314 ( .A(n_140), .Y(n_314) );
AND2x2_ASAP7_75t_L g318 ( .A(n_140), .B(n_209), .Y(n_318) );
AND2x2_ASAP7_75t_L g399 ( .A(n_140), .B(n_208), .Y(n_399) );
AO21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .B(n_175), .Y(n_140) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_141), .A2(n_530), .B(n_536), .Y(n_529) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_141), .A2(n_557), .B(n_563), .Y(n_556) );
AO21x2_ASAP7_75t_L g594 ( .A1(n_141), .A2(n_530), .B(n_536), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_142), .Y(n_141) );
OA21x2_ASAP7_75t_L g586 ( .A1(n_142), .A2(n_587), .B(n_591), .Y(n_586) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x4_ASAP7_75t_L g187 ( .A(n_144), .B(n_145), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_157), .Y(n_146) );
INVx1_ASAP7_75t_L g264 ( .A(n_148), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_148), .A2(n_158), .B1(n_506), .B2(n_508), .Y(n_505) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_154), .Y(n_148) );
INVx1_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
OR2x6_ASAP7_75t_L g166 ( .A(n_150), .B(n_162), .Y(n_166) );
INVxp33_ASAP7_75t_L g236 ( .A(n_150), .Y(n_236) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g163 ( .A(n_151), .B(n_153), .Y(n_163) );
AND2x4_ASAP7_75t_L g222 ( .A(n_151), .B(n_171), .Y(n_222) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x6_ASAP7_75t_L g513 ( .A(n_155), .B(n_163), .Y(n_513) );
INVx2_ASAP7_75t_L g162 ( .A(n_156), .Y(n_162) );
AND2x6_ASAP7_75t_L g219 ( .A(n_156), .B(n_169), .Y(n_219) );
INVxp67_ASAP7_75t_L g262 ( .A(n_158), .Y(n_262) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_163), .Y(n_158) );
NOR2x1p5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx1_ASAP7_75t_L g237 ( .A(n_161), .Y(n_237) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_173), .Y(n_164) );
INVx2_ASAP7_75t_L g192 ( .A(n_166), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_166), .A2(n_173), .B(n_201), .C(n_202), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_166), .A2(n_213), .B1(n_214), .B2(n_215), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g243 ( .A1(n_166), .A2(n_173), .B(n_244), .C(n_245), .Y(n_243) );
INVxp67_ASAP7_75t_L g252 ( .A(n_166), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g283 ( .A1(n_166), .A2(n_173), .B(n_284), .C(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g215 ( .A(n_168), .Y(n_215) );
AND2x4_ASAP7_75t_L g525 ( .A(n_168), .B(n_174), .Y(n_525) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_171), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_173), .A2(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_173), .B(n_187), .Y(n_223) );
INVx1_ASAP7_75t_L g233 ( .A(n_173), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_173), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_173), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_173), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_173), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_173), .A2(n_581), .B(n_582), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_173), .A2(n_589), .B(n_590), .Y(n_588) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_174), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_176), .A2(n_251), .B1(n_256), .B2(n_257), .Y(n_250) );
INVx3_ASAP7_75t_L g257 ( .A(n_176), .Y(n_257) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_177), .B(n_260), .Y(n_259) );
AOI21x1_ASAP7_75t_L g518 ( .A1(n_177), .A2(n_519), .B(n_526), .Y(n_518) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx4f_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
AND2x4_ASAP7_75t_SL g179 ( .A(n_180), .B(n_195), .Y(n_179) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g224 ( .A(n_181), .Y(n_224) );
AND2x2_ASAP7_75t_L g268 ( .A(n_181), .B(n_209), .Y(n_268) );
AND2x2_ASAP7_75t_L g289 ( .A(n_181), .B(n_196), .Y(n_289) );
INVx1_ASAP7_75t_L g312 ( .A(n_181), .Y(n_312) );
AND2x4_ASAP7_75t_L g379 ( .A(n_181), .B(n_208), .Y(n_379) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_188), .Y(n_181) );
NOR3xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .C(n_186), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_187), .A2(n_199), .B(n_203), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_187), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_187), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_187), .B(n_512), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_187), .B(n_215), .C(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_187), .A2(n_544), .B(n_545), .Y(n_543) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_193), .A2(n_231), .B(n_239), .Y(n_230) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_193), .A2(n_231), .B(n_239), .Y(n_294) );
AOI21x1_ASAP7_75t_L g551 ( .A1(n_193), .A2(n_552), .B(n_555), .Y(n_551) );
INVx2_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_194), .A2(n_242), .B(n_246), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_194), .A2(n_578), .B(n_579), .Y(n_577) );
AND2x4_ASAP7_75t_L g395 ( .A(n_195), .B(n_312), .Y(n_395) );
OR2x2_ASAP7_75t_L g436 ( .A(n_195), .B(n_437), .Y(n_436) );
NOR2xp67_ASAP7_75t_SL g455 ( .A(n_195), .B(n_328), .Y(n_455) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_195), .B(n_387), .Y(n_473) );
INVx4_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2x1_ASAP7_75t_SL g273 ( .A(n_196), .B(n_209), .Y(n_273) );
AND2x4_ASAP7_75t_L g311 ( .A(n_196), .B(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_196), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_196), .B(n_271), .Y(n_349) );
INVx2_ASAP7_75t_L g363 ( .A(n_196), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_196), .B(n_315), .Y(n_385) );
AND2x2_ASAP7_75t_L g477 ( .A(n_196), .B(n_335), .Y(n_477) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2x1_ASAP7_75t_L g205 ( .A(n_206), .B(n_225), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_207), .B(n_314), .Y(n_328) );
AND2x2_ASAP7_75t_SL g337 ( .A(n_207), .B(n_317), .Y(n_337) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_224), .Y(n_207) );
INVx1_ASAP7_75t_L g315 ( .A(n_208), .Y(n_315) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g335 ( .A(n_209), .Y(n_335) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_216), .B(n_223), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_215), .B(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B1(n_220), .B2(n_221), .Y(n_216) );
INVxp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVxp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g368 ( .A(n_224), .Y(n_368) );
INVx2_ASAP7_75t_SL g413 ( .A(n_225), .Y(n_413) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_247), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_228), .B(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g359 ( .A(n_228), .Y(n_359) );
AND2x2_ASAP7_75t_L g483 ( .A(n_228), .B(n_308), .Y(n_483) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_240), .Y(n_228) );
AND2x4_ASAP7_75t_L g296 ( .A(n_229), .B(n_278), .Y(n_296) );
INVx1_ASAP7_75t_L g307 ( .A(n_229), .Y(n_307) );
AND2x2_ASAP7_75t_L g338 ( .A(n_229), .B(n_293), .Y(n_338) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_230), .B(n_241), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_230), .B(n_279), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_232), .B(n_238), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVxp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g276 ( .A(n_241), .Y(n_276) );
AND2x4_ASAP7_75t_L g344 ( .A(n_241), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g356 ( .A(n_241), .Y(n_356) );
INVx1_ASAP7_75t_L g398 ( .A(n_241), .Y(n_398) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_241), .Y(n_410) );
AND2x2_ASAP7_75t_L g426 ( .A(n_241), .B(n_249), .Y(n_426) );
BUFx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g373 ( .A(n_248), .B(n_331), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_248), .Y(n_375) );
AND2x2_ASAP7_75t_L g396 ( .A(n_248), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g275 ( .A(n_249), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g303 ( .A(n_249), .Y(n_303) );
INVx2_ASAP7_75t_L g309 ( .A(n_249), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_249), .B(n_279), .Y(n_324) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_258), .Y(n_249) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_257), .A2(n_280), .B(n_286), .Y(n_279) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_257), .A2(n_280), .B(n_286), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B1(n_263), .B2(n_264), .Y(n_258) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .B(n_274), .Y(n_265) );
INVx1_ASAP7_75t_L g405 ( .A(n_266), .Y(n_405) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g325 ( .A(n_268), .Y(n_325) );
AND2x2_ASAP7_75t_L g381 ( .A(n_268), .B(n_317), .Y(n_381) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
INVx1_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_270), .B(n_311), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_270), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g402 ( .A(n_270), .B(n_395), .Y(n_402) );
AND2x2_ASAP7_75t_L g476 ( .A(n_270), .B(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_271), .Y(n_464) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_272), .Y(n_384) );
AND2x2_ASAP7_75t_L g297 ( .A(n_273), .B(n_298), .Y(n_297) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_273), .A2(n_486), .B(n_488), .Y(n_485) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx3_ASAP7_75t_L g371 ( .A(n_275), .Y(n_371) );
NAND2x1_ASAP7_75t_SL g415 ( .A(n_275), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g418 ( .A(n_275), .B(n_296), .Y(n_418) );
AND2x2_ASAP7_75t_L g330 ( .A(n_277), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g467 ( .A(n_277), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g478 ( .A(n_277), .B(n_426), .Y(n_478) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_278), .B(n_355), .Y(n_354) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g409 ( .A(n_279), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_301), .B(n_304), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B1(n_296), .B2(n_297), .Y(n_288) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_289), .Y(n_346) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g425 ( .A(n_291), .B(n_426), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_291), .A2(n_444), .B1(n_445), .B2(n_446), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_291), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_293), .B(n_309), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g389 ( .A(n_293), .B(n_309), .Y(n_389) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_293), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g345 ( .A(n_294), .Y(n_345) );
AND2x2_ASAP7_75t_L g353 ( .A(n_294), .B(n_309), .Y(n_353) );
INVx1_ASAP7_75t_L g416 ( .A(n_294), .Y(n_416) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2x1_ASAP7_75t_L g334 ( .A(n_299), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g446 ( .A(n_302), .B(n_331), .Y(n_446) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
AND2x2_ASAP7_75t_L g343 ( .A(n_303), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g431 ( .A(n_303), .B(n_338), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_310), .B1(n_316), .B2(n_319), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g439 ( .A(n_306), .B(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g469 ( .A(n_309), .B(n_356), .Y(n_469) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx2_ASAP7_75t_L g336 ( .A(n_311), .Y(n_336) );
OAI21xp33_ASAP7_75t_SL g482 ( .A1(n_311), .A2(n_483), .B(n_484), .Y(n_482) );
AND2x4_ASAP7_75t_SL g313 ( .A(n_314), .B(n_315), .Y(n_313) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_314), .Y(n_472) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_SL g414 ( .A1(n_317), .A2(n_415), .B(n_417), .C(n_419), .Y(n_414) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_318), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g419 ( .A(n_318), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_318), .B(n_395), .Y(n_459) );
INVx1_ASAP7_75t_SL g326 ( .A(n_319), .Y(n_326) );
AND2x2_ASAP7_75t_L g407 ( .A(n_320), .B(n_344), .Y(n_407) );
INVx1_ASAP7_75t_L g452 ( .A(n_320), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B1(n_326), .B2(n_327), .C(n_329), .Y(n_321) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_322), .Y(n_441) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g489 ( .A(n_324), .B(n_332), .Y(n_489) );
OR2x2_ASAP7_75t_L g348 ( .A(n_325), .B(n_349), .Y(n_348) );
NOR2x1_ASAP7_75t_L g361 ( .A(n_325), .B(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_325), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g487 ( .A(n_325), .B(n_384), .Y(n_487) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI32xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .A3(n_336), .B1(n_337), .B2(n_338), .Y(n_329) );
INVx1_ASAP7_75t_L g350 ( .A(n_331), .Y(n_350) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_333), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g445 ( .A(n_334), .Y(n_445) );
OAI22xp33_ASAP7_75t_SL g427 ( .A1(n_336), .A2(n_428), .B1(n_430), .B2(n_432), .Y(n_427) );
INVx1_ASAP7_75t_L g458 ( .A(n_337), .Y(n_458) );
AOI211x1_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_346), .B(n_347), .C(n_364), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_341), .B(n_426), .Y(n_432) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g388 ( .A(n_344), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g454 ( .A(n_344), .Y(n_454) );
OAI222xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B1(n_351), .B2(n_357), .C1(n_358), .C2(n_360), .Y(n_347) );
INVxp67_ASAP7_75t_L g444 ( .A(n_348), .Y(n_444) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_352), .B(n_437), .Y(n_484) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g400 ( .A(n_353), .B(n_397), .Y(n_400) );
INVx3_ASAP7_75t_L g440 ( .A(n_355), .Y(n_440) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g378 ( .A(n_363), .B(n_379), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B1(n_372), .B2(n_377), .C(n_380), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_366), .A2(n_423), .B(n_425), .Y(n_422) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g376 ( .A(n_370), .Y(n_376) );
OR2x2_ASAP7_75t_L g480 ( .A(n_371), .B(n_416), .Y(n_480) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_374), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_377), .A2(n_406), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_378), .A2(n_450), .B(n_457), .Y(n_456) );
INVx4_ASAP7_75t_L g387 ( .A(n_379), .Y(n_387) );
OAI31xp33_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_382), .A3(n_386), .B(n_388), .Y(n_380) );
INVx1_ASAP7_75t_L g438 ( .A(n_382), .Y(n_438) );
NOR2x1_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g412 ( .A(n_387), .Y(n_412) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_403), .Y(n_390) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_391), .B(n_403), .C(n_422), .D(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_401), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_399), .B2(n_400), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g463 ( .A(n_395), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_396), .B(n_416), .Y(n_424) );
INVx1_ASAP7_75t_SL g437 ( .A(n_399), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_414), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_408), .B2(n_411), .Y(n_404) );
INVx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_413), .A2(n_476), .B1(n_478), .B2(n_479), .Y(n_475) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_427), .C(n_433), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g492 ( .A(n_427), .Y(n_492) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_433), .A2(n_494), .B(n_495), .Y(n_493) );
INVxp33_ASAP7_75t_L g494 ( .A(n_434), .Y(n_494) );
AND2x2_ASAP7_75t_L g803 ( .A(n_434), .B(n_460), .Y(n_803) );
NOR2xp67_ASAP7_75t_L g434 ( .A(n_435), .B(n_442), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B1(n_439), .B2(n_441), .Y(n_435) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_439), .A2(n_462), .B(n_465), .Y(n_461) );
INVx2_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_447), .C(n_456), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B1(n_453), .B2(n_455), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVxp33_ASAP7_75t_SL g495 ( .A(n_460), .Y(n_495) );
NOR3x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_474), .C(n_481), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_482), .B(n_485), .Y(n_481) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g805 ( .A(n_491), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_663), .Y(n_499) );
NOR4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_606), .C(n_645), .D(n_652), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_527), .B1(n_564), .B2(n_573), .C(n_592), .Y(n_501) );
OR2x2_ASAP7_75t_L g736 ( .A(n_502), .B(n_598), .Y(n_736) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g651 ( .A(n_503), .B(n_576), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_503), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_SL g716 ( .A(n_503), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_516), .Y(n_503) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_504), .B(n_576), .Y(n_575) );
INVx3_ASAP7_75t_L g597 ( .A(n_504), .Y(n_597) );
AND2x2_ASAP7_75t_L g632 ( .A(n_504), .B(n_605), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_504), .B(n_517), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_504), .B(n_599), .Y(n_684) );
OR2x2_ASAP7_75t_L g762 ( .A(n_504), .B(n_576), .Y(n_762) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .Y(n_504) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g584 ( .A(n_517), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_517), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g610 ( .A(n_517), .Y(n_610) );
OR2x2_ASAP7_75t_L g615 ( .A(n_517), .B(n_599), .Y(n_615) );
AND2x2_ASAP7_75t_L g628 ( .A(n_517), .B(n_586), .Y(n_628) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_517), .Y(n_631) );
INVx1_ASAP7_75t_L g643 ( .A(n_517), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_517), .B(n_597), .Y(n_708) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_528), .B(n_537), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g572 ( .A(n_529), .B(n_556), .Y(n_572) );
AND2x4_ASAP7_75t_L g602 ( .A(n_529), .B(n_541), .Y(n_602) );
INVx2_ASAP7_75t_L g636 ( .A(n_529), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_529), .B(n_556), .Y(n_694) );
AND2x2_ASAP7_75t_L g741 ( .A(n_529), .B(n_570), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g729 ( .A1(n_537), .A2(n_601), .B1(n_644), .B2(n_704), .C1(n_730), .C2(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_549), .Y(n_538) );
AND2x2_ASAP7_75t_L g648 ( .A(n_539), .B(n_568), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_539), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g777 ( .A(n_539), .B(n_617), .Y(n_777) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_540), .A2(n_608), .B(n_612), .Y(n_607) );
AND2x2_ASAP7_75t_L g688 ( .A(n_540), .B(n_571), .Y(n_688) );
OR2x2_ASAP7_75t_L g713 ( .A(n_540), .B(n_572), .Y(n_713) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx5_ASAP7_75t_L g567 ( .A(n_541), .Y(n_567) );
AND2x2_ASAP7_75t_L g654 ( .A(n_541), .B(n_636), .Y(n_654) );
AND2x2_ASAP7_75t_L g680 ( .A(n_541), .B(n_556), .Y(n_680) );
OR2x2_ASAP7_75t_L g683 ( .A(n_541), .B(n_570), .Y(n_683) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_541), .Y(n_701) );
AND2x4_ASAP7_75t_SL g758 ( .A(n_541), .B(n_635), .Y(n_758) );
OR2x2_ASAP7_75t_L g767 ( .A(n_541), .B(n_594), .Y(n_767) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g600 ( .A(n_549), .Y(n_600) );
AOI221xp5_ASAP7_75t_SL g718 ( .A1(n_549), .A2(n_602), .B1(n_719), .B2(n_721), .C(n_722), .Y(n_718) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_556), .Y(n_549) );
OR2x2_ASAP7_75t_L g657 ( .A(n_550), .B(n_627), .Y(n_657) );
OR2x2_ASAP7_75t_L g667 ( .A(n_550), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g693 ( .A(n_550), .B(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g699 ( .A(n_550), .B(n_618), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_550), .B(n_682), .Y(n_711) );
INVx2_ASAP7_75t_L g724 ( .A(n_550), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_550), .B(n_602), .Y(n_745) );
AND2x2_ASAP7_75t_L g749 ( .A(n_550), .B(n_571), .Y(n_749) );
AND2x2_ASAP7_75t_L g757 ( .A(n_550), .B(n_758), .Y(n_757) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g570 ( .A(n_551), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_556), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g601 ( .A(n_556), .B(n_570), .Y(n_601) );
INVx2_ASAP7_75t_L g618 ( .A(n_556), .Y(n_618) );
AND2x4_ASAP7_75t_L g635 ( .A(n_556), .B(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_556), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g747 ( .A(n_566), .B(n_569), .Y(n_747) );
AND2x4_ASAP7_75t_L g593 ( .A(n_567), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g634 ( .A(n_567), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g661 ( .A(n_567), .B(n_601), .Y(n_661) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g765 ( .A(n_569), .B(n_766), .Y(n_765) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g617 ( .A(n_570), .B(n_618), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_571), .A2(n_638), .B(n_644), .Y(n_637) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_584), .Y(n_574) );
INVx1_ASAP7_75t_SL g691 ( .A(n_575), .Y(n_691) );
AND2x2_ASAP7_75t_L g721 ( .A(n_575), .B(n_631), .Y(n_721) );
AND2x4_ASAP7_75t_L g732 ( .A(n_575), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g598 ( .A(n_576), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g605 ( .A(n_576), .Y(n_605) );
AND2x4_ASAP7_75t_L g611 ( .A(n_576), .B(n_597), .Y(n_611) );
INVx2_ASAP7_75t_L g622 ( .A(n_576), .Y(n_622) );
INVx1_ASAP7_75t_L g671 ( .A(n_576), .Y(n_671) );
OR2x2_ASAP7_75t_L g692 ( .A(n_576), .B(n_676), .Y(n_692) );
OR2x2_ASAP7_75t_L g706 ( .A(n_576), .B(n_586), .Y(n_706) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_576), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_576), .B(n_628), .Y(n_778) );
OR2x6_ASAP7_75t_L g576 ( .A(n_577), .B(n_583), .Y(n_576) );
INVx1_ASAP7_75t_L g623 ( .A(n_584), .Y(n_623) );
AND2x2_ASAP7_75t_L g756 ( .A(n_584), .B(n_622), .Y(n_756) );
AND2x2_ASAP7_75t_L g781 ( .A(n_584), .B(n_611), .Y(n_781) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g599 ( .A(n_586), .Y(n_599) );
BUFx3_ASAP7_75t_L g641 ( .A(n_586), .Y(n_641) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_586), .Y(n_668) );
INVx1_ASAP7_75t_L g677 ( .A(n_586), .Y(n_677) );
AOI33xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .A3(n_600), .B1(n_601), .B2(n_602), .B3(n_603), .Y(n_592) );
AOI21x1_ASAP7_75t_SL g695 ( .A1(n_593), .A2(n_617), .B(n_679), .Y(n_695) );
INVx2_ASAP7_75t_L g725 ( .A(n_593), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_593), .B(n_724), .Y(n_731) );
AND2x2_ASAP7_75t_L g679 ( .A(n_594), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AND2x2_ASAP7_75t_L g642 ( .A(n_597), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g743 ( .A(n_598), .Y(n_743) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_599), .Y(n_733) );
OAI32xp33_ASAP7_75t_L g782 ( .A1(n_600), .A2(n_602), .A3(n_778), .B1(n_783), .B2(n_785), .Y(n_782) );
AND2x2_ASAP7_75t_L g700 ( .A(n_601), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g690 ( .A(n_602), .Y(n_690) );
AND2x2_ASAP7_75t_L g755 ( .A(n_602), .B(n_699), .Y(n_755) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_616), .B1(n_619), .B2(n_633), .C(n_637), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_610), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_611), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_611), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_611), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g660 ( .A(n_615), .Y(n_660) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_624), .C(n_629), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_621), .A2(n_683), .B1(n_723), .B2(n_726), .Y(n_722) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g626 ( .A(n_622), .Y(n_626) );
NOR2x1p5_ASAP7_75t_L g640 ( .A(n_622), .B(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI322xp33_ASAP7_75t_L g689 ( .A1(n_625), .A2(n_667), .A3(n_690), .B1(n_691), .B2(n_692), .C1(n_693), .C2(n_695), .Y(n_689) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_627), .A2(n_646), .B(n_647), .C(n_649), .Y(n_645) );
OR2x2_ASAP7_75t_L g737 ( .A(n_627), .B(n_691), .Y(n_737) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g644 ( .A(n_628), .B(n_632), .Y(n_644) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g650 ( .A(n_634), .B(n_651), .Y(n_650) );
INVx3_ASAP7_75t_SL g682 ( .A(n_635), .Y(n_682) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_639), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_SL g686 ( .A(n_642), .Y(n_686) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_643), .Y(n_728) );
OR2x6_ASAP7_75t_SL g783 ( .A(n_646), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g773 ( .A1(n_651), .A2(n_774), .B(n_775), .C(n_782), .Y(n_773) );
O2A1O1Ixp33_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_655), .B(n_658), .C(n_662), .Y(n_652) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_653), .A2(n_665), .B(n_672), .C(n_696), .Y(n_664) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_709), .C(n_753), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_668), .Y(n_760) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g715 ( .A(n_671), .Y(n_715) );
NOR3xp33_ASAP7_75t_SL g672 ( .A(n_673), .B(n_685), .C(n_689), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_678), .B1(n_681), .B2(n_684), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g717 ( .A(n_677), .Y(n_717) );
INVxp67_ASAP7_75t_SL g784 ( .A(n_677), .Y(n_784) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_SL g770 ( .A(n_683), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
OR2x2_ASAP7_75t_L g720 ( .A(n_686), .B(n_706), .Y(n_720) );
OR2x2_ASAP7_75t_L g771 ( .A(n_686), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g769 ( .A(n_694), .Y(n_769) );
OR2x2_ASAP7_75t_L g785 ( .A(n_694), .B(n_724), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_700), .B(n_702), .Y(n_696) );
OAI31xp33_ASAP7_75t_L g710 ( .A1(n_697), .A2(n_711), .A3(n_712), .B(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g742 ( .A(n_707), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND4xp25_ASAP7_75t_SL g709 ( .A(n_710), .B(n_718), .C(n_729), .D(n_734), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_717), .Y(n_752) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_738), .B1(n_742), .B2(n_744), .C(n_746), .Y(n_734) );
NAND2xp33_ASAP7_75t_SL g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g779 ( .A(n_738), .Y(n_779) );
AND2x2_ASAP7_75t_SL g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g774 ( .A(n_748), .Y(n_774) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_773), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_757), .B2(n_759), .C(n_763), .Y(n_754) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
AOI21xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_768), .B(n_771), .Y(n_763) );
INVxp33_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_787), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OAI22xp33_ASAP7_75t_SL g799 ( .A1(n_800), .A2(n_801), .B1(n_806), .B2(n_807), .Y(n_799) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND3x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .C(n_805), .Y(n_802) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
endmodule