module fake_ariane_915_n_1405 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_1405);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_1405;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_96;
wire n_319;
wire n_49;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_72;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_57;
wire n_117;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_137;
wire n_1298;
wire n_1366;
wire n_232;
wire n_52;
wire n_568;
wire n_1088;
wire n_77;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_54;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_69;
wire n_259;
wire n_953;
wire n_1364;
wire n_143;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_93;
wire n_1074;
wire n_859;
wire n_108;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_136;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_104;
wire n_438;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_1391;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_94;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_65;
wire n_123;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_135;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_102;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_78;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_306;
wire n_92;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_111;
wire n_274;
wire n_1083;
wire n_967;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_76;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_80;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_124;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_133;
wire n_66;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_776;
wire n_424;
wire n_85;
wire n_130;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_138;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_73;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_59;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_90;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_120;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_129;
wire n_126;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_86;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_46;
wire n_84;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_70;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_61;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_55;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_134;
wire n_1257;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_211;
wire n_642;
wire n_97;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1305;
wire n_180;
wire n_64;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_71;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_87;
wire n_714;
wire n_790;
wire n_354;
wire n_140;
wire n_725;
wire n_151;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_75;
wire n_1047;
wire n_95;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_106;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_62;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_128;
wire n_224;
wire n_82;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_81;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_141;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_305;
wire n_312;
wire n_56;
wire n_60;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_89;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_74;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_107;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_58;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_125;
wire n_820;
wire n_43;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_99;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_67;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_114;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_132;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_121;
wire n_118;
wire n_353;
wire n_1361;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_828;
wire n_322;
wire n_1359;
wire n_558;
wire n_116;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_160;
wire n_119;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_109;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_50;
wire n_318;
wire n_103;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_139;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_122;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_47;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_115;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_79;
wire n_759;
wire n_567;
wire n_91;
wire n_240;
wire n_369;
wire n_44;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_48;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_88;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_53;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_68;
wire n_415;
wire n_63;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_83;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_110;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_98;
wire n_946;
wire n_757;
wire n_375;
wire n_113;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_156;
wire n_174;
wire n_275;
wire n_100;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_51;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_105;
wire n_1051;
wire n_719;
wire n_131;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_101;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_112;
wire n_45;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_127;
wire n_531;
wire n_1374;
wire n_675;

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_23),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_11),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_5),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_28),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_27),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_7),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_48),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_0),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_R g104 ( 
.A(n_87),
.B(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_91),
.B1(n_95),
.B2(n_65),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_R g134 ( 
.A(n_114),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_91),
.B1(n_95),
.B2(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_93),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_71),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_93),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_107),
.B(n_97),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_68),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_123),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

BUFx4f_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_99),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_116),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_115),
.A2(n_95),
.B1(n_68),
.B2(n_83),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_104),
.B(n_116),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_111),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_71),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_74),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_121),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_117),
.A2(n_80),
.B1(n_66),
.B2(n_74),
.Y(n_176)
);

CKINVDCx8_ASAP7_75t_R g177 ( 
.A(n_119),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_74),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_58),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_52),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_110),
.B(n_100),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_124),
.B(n_125),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_129),
.B(n_128),
.C(n_120),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_66),
.B1(n_80),
.B2(n_124),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_125),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_127),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_127),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_104),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_121),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_121),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_126),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_102),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_181),
.B1(n_166),
.B2(n_131),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_131),
.C(n_137),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_51),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_129),
.C(n_128),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_128),
.Y(n_213)
);

BUFx8_ASAP7_75t_SL g214 ( 
.A(n_136),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_129),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_144),
.A2(n_58),
.B(n_52),
.C(n_68),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_159),
.A2(n_52),
.B1(n_68),
.B2(n_83),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_148),
.B(n_130),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_154),
.B(n_102),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_159),
.A2(n_83),
.B1(n_62),
.B2(n_84),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_130),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_177),
.B(n_51),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_130),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_151),
.B(n_100),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_100),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_L g228 ( 
.A(n_159),
.B(n_134),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_157),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_151),
.B(n_101),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_159),
.A2(n_73),
.B1(n_72),
.B2(n_75),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_177),
.B(n_53),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_151),
.B(n_171),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_151),
.B(n_101),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_151),
.B(n_101),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_177),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_118),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_168),
.B(n_53),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_176),
.A2(n_118),
.B1(n_113),
.B2(n_55),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_159),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_180),
.B(n_113),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_180),
.A2(n_43),
.B1(n_45),
.B2(n_84),
.Y(n_248)
);

AND2x6_ASAP7_75t_SL g249 ( 
.A(n_178),
.B(n_70),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_151),
.B(n_103),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_61),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_176),
.A2(n_185),
.B1(n_136),
.B2(n_165),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_178),
.A2(n_70),
.B1(n_54),
.B2(n_46),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_180),
.B(n_61),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_168),
.B(n_59),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_163),
.A2(n_103),
.B(n_54),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_171),
.B(n_103),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_187),
.B(n_85),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_185),
.B(n_176),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_157),
.A2(n_77),
.B(n_55),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_182),
.Y(n_263)
);

NAND2x1_ASAP7_75t_L g264 ( 
.A(n_141),
.B(n_182),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_182),
.A2(n_76),
.B1(n_82),
.B2(n_81),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_187),
.B(n_85),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_171),
.B(n_77),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_L g269 ( 
.A(n_150),
.B(n_0),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_173),
.B(n_64),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_173),
.B(n_64),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_173),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_205),
.Y(n_274)
);

AO22x1_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_165),
.B1(n_173),
.B2(n_178),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_195),
.B(n_178),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_190),
.B(n_178),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_206),
.A2(n_186),
.B1(n_150),
.B2(n_152),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_205),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_204),
.Y(n_284)
);

OR2x6_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_186),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_190),
.B(n_135),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_195),
.B(n_178),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_204),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_192),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_203),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_203),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_234),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_190),
.B(n_135),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_207),
.A2(n_188),
.B1(n_135),
.B2(n_140),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_214),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_209),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_201),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_190),
.B(n_199),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_212),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_138),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_207),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_199),
.B(n_138),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_212),
.B(n_139),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_231),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_246),
.B(n_189),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_194),
.B(n_134),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_224),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_224),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_201),
.Y(n_318)
);

BUFx4f_ASAP7_75t_L g319 ( 
.A(n_237),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_189),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_239),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_SL g322 ( 
.A(n_253),
.B(n_59),
.C(n_60),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_152),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_196),
.B(n_132),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_197),
.B(n_132),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_233),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_217),
.B(n_132),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_233),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_230),
.B(n_140),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_230),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_SL g335 ( 
.A(n_247),
.B(n_56),
.C(n_60),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_238),
.B(n_155),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_261),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_263),
.B(n_139),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_267),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_SL g342 ( 
.A(n_252),
.B(n_56),
.C(n_78),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_270),
.B(n_188),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_189),
.B(n_186),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_189),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_227),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_267),
.B(n_150),
.Y(n_347)
);

BUFx4f_ASAP7_75t_L g348 ( 
.A(n_251),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_189),
.B(n_152),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_206),
.A2(n_164),
.B1(n_155),
.B2(n_79),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_215),
.B(n_164),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_SL g354 ( 
.A(n_281),
.B(n_189),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_284),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_351),
.A2(n_228),
.B(n_219),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_326),
.A2(n_219),
.B(n_257),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_351),
.A2(n_225),
.B(n_222),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_273),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_270),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_271),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_321),
.B(n_271),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g363 ( 
.A1(n_322),
.A2(n_260),
.B1(n_242),
.B2(n_248),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

AO21x2_ASAP7_75t_L g365 ( 
.A1(n_324),
.A2(n_269),
.B(n_191),
.Y(n_365)
);

AOI21x1_ASAP7_75t_SL g366 ( 
.A1(n_343),
.A2(n_211),
.B(n_213),
.Y(n_366)
);

AOI21x1_ASAP7_75t_L g367 ( 
.A1(n_280),
.A2(n_264),
.B(n_269),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_321),
.B(n_255),
.Y(n_368)
);

O2A1O1Ixp5_ASAP7_75t_L g369 ( 
.A1(n_314),
.A2(n_337),
.B(n_244),
.C(n_256),
.Y(n_369)
);

OAI211xp5_ASAP7_75t_L g370 ( 
.A1(n_342),
.A2(n_259),
.B(n_266),
.C(n_193),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_276),
.B(n_288),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_308),
.A2(n_163),
.B(n_264),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_295),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_278),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_277),
.B(n_227),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_338),
.A2(n_245),
.B1(n_220),
.B2(n_193),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_310),
.B(n_249),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_285),
.Y(n_379)
);

AO21x1_ASAP7_75t_L g380 ( 
.A1(n_280),
.A2(n_235),
.B(n_248),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_305),
.A2(n_210),
.B(n_202),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_305),
.A2(n_210),
.B(n_200),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g383 ( 
.A1(n_297),
.A2(n_184),
.B(n_149),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g384 ( 
.A1(n_297),
.A2(n_184),
.B(n_149),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_306),
.B(n_311),
.Y(n_385)
);

AOI21x1_ASAP7_75t_L g386 ( 
.A1(n_308),
.A2(n_184),
.B(n_153),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_198),
.B(n_163),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_302),
.B(n_258),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_322),
.A2(n_275),
.B1(n_342),
.B2(n_277),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_277),
.B(n_226),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_302),
.B(n_254),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_284),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_332),
.A2(n_340),
.B(n_347),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_332),
.A2(n_163),
.B(n_251),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_340),
.A2(n_184),
.B(n_133),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_313),
.B(n_251),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_323),
.A2(n_235),
.B1(n_232),
.B2(n_240),
.Y(n_398)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_331),
.A2(n_175),
.B(n_149),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_347),
.A2(n_163),
.B(n_250),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_282),
.B(n_318),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_323),
.B(n_275),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_319),
.A2(n_163),
.B(n_241),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_350),
.A2(n_169),
.B(n_133),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_306),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_313),
.B(n_208),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_286),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_282),
.B(n_249),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_343),
.B(n_268),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_331),
.A2(n_175),
.B(n_153),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_286),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_343),
.B(n_218),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_312),
.B(n_265),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_306),
.B(n_236),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_301),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_331),
.A2(n_156),
.B(n_149),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_301),
.B(n_304),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_306),
.B(n_223),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_286),
.A2(n_156),
.B(n_153),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_304),
.B(n_265),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_273),
.Y(n_421)
);

OAI21x1_ASAP7_75t_L g422 ( 
.A1(n_289),
.A2(n_169),
.B(n_153),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_304),
.B(n_262),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_307),
.B(n_262),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_319),
.A2(n_348),
.B(n_307),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_282),
.B(n_216),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_290),
.Y(n_427)
);

BUFx12f_ASAP7_75t_L g428 ( 
.A(n_299),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_319),
.A2(n_145),
.B(n_158),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_289),
.A2(n_169),
.B(n_133),
.Y(n_430)
);

AND3x2_ASAP7_75t_L g431 ( 
.A(n_325),
.B(n_221),
.C(n_175),
.Y(n_431)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_290),
.A2(n_175),
.B(n_133),
.Y(n_432)
);

OA21x2_ASAP7_75t_L g433 ( 
.A1(n_289),
.A2(n_169),
.B(n_167),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g434 ( 
.A1(n_315),
.A2(n_167),
.B(n_156),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_274),
.Y(n_435)
);

AO22x2_ASAP7_75t_L g436 ( 
.A1(n_341),
.A2(n_156),
.B1(n_167),
.B2(n_160),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_315),
.A2(n_167),
.B(n_146),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_315),
.A2(n_146),
.B(n_145),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_313),
.B(n_160),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_291),
.B(n_146),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_319),
.A2(n_158),
.B(n_145),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_316),
.A2(n_146),
.B(n_160),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_316),
.A2(n_146),
.B(n_160),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_348),
.A2(n_158),
.B(n_145),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_291),
.Y(n_445)
);

AO31x2_ASAP7_75t_L g446 ( 
.A1(n_341),
.A2(n_158),
.A3(n_145),
.B(n_160),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_285),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_292),
.B(n_146),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_356),
.A2(n_344),
.B(n_287),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_394),
.A2(n_358),
.B(n_425),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_377),
.A2(n_335),
.B1(n_285),
.B2(n_282),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_377),
.A2(n_285),
.B1(n_325),
.B2(n_344),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

AO21x2_ASAP7_75t_L g456 ( 
.A1(n_367),
.A2(n_300),
.B(n_303),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_353),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_370),
.A2(n_335),
.B(n_348),
.C(n_344),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_371),
.A2(n_348),
.B(n_334),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_344),
.B(n_287),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_L g461 ( 
.A1(n_389),
.A2(n_368),
.B1(n_362),
.B2(n_420),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_396),
.A2(n_317),
.B(n_316),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_396),
.A2(n_317),
.B(n_327),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_352),
.B(n_281),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_355),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_373),
.B(n_306),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_408),
.B(n_401),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_355),
.Y(n_471)
);

O2A1O1Ixp33_ASAP7_75t_SL g472 ( 
.A1(n_388),
.A2(n_328),
.B(n_296),
.C(n_334),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_363),
.A2(n_285),
.B1(n_344),
.B2(n_311),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

OA21x2_ASAP7_75t_L g475 ( 
.A1(n_357),
.A2(n_300),
.B(n_292),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_355),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_373),
.B(n_397),
.Y(n_477)
);

OAI211xp5_ASAP7_75t_L g478 ( 
.A1(n_389),
.A2(n_336),
.B(n_293),
.C(n_309),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_427),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_363),
.A2(n_285),
.B1(n_311),
.B2(n_295),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_387),
.A2(n_296),
.B(n_349),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g482 ( 
.A1(n_357),
.A2(n_309),
.B(n_293),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_373),
.B(n_311),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_427),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_387),
.A2(n_349),
.B(n_303),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_437),
.A2(n_336),
.B(n_341),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_372),
.A2(n_330),
.B(n_327),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_386),
.A2(n_327),
.B(n_317),
.Y(n_492)
);

OAI221xp5_ASAP7_75t_L g493 ( 
.A1(n_378),
.A2(n_339),
.B1(n_294),
.B2(n_298),
.C(n_333),
.Y(n_493)
);

AOI221x1_ASAP7_75t_L g494 ( 
.A1(n_363),
.A2(n_329),
.B1(n_330),
.B2(n_349),
.C(n_333),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_375),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_386),
.A2(n_330),
.B(n_329),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_369),
.A2(n_402),
.B(n_426),
.C(n_409),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_375),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_388),
.B(n_391),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_363),
.A2(n_311),
.B1(n_295),
.B2(n_313),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_395),
.A2(n_329),
.B(n_283),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_367),
.A2(n_279),
.B(n_294),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_379),
.B(n_311),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g506 ( 
.A1(n_413),
.A2(n_274),
.B1(n_295),
.B2(n_281),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_435),
.Y(n_507)
);

AOI221xp5_ASAP7_75t_L g508 ( 
.A1(n_380),
.A2(n_349),
.B1(n_339),
.B2(n_294),
.C(n_333),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_432),
.A2(n_279),
.B(n_333),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_375),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_432),
.A2(n_279),
.B(n_298),
.Y(n_511)
);

AOI21x1_ASAP7_75t_L g512 ( 
.A1(n_436),
.A2(n_349),
.B(n_283),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_393),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_393),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

AOI21xp33_ASAP7_75t_L g516 ( 
.A1(n_380),
.A2(n_311),
.B(n_298),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_360),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_436),
.A2(n_283),
.B(n_160),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_391),
.B(n_412),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_361),
.B(n_281),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_405),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_407),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_397),
.B(n_345),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_412),
.B(n_298),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_442),
.A2(n_443),
.B(n_437),
.Y(n_526)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_428),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_398),
.A2(n_274),
.B1(n_294),
.B2(n_273),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_406),
.B(n_279),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_442),
.A2(n_160),
.B(n_172),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_379),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_381),
.B(n_132),
.C(n_161),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_376),
.B(n_281),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_381),
.A2(n_145),
.B(n_158),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_411),
.Y(n_538)
);

O2A1O1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_382),
.A2(n_345),
.B(n_172),
.C(n_0),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_443),
.A2(n_160),
.B(n_172),
.Y(n_540)
);

AO21x2_ASAP7_75t_L g541 ( 
.A1(n_404),
.A2(n_172),
.B(n_141),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_406),
.B(n_273),
.Y(n_542)
);

AO21x2_ASAP7_75t_L g543 ( 
.A1(n_404),
.A2(n_141),
.B(n_132),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_428),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_399),
.A2(n_320),
.B(n_141),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_440),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_406),
.B(n_345),
.Y(n_547)
);

AO21x2_ASAP7_75t_L g548 ( 
.A1(n_382),
.A2(n_141),
.B(n_132),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_383),
.A2(n_158),
.B(n_281),
.Y(n_549)
);

O2A1O1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_398),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_399),
.A2(n_416),
.B(n_410),
.Y(n_551)
);

AOI22x1_ASAP7_75t_L g552 ( 
.A1(n_429),
.A2(n_183),
.B1(n_161),
.B2(n_132),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_534),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_452),
.A2(n_406),
.B1(n_392),
.B2(n_447),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_468),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_447),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_468),
.Y(n_557)
);

AO22x1_ASAP7_75t_SL g558 ( 
.A1(n_527),
.A2(n_428),
.B1(n_397),
.B2(n_439),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g559 ( 
.A1(n_451),
.A2(n_365),
.B(n_424),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_469),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_528),
.A2(n_423),
.B1(n_435),
.B2(n_281),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_534),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_519),
.B(n_352),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_471),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_471),
.Y(n_567)
);

CKINVDCx11_ASAP7_75t_R g568 ( 
.A(n_527),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_475),
.Y(n_570)
);

OAI221xp5_ASAP7_75t_L g571 ( 
.A1(n_452),
.A2(n_414),
.B1(n_418),
.B2(n_448),
.C(n_403),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_528),
.A2(n_435),
.B1(n_397),
.B2(n_421),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_461),
.A2(n_431),
.B1(n_436),
.B2(n_365),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_470),
.A2(n_493),
.B1(n_501),
.B2(n_458),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_455),
.Y(n_575)
);

OAI211xp5_ASAP7_75t_L g576 ( 
.A1(n_550),
.A2(n_478),
.B(n_539),
.C(n_499),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_466),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_517),
.A2(n_436),
.B1(n_365),
.B2(n_364),
.Y(n_578)
);

AOI211xp5_ASAP7_75t_L g579 ( 
.A1(n_501),
.A2(n_516),
.B(n_463),
.C(n_479),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_454),
.A2(n_385),
.B1(n_439),
.B2(n_354),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_477),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_494),
.A2(n_405),
.B1(n_352),
.B2(n_364),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_476),
.Y(n_584)
);

AOI21xp33_ASAP7_75t_L g585 ( 
.A1(n_546),
.A2(n_364),
.B(n_433),
.Y(n_585)
);

AOI222xp33_ASAP7_75t_L g586 ( 
.A1(n_473),
.A2(n_430),
.B1(n_439),
.B2(n_438),
.C1(n_384),
.C2(n_383),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_SL g587 ( 
.A(n_544),
.B(n_444),
.C(n_441),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_527),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_497),
.B(n_439),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_525),
.B(n_430),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_455),
.B(n_359),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_525),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_450),
.B(n_433),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_475),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_475),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_455),
.B(n_359),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_433),
.Y(n_597)
);

AO31x2_ASAP7_75t_L g598 ( 
.A1(n_494),
.A2(n_446),
.A3(n_366),
.B(n_433),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_457),
.B(n_421),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_469),
.Y(n_600)
);

CKINVDCx6p67_ASAP7_75t_R g601 ( 
.A(n_490),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_476),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_490),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_482),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_490),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_542),
.A2(n_354),
.B1(n_438),
.B2(n_359),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_536),
.A2(n_485),
.B1(n_505),
.B2(n_481),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_485),
.A2(n_359),
.B1(n_421),
.B2(n_320),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_491),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_482),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_508),
.A2(n_421),
.B1(n_320),
.B2(n_141),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_502),
.A2(n_384),
.B1(n_320),
.B2(n_416),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_482),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_491),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_477),
.B(n_524),
.Y(n_615)
);

NAND2x1_ASAP7_75t_L g616 ( 
.A(n_453),
.B(n_141),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_457),
.B(n_1),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_530),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_469),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_491),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_505),
.A2(n_481),
.B1(n_546),
.B2(n_474),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_480),
.A2(n_320),
.B1(n_410),
.B2(n_132),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_463),
.B(n_446),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_477),
.B(n_446),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_482),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_500),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_477),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_520),
.A2(n_320),
.B1(n_132),
.B2(n_183),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_547),
.A2(n_320),
.B1(n_161),
.B2(n_183),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_552),
.A2(n_434),
.B(n_422),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_500),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_474),
.B(n_2),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_479),
.B(n_446),
.Y(n_634)
);

AO31x2_ASAP7_75t_L g635 ( 
.A1(n_488),
.A2(n_529),
.A3(n_500),
.B(n_496),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_484),
.B(n_4),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_469),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_483),
.B(n_547),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_552),
.A2(n_434),
.B(n_422),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_SL g640 ( 
.A1(n_459),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_460),
.A2(n_419),
.B1(n_446),
.B2(n_183),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_483),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_460),
.A2(n_419),
.B1(n_446),
.B2(n_183),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_568),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_563),
.B(n_484),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_576),
.A2(n_507),
.B1(n_453),
.B2(n_535),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_593),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_565),
.B(n_487),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_561),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_577),
.B(n_487),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_574),
.A2(n_554),
.B1(n_573),
.B2(n_578),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_573),
.A2(n_483),
.B1(n_524),
.B2(n_516),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_565),
.B(n_489),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_606),
.A2(n_507),
.B1(n_453),
.B2(n_535),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_593),
.Y(n_655)
);

BUFx12f_ASAP7_75t_L g656 ( 
.A(n_614),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_562),
.A2(n_472),
.B(n_449),
.Y(n_657)
);

OA21x2_ASAP7_75t_L g658 ( 
.A1(n_631),
.A2(n_551),
.B(n_526),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_635),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_553),
.B(n_489),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_SL g661 ( 
.A1(n_581),
.A2(n_483),
.B1(n_524),
.B2(n_541),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_625),
.A2(n_524),
.B1(n_510),
.B2(n_531),
.Y(n_662)
);

BUFx12f_ASAP7_75t_L g663 ( 
.A(n_614),
.Y(n_663)
);

AOI21xp33_ASAP7_75t_SL g664 ( 
.A1(n_617),
.A2(n_6),
.B(n_8),
.Y(n_664)
);

AOI21xp33_ASAP7_75t_SL g665 ( 
.A1(n_633),
.A2(n_9),
.B(n_11),
.Y(n_665)
);

AOI21xp33_ASAP7_75t_L g666 ( 
.A1(n_579),
.A2(n_513),
.B(n_510),
.Y(n_666)
);

NAND2x1_ASAP7_75t_L g667 ( 
.A(n_591),
.B(n_507),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_621),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_555),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_625),
.A2(n_513),
.B1(n_496),
.B2(n_514),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_635),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_625),
.A2(n_514),
.B1(n_531),
.B2(n_523),
.Y(n_672)
);

OAI221xp5_ASAP7_75t_L g673 ( 
.A1(n_640),
.A2(n_449),
.B1(n_521),
.B2(n_495),
.C(n_503),
.Y(n_673)
);

OAI221xp5_ASAP7_75t_L g674 ( 
.A1(n_636),
.A2(n_521),
.B1(n_495),
.B2(n_538),
.C(n_533),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_556),
.A2(n_515),
.B1(n_522),
.B2(n_533),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_572),
.A2(n_506),
.B(n_456),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_635),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_561),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_556),
.B(n_515),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_605),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_555),
.Y(n_681)
);

AOI221xp5_ASAP7_75t_L g682 ( 
.A1(n_622),
.A2(n_523),
.B1(n_522),
.B2(n_538),
.C(n_456),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_606),
.A2(n_507),
.B1(n_453),
.B2(n_495),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_588),
.A2(n_537),
.B1(n_512),
.B2(n_549),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_605),
.B(n_512),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_635),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_588),
.A2(n_537),
.B1(n_549),
.B2(n_467),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_SL g688 ( 
.A1(n_581),
.A2(n_541),
.B1(n_456),
.B2(n_548),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_557),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_635),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_624),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_624),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_589),
.A2(n_529),
.B1(n_456),
.B2(n_541),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_621),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_592),
.A2(n_634),
.B1(n_571),
.B2(n_628),
.Y(n_695)
);

OAI211xp5_ASAP7_75t_L g696 ( 
.A1(n_553),
.A2(n_486),
.B(n_504),
.C(n_518),
.Y(n_696)
);

OAI33xp33_ASAP7_75t_L g697 ( 
.A1(n_607),
.A2(n_9),
.A3(n_12),
.B1(n_13),
.B2(n_16),
.B3(n_18),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_634),
.A2(n_529),
.B1(n_541),
.B2(n_548),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_L g699 ( 
.A1(n_580),
.A2(n_518),
.B1(n_467),
.B2(n_486),
.Y(n_699)
);

OAI211xp5_ASAP7_75t_L g700 ( 
.A1(n_564),
.A2(n_486),
.B(n_504),
.C(n_509),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_564),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_597),
.B(n_548),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_601),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_581),
.A2(n_548),
.B1(n_543),
.B2(n_486),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_557),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_560),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_601),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_638),
.A2(n_543),
.B1(n_492),
.B2(n_498),
.Y(n_708)
);

OAI211xp5_ASAP7_75t_L g709 ( 
.A1(n_599),
.A2(n_511),
.B(n_509),
.C(n_465),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_608),
.A2(n_467),
.B1(n_183),
.B2(n_161),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_560),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_580),
.A2(n_183),
.B1(n_161),
.B2(n_162),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_638),
.B(n_543),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_638),
.A2(n_543),
.B1(n_498),
.B2(n_492),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_603),
.B(n_465),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_603),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_600),
.A2(n_462),
.B1(n_511),
.B2(n_545),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_566),
.Y(n_718)
);

AOI21x1_ASAP7_75t_L g719 ( 
.A1(n_639),
.A2(n_551),
.B(n_526),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_609),
.B(n_462),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_566),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_569),
.A2(n_545),
.A3(n_540),
.B(n_532),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_R g723 ( 
.A1(n_591),
.A2(n_12),
.B(n_19),
.Y(n_723)
);

OAI211xp5_ASAP7_75t_L g724 ( 
.A1(n_609),
.A2(n_20),
.B(n_22),
.C(n_24),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_600),
.A2(n_183),
.B1(n_161),
.B2(n_540),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_558),
.Y(n_726)
);

AOI222xp33_ASAP7_75t_L g727 ( 
.A1(n_590),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.C1(n_28),
.C2(n_29),
.Y(n_727)
);

AOI222xp33_ASAP7_75t_L g728 ( 
.A1(n_582),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.C1(n_36),
.C2(n_37),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_647),
.B(n_595),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_647),
.B(n_595),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_685),
.B(n_594),
.Y(n_731)
);

AND2x4_ASAP7_75t_SL g732 ( 
.A(n_713),
.B(n_642),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_659),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_655),
.B(n_594),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_685),
.B(n_569),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_655),
.B(n_570),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_691),
.B(n_604),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_691),
.B(n_604),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_692),
.B(n_610),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_716),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_692),
.B(n_610),
.Y(n_741)
);

INVxp67_ASAP7_75t_R g742 ( 
.A(n_684),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_680),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_713),
.B(n_570),
.Y(n_744)
);

AO21x2_ASAP7_75t_L g745 ( 
.A1(n_676),
.A2(n_613),
.B(n_626),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_659),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_671),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_648),
.B(n_613),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_671),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_685),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_677),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_648),
.B(n_626),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_715),
.B(n_559),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_653),
.B(n_559),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_701),
.Y(n_755)
);

OAI222xp33_ASAP7_75t_L g756 ( 
.A1(n_651),
.A2(n_612),
.B1(n_637),
.B2(n_561),
.C1(n_619),
.C2(n_575),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_677),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_686),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_686),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_690),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_653),
.B(n_559),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_658),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_660),
.B(n_598),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_716),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_690),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_660),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_705),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_705),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_715),
.B(n_642),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_711),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_720),
.B(n_598),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_718),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_718),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_721),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_721),
.B(n_600),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_702),
.B(n_598),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_723),
.A2(n_612),
.B1(n_581),
.B2(n_641),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_658),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_658),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_680),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_720),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_704),
.B(n_598),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_658),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_688),
.B(n_598),
.Y(n_785)
);

AND2x2_ASAP7_75t_SL g786 ( 
.A(n_682),
.B(n_619),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_719),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_702),
.B(n_575),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_669),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_719),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_698),
.B(n_708),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_657),
.B(n_643),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_645),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_679),
.B(n_619),
.Y(n_794)
);

OR2x6_ASAP7_75t_SL g795 ( 
.A(n_703),
.B(n_602),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_680),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_697),
.A2(n_587),
.B1(n_615),
.B2(n_611),
.C(n_596),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_650),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_668),
.B(n_618),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_668),
.B(n_694),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_791),
.A2(n_726),
.B1(n_728),
.B2(n_727),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_782),
.B(n_744),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_SL g803 ( 
.A1(n_791),
.A2(n_726),
.B1(n_724),
.B2(n_674),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_796),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_750),
.B(n_680),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_782),
.B(n_680),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_798),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_798),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_792),
.B(n_665),
.C(n_793),
.Y(n_809)
);

AOI222xp33_ASAP7_75t_L g810 ( 
.A1(n_791),
.A2(n_695),
.B1(n_652),
.B2(n_693),
.C1(n_699),
.C2(n_712),
.Y(n_810)
);

AOI221xp5_ASAP7_75t_L g811 ( 
.A1(n_785),
.A2(n_665),
.B1(n_664),
.B2(n_666),
.C(n_675),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_793),
.B(n_668),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_755),
.Y(n_813)
);

OAI33xp33_ASAP7_75t_L g814 ( 
.A1(n_766),
.A2(n_646),
.A3(n_687),
.B1(n_644),
.B2(n_703),
.B3(n_707),
.Y(n_814)
);

OAI211xp5_ASAP7_75t_L g815 ( 
.A1(n_792),
.A2(n_694),
.B(n_707),
.C(n_700),
.Y(n_815)
);

NOR2x1_ASAP7_75t_L g816 ( 
.A(n_799),
.B(n_694),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_750),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_771),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_771),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_791),
.A2(n_661),
.B1(n_662),
.B2(n_670),
.Y(n_820)
);

AOI33xp33_ASAP7_75t_L g821 ( 
.A1(n_772),
.A2(n_33),
.A3(n_34),
.B1(n_36),
.B2(n_37),
.B3(n_38),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_771),
.Y(n_822)
);

AOI222xp33_ASAP7_75t_L g823 ( 
.A1(n_792),
.A2(n_672),
.B1(n_710),
.B2(n_673),
.C1(n_681),
.C2(n_706),
.Y(n_823)
);

OAI31xp33_ASAP7_75t_L g824 ( 
.A1(n_778),
.A2(n_696),
.A3(n_654),
.B(n_709),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_766),
.B(n_649),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_740),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_771),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_755),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_742),
.A2(n_656),
.B1(n_663),
.B2(n_644),
.Y(n_829)
);

OAI33xp33_ASAP7_75t_L g830 ( 
.A1(n_764),
.A2(n_683),
.A3(n_41),
.B1(n_39),
.B2(n_689),
.B3(n_706),
.Y(n_830)
);

OAI211xp5_ASAP7_75t_SL g831 ( 
.A1(n_764),
.A2(n_678),
.B(n_649),
.C(n_717),
.Y(n_831)
);

NOR4xp25_ASAP7_75t_SL g832 ( 
.A(n_796),
.B(n_663),
.C(n_656),
.D(n_585),
.Y(n_832)
);

OR2x6_ASAP7_75t_L g833 ( 
.A(n_750),
.B(n_778),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_740),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_796),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_740),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_754),
.B(n_689),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_754),
.B(n_649),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_742),
.A2(n_667),
.B(n_616),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_771),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_774),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_742),
.A2(n_637),
.B1(n_667),
.B2(n_678),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_R g843 ( 
.A(n_799),
.B(n_800),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_774),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_744),
.B(n_714),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_744),
.B(n_678),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_774),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_750),
.B(n_637),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_774),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_774),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_743),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_736),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_767),
.Y(n_853)
);

OAI211xp5_ASAP7_75t_SL g854 ( 
.A1(n_797),
.A2(n_586),
.B(n_41),
.C(n_630),
.Y(n_854)
);

OAI21xp33_ASAP7_75t_L g855 ( 
.A1(n_785),
.A2(n_623),
.B(n_629),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_795),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_775),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_767),
.Y(n_858)
);

NAND4xp25_ASAP7_75t_L g859 ( 
.A(n_800),
.B(n_596),
.C(n_591),
.D(n_725),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_767),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_744),
.B(n_722),
.Y(n_861)
);

OR2x2_ASAP7_75t_SL g862 ( 
.A(n_763),
.B(n_600),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_747),
.B(n_642),
.C(n_600),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_797),
.B(n_616),
.C(n_596),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_775),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_SL g866 ( 
.A1(n_785),
.A2(n_642),
.B1(n_618),
.B2(n_669),
.Y(n_866)
);

AO21x2_ASAP7_75t_L g867 ( 
.A1(n_787),
.A2(n_681),
.B(n_602),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_775),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_775),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_786),
.A2(n_532),
.B(n_642),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_785),
.A2(n_618),
.B1(n_632),
.B2(n_627),
.Y(n_871)
);

OAI33xp33_ASAP7_75t_L g872 ( 
.A1(n_763),
.A2(n_584),
.A3(n_632),
.B1(n_627),
.B2(n_567),
.B3(n_583),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_775),
.Y(n_873)
);

AOI221xp5_ASAP7_75t_L g874 ( 
.A1(n_783),
.A2(n_583),
.B1(n_620),
.B2(n_584),
.C(n_567),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_778),
.A2(n_620),
.B1(n_722),
.B2(n_183),
.Y(n_875)
);

NOR4xp25_ASAP7_75t_SL g876 ( 
.A(n_747),
.B(n_722),
.C(n_161),
.D(n_162),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_768),
.Y(n_877)
);

OAI211xp5_ASAP7_75t_L g878 ( 
.A1(n_797),
.A2(n_722),
.B(n_162),
.C(n_161),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_750),
.B(n_722),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_783),
.A2(n_161),
.B1(n_162),
.B2(n_786),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_783),
.A2(n_162),
.B1(n_786),
.B2(n_754),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_733),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_786),
.A2(n_162),
.B1(n_795),
.B2(n_794),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_772),
.B(n_162),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_794),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_783),
.A2(n_162),
.B1(n_786),
.B2(n_754),
.Y(n_886)
);

AOI221xp5_ASAP7_75t_L g887 ( 
.A1(n_772),
.A2(n_162),
.B1(n_761),
.B2(n_753),
.C(n_756),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_795),
.A2(n_162),
.B1(n_794),
.B2(n_763),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_802),
.B(n_772),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_867),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_808),
.B(n_761),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_861),
.B(n_761),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_861),
.B(n_761),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_829),
.B(n_794),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_802),
.B(n_731),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_846),
.B(n_731),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_852),
.B(n_748),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_856),
.B(n_748),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_856),
.B(n_748),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_853),
.Y(n_900)
);

OAI31xp33_ASAP7_75t_L g901 ( 
.A1(n_801),
.A2(n_756),
.A3(n_763),
.B(n_777),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_846),
.B(n_731),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_807),
.B(n_748),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_858),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_879),
.B(n_735),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_885),
.B(n_777),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_860),
.Y(n_907)
);

AND2x2_ASAP7_75t_SL g908 ( 
.A(n_821),
.B(n_795),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_839),
.B(n_848),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_877),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_879),
.B(n_735),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_867),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_879),
.B(n_735),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_813),
.B(n_752),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_809),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_879),
.B(n_735),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_867),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_819),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_834),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_836),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_828),
.B(n_777),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_819),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_817),
.B(n_735),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_817),
.B(n_735),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_817),
.B(n_735),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_818),
.B(n_752),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_838),
.B(n_777),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_882),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_882),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_822),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_826),
.B(n_788),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_833),
.B(n_753),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_803),
.A2(n_753),
.B1(n_776),
.B2(n_731),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_845),
.B(n_731),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_818),
.B(n_752),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_827),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_811),
.A2(n_749),
.B(n_753),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_827),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_804),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_841),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_845),
.B(n_731),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_806),
.B(n_731),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_806),
.B(n_752),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_804),
.B(n_770),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_SL g945 ( 
.A(n_814),
.B(n_760),
.C(n_747),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_841),
.B(n_849),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_822),
.B(n_753),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_849),
.B(n_745),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_840),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_837),
.B(n_788),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_857),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_837),
.B(n_788),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_857),
.B(n_745),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_843),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_840),
.B(n_753),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_844),
.B(n_753),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_844),
.B(n_847),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_847),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_869),
.B(n_745),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_850),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_851),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_850),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_833),
.B(n_805),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_825),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_865),
.B(n_739),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_865),
.B(n_739),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_868),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_862),
.B(n_788),
.Y(n_968)
);

AND2x4_ASAP7_75t_SL g969 ( 
.A(n_848),
.B(n_770),
.Y(n_969)
);

NOR2x1p5_ASAP7_75t_L g970 ( 
.A(n_859),
.B(n_736),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_812),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_869),
.B(n_745),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_868),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_833),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_873),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_804),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_892),
.B(n_833),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_900),
.Y(n_978)
);

INVx3_ASAP7_75t_R g979 ( 
.A(n_963),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_900),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_904),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_892),
.B(n_873),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_904),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_907),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_911),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_915),
.B(n_824),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_937),
.B(n_875),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_915),
.B(n_823),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_890),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_934),
.B(n_805),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_893),
.B(n_736),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_907),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_910),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_893),
.B(n_736),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_891),
.B(n_737),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_890),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_910),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_891),
.B(n_737),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_945),
.B(n_835),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_890),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_921),
.B(n_737),
.Y(n_1001)
);

NAND2x1_ASAP7_75t_SL g1002 ( 
.A(n_963),
.B(n_816),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_934),
.B(n_941),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_912),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_954),
.B(n_830),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_934),
.B(n_805),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_921),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_914),
.B(n_741),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_918),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_941),
.B(n_835),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_908),
.B(n_848),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_918),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_912),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_912),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_945),
.B(n_835),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_903),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_941),
.B(n_851),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_922),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_922),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_889),
.B(n_739),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_917),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_917),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_971),
.B(n_729),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_903),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_963),
.B(n_911),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_971),
.B(n_729),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_969),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_914),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_917),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_889),
.B(n_739),
.Y(n_1030)
);

NAND4xp25_ASAP7_75t_L g1031 ( 
.A(n_937),
.B(n_821),
.C(n_815),
.D(n_864),
.Y(n_1031)
);

INVxp67_ASAP7_75t_SL g1032 ( 
.A(n_970),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_963),
.B(n_863),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_919),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_894),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_901),
.A2(n_854),
.B(n_878),
.C(n_883),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_906),
.B(n_738),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_906),
.B(n_738),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_930),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_909),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_911),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_908),
.A2(n_810),
.B1(n_855),
.B2(n_820),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_889),
.B(n_741),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_954),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_964),
.B(n_729),
.Y(n_1045)
);

AND3x2_ASAP7_75t_L g1046 ( 
.A(n_901),
.B(n_887),
.C(n_884),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_970),
.B(n_927),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_895),
.B(n_741),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_969),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_928),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_908),
.A2(n_886),
.B(n_881),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_1007),
.B(n_927),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_986),
.B(n_831),
.C(n_974),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_989),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1007),
.B(n_897),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_988),
.B(n_920),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_1044),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_980),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_980),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_981),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1003),
.B(n_969),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1003),
.B(n_895),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1032),
.B(n_1027),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_981),
.Y(n_1064)
);

NAND4xp25_ASAP7_75t_L g1065 ( 
.A(n_1031),
.B(n_933),
.C(n_976),
.D(n_939),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1027),
.B(n_895),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_989),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_983),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1049),
.B(n_898),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1049),
.B(n_898),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_1028),
.B(n_897),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_996),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_983),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_996),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_1005),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_SL g1076 ( 
.A1(n_1011),
.A2(n_932),
.B1(n_909),
.B2(n_880),
.Y(n_1076)
);

NAND4xp75_ASAP7_75t_SL g1077 ( 
.A(n_1010),
.B(n_899),
.C(n_944),
.D(n_925),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1042),
.A2(n_974),
.B1(n_932),
.B2(n_888),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_987),
.A2(n_932),
.B1(n_911),
.B2(n_913),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_984),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_1025),
.B(n_905),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1011),
.B(n_899),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1000),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1035),
.B(n_965),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1011),
.B(n_896),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1034),
.B(n_965),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_1016),
.B(n_950),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_984),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_992),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1024),
.B(n_965),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_990),
.B(n_896),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_990),
.B(n_896),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_991),
.B(n_950),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_992),
.Y(n_1094)
);

AO22x1_ASAP7_75t_L g1095 ( 
.A1(n_999),
.A2(n_905),
.B1(n_913),
.B2(n_916),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1015),
.B(n_966),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_993),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_987),
.A2(n_932),
.B1(n_913),
.B2(n_916),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_978),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_1040),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_991),
.B(n_952),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1025),
.B(n_905),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_1040),
.Y(n_1103)
);

NAND2x1_ASAP7_75t_L g1104 ( 
.A(n_985),
.B(n_939),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1047),
.B(n_966),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1023),
.B(n_966),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_993),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1006),
.B(n_902),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1026),
.B(n_1020),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1020),
.B(n_947),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_SL g1111 ( 
.A1(n_1051),
.A2(n_931),
.B(n_968),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_994),
.B(n_1008),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_994),
.B(n_952),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1006),
.B(n_902),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1008),
.B(n_926),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1030),
.B(n_902),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1001),
.B(n_926),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_987),
.A2(n_932),
.B(n_959),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_1002),
.Y(n_1119)
);

AOI211xp5_ASAP7_75t_L g1120 ( 
.A1(n_1065),
.A2(n_1036),
.B(n_916),
.C(n_1033),
.Y(n_1120)
);

AOI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_1075),
.A2(n_987),
.B(n_1050),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_1057),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_SL g1123 ( 
.A1(n_1056),
.A2(n_931),
.B(n_977),
.C(n_1001),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1053),
.B(n_1030),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_1104),
.A2(n_977),
.B(n_985),
.C(n_1041),
.Y(n_1125)
);

AOI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_1119),
.A2(n_1111),
.B(n_1103),
.Y(n_1126)
);

NAND4xp25_ASAP7_75t_SL g1127 ( 
.A(n_1098),
.B(n_1010),
.C(n_1017),
.D(n_1043),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1099),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1079),
.A2(n_1076),
.B1(n_1118),
.B2(n_1078),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1064),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1111),
.A2(n_1033),
.B(n_932),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1064),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1095),
.A2(n_972),
.B1(n_948),
.B2(n_959),
.C(n_953),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1094),
.Y(n_1134)
);

NAND4xp75_ASAP7_75t_L g1135 ( 
.A(n_1063),
.B(n_1082),
.C(n_1085),
.D(n_1054),
.Y(n_1135)
);

OAI222xp33_ASAP7_75t_L g1136 ( 
.A1(n_1063),
.A2(n_1046),
.B1(n_968),
.B2(n_1033),
.C1(n_1041),
.C2(n_985),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1084),
.B(n_1043),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1094),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1058),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_1096),
.A2(n_1002),
.B(n_1041),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1061),
.B(n_1048),
.Y(n_1141)
);

AOI322xp5_ASAP7_75t_L g1142 ( 
.A1(n_1105),
.A2(n_972),
.A3(n_953),
.B1(n_948),
.B2(n_947),
.C1(n_955),
.C2(n_956),
.Y(n_1142)
);

OAI21xp33_ASAP7_75t_L g1143 ( 
.A1(n_1086),
.A2(n_997),
.B(n_1045),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1059),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1095),
.A2(n_871),
.B1(n_866),
.B2(n_1050),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1061),
.B(n_1048),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1100),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1060),
.Y(n_1148)
);

OA211x2_ASAP7_75t_L g1149 ( 
.A1(n_1104),
.A2(n_979),
.B(n_935),
.C(n_1025),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1068),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_1081),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1082),
.B(n_1017),
.Y(n_1152)
);

AOI221x1_ASAP7_75t_L g1153 ( 
.A1(n_1073),
.A2(n_997),
.B1(n_1039),
.B2(n_1009),
.C(n_1012),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1081),
.A2(n_976),
.B(n_1019),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1080),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1085),
.B(n_923),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1052),
.A2(n_947),
.B1(n_955),
.B2(n_956),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1088),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1054),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1089),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_SL g1161 ( 
.A1(n_1081),
.A2(n_909),
.B(n_842),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1097),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1052),
.A2(n_955),
.B1(n_956),
.B2(n_776),
.Y(n_1163)
);

AOI221xp5_ASAP7_75t_L g1164 ( 
.A1(n_1107),
.A2(n_1039),
.B1(n_1009),
.B2(n_1018),
.C(n_1012),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1102),
.B(n_923),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1055),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1055),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1069),
.B(n_832),
.C(n_909),
.Y(n_1168)
);

INVxp67_ASAP7_75t_SL g1169 ( 
.A(n_1067),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1102),
.A2(n_776),
.B1(n_872),
.B2(n_1018),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1102),
.B(n_1019),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_1122),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1151),
.B(n_1093),
.Y(n_1173)
);

OAI21xp33_ASAP7_75t_SL g1174 ( 
.A1(n_1135),
.A2(n_1077),
.B(n_1062),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1120),
.B(n_1069),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1147),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1130),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1136),
.A2(n_1070),
.B(n_1090),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1132),
.Y(n_1179)
);

OAI221xp5_ASAP7_75t_SL g1180 ( 
.A1(n_1124),
.A2(n_1112),
.B1(n_1093),
.B2(n_1113),
.C(n_1101),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1166),
.B(n_1070),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_1121),
.A2(n_1071),
.B(n_1112),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1152),
.B(n_1091),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1151),
.B(n_1101),
.Y(n_1184)
);

AOI322xp5_ASAP7_75t_L g1185 ( 
.A1(n_1169),
.A2(n_1109),
.A3(n_1067),
.B1(n_1072),
.B2(n_1074),
.C1(n_1083),
.C2(n_1106),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1167),
.B(n_1116),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1129),
.A2(n_1072),
.B1(n_1074),
.B2(n_1083),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1134),
.Y(n_1188)
);

O2A1O1Ixp5_ASAP7_75t_L g1189 ( 
.A1(n_1126),
.A2(n_1066),
.B(n_1071),
.C(n_1062),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1123),
.A2(n_1087),
.B(n_1113),
.C(n_1110),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1149),
.A2(n_1161),
.B1(n_1145),
.B2(n_1131),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1152),
.Y(n_1192)
);

O2A1O1Ixp5_ASAP7_75t_SL g1193 ( 
.A1(n_1138),
.A2(n_930),
.B(n_975),
.C(n_949),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1123),
.A2(n_1087),
.B(n_1066),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1139),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1157),
.A2(n_1091),
.B1(n_1092),
.B2(n_1114),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1153),
.A2(n_1114),
.B(n_1108),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1128),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1144),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1148),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_SL g1201 ( 
.A(n_1140),
.B(n_961),
.Y(n_1201)
);

OAI21xp33_ASAP7_75t_L g1202 ( 
.A1(n_1127),
.A2(n_1115),
.B(n_1117),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1150),
.Y(n_1203)
);

AO22x2_ASAP7_75t_L g1204 ( 
.A1(n_1169),
.A2(n_1029),
.B1(n_1000),
.B2(n_1004),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1171),
.B(n_1116),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1170),
.A2(n_1168),
.B1(n_1159),
.B2(n_1171),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1155),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1158),
.Y(n_1208)
);

AOI322xp5_ASAP7_75t_L g1209 ( 
.A1(n_1133),
.A2(n_1021),
.A3(n_1013),
.B1(n_1014),
.B2(n_1029),
.C1(n_1022),
.C2(n_1004),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_L g1210 ( 
.A1(n_1160),
.A2(n_1108),
.B(n_1092),
.C(n_1022),
.Y(n_1210)
);

AOI21xp33_ASAP7_75t_L g1211 ( 
.A1(n_1162),
.A2(n_1021),
.B(n_1014),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1159),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1154),
.A2(n_1115),
.B(n_1117),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1171),
.B(n_961),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1137),
.B(n_979),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1141),
.Y(n_1216)
);

OAI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1163),
.A2(n_1038),
.B1(n_1037),
.B2(n_982),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1143),
.A2(n_982),
.B(n_961),
.Y(n_1218)
);

XNOR2xp5_ASAP7_75t_L g1219 ( 
.A(n_1172),
.B(n_1187),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1172),
.A2(n_1164),
.B(n_1165),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_SL g1221 ( 
.A(n_1180),
.B(n_1125),
.C(n_1165),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1176),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1212),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1177),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1183),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_SL g1226 ( 
.A(n_1192),
.B(n_1141),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1173),
.B(n_1146),
.Y(n_1227)
);

XNOR2x1_ASAP7_75t_L g1228 ( 
.A(n_1191),
.B(n_1204),
.Y(n_1228)
);

AOI322xp5_ASAP7_75t_L g1229 ( 
.A1(n_1175),
.A2(n_1142),
.A3(n_1156),
.B1(n_1146),
.B2(n_1013),
.C1(n_874),
.C2(n_1125),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1189),
.B(n_1156),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1179),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1189),
.B(n_923),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_SL g1233 ( 
.A(n_1180),
.B(n_958),
.C(n_949),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1185),
.B(n_762),
.C(n_884),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1188),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1195),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1204),
.Y(n_1237)
);

XNOR2x1_ASAP7_75t_L g1238 ( 
.A(n_1204),
.B(n_1038),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1198),
.B(n_1037),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1186),
.B(n_998),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1216),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1210),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1181),
.B(n_998),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1200),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1203),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1207),
.Y(n_1246)
);

NAND2xp33_ASAP7_75t_SL g1247 ( 
.A(n_1208),
.B(n_995),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1184),
.B(n_942),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_R g1249 ( 
.A(n_1194),
.B(n_876),
.Y(n_1249)
);

NOR2x1_ASAP7_75t_L g1250 ( 
.A(n_1214),
.B(n_923),
.Y(n_1250)
);

XNOR2x1_ASAP7_75t_L g1251 ( 
.A(n_1206),
.B(n_995),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1199),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1205),
.B(n_935),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1182),
.B(n_943),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1199),
.B(n_943),
.Y(n_1255)
);

BUFx5_ASAP7_75t_L g1256 ( 
.A(n_1193),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1190),
.A2(n_946),
.B(n_940),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1215),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1210),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1174),
.B(n_762),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1178),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1196),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1202),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1220),
.A2(n_1228),
.B(n_1219),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1222),
.B(n_1213),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1261),
.A2(n_1211),
.B(n_1201),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1256),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_1225),
.B(n_1197),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1261),
.A2(n_1218),
.B1(n_1217),
.B2(n_1209),
.Y(n_1269)
);

OA22x2_ASAP7_75t_L g1270 ( 
.A1(n_1263),
.A2(n_924),
.B1(n_925),
.B2(n_944),
.Y(n_1270)
);

NOR3xp33_ASAP7_75t_L g1271 ( 
.A(n_1258),
.B(n_1252),
.C(n_1230),
.Y(n_1271)
);

NOR3xp33_ASAP7_75t_L g1272 ( 
.A(n_1230),
.B(n_946),
.C(n_928),
.Y(n_1272)
);

AOI211xp5_ASAP7_75t_L g1273 ( 
.A1(n_1242),
.A2(n_762),
.B(n_784),
.C(n_779),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1242),
.A2(n_762),
.B1(n_784),
.B2(n_779),
.C(n_780),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1237),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1221),
.B(n_1226),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1221),
.B(n_1256),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1239),
.B(n_943),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1233),
.A2(n_925),
.B(n_924),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_1241),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1239),
.B(n_957),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1259),
.A2(n_779),
.B(n_784),
.C(n_780),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1233),
.A2(n_924),
.B(n_957),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1248),
.B(n_942),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1229),
.A2(n_957),
.B(n_973),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1256),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1236),
.B(n_973),
.Y(n_1287)
);

NOR2x1_ASAP7_75t_L g1288 ( 
.A(n_1236),
.B(n_973),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1241),
.B(n_1227),
.Y(n_1289)
);

AOI211xp5_ASAP7_75t_L g1290 ( 
.A1(n_1260),
.A2(n_762),
.B(n_779),
.C(n_780),
.Y(n_1290)
);

AND2x2_ASAP7_75t_SL g1291 ( 
.A(n_1244),
.B(n_762),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1262),
.B(n_942),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1223),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1245),
.B(n_975),
.Y(n_1294)
);

NOR4xp25_ASAP7_75t_L g1295 ( 
.A(n_1246),
.B(n_967),
.C(n_962),
.D(n_960),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1250),
.B(n_967),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1280),
.B(n_1231),
.Y(n_1297)
);

OAI222xp33_ASAP7_75t_L g1298 ( 
.A1(n_1277),
.A2(n_1264),
.B1(n_1269),
.B2(n_1266),
.C1(n_1276),
.C2(n_1260),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1289),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_SL g1300 ( 
.A(n_1277),
.B(n_1224),
.C(n_1235),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1268),
.A2(n_1238),
.B1(n_1256),
.B2(n_1251),
.Y(n_1301)
);

OAI32xp33_ASAP7_75t_L g1302 ( 
.A1(n_1276),
.A2(n_1249),
.A3(n_1247),
.B1(n_1232),
.B2(n_1234),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1267),
.A2(n_1247),
.B1(n_1257),
.B2(n_1232),
.C(n_1254),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1275),
.Y(n_1304)
);

OAI211xp5_ASAP7_75t_L g1305 ( 
.A1(n_1271),
.A2(n_1255),
.B(n_1256),
.C(n_1243),
.Y(n_1305)
);

NAND4xp25_ASAP7_75t_L g1306 ( 
.A(n_1265),
.B(n_1249),
.C(n_1240),
.D(n_1253),
.Y(n_1306)
);

NAND4xp25_ASAP7_75t_L g1307 ( 
.A(n_1267),
.B(n_1256),
.C(n_962),
.D(n_960),
.Y(n_1307)
);

O2A1O1Ixp5_ASAP7_75t_L g1308 ( 
.A1(n_1286),
.A2(n_958),
.B(n_951),
.C(n_940),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1272),
.A2(n_951),
.B1(n_940),
.B2(n_938),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_SL g1310 ( 
.A(n_1293),
.B(n_870),
.C(n_765),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1273),
.B(n_762),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1286),
.A2(n_951),
.B(n_938),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1288),
.A2(n_938),
.B(n_936),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1285),
.A2(n_779),
.B(n_784),
.C(n_780),
.Y(n_1314)
);

AOI321xp33_ASAP7_75t_L g1315 ( 
.A1(n_1290),
.A2(n_780),
.A3(n_784),
.B1(n_749),
.B2(n_760),
.C(n_757),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1292),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1278),
.A2(n_1270),
.B1(n_1281),
.B2(n_1292),
.Y(n_1317)
);

AOI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1295),
.A2(n_1274),
.B1(n_1282),
.B2(n_1287),
.C(n_1294),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1287),
.B(n_1284),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1270),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1283),
.A2(n_762),
.B1(n_929),
.B2(n_928),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1279),
.A2(n_745),
.B(n_929),
.C(n_936),
.Y(n_1322)
);

AOI221xp5_ASAP7_75t_L g1323 ( 
.A1(n_1296),
.A2(n_762),
.B1(n_745),
.B2(n_936),
.C(n_929),
.Y(n_1323)
);

AOI221xp5_ASAP7_75t_L g1324 ( 
.A1(n_1296),
.A2(n_762),
.B1(n_790),
.B2(n_787),
.C(n_765),
.Y(n_1324)
);

OAI211xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1291),
.A2(n_787),
.B(n_790),
.C(n_781),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1316),
.Y(n_1326)
);

NAND4xp25_ASAP7_75t_L g1327 ( 
.A(n_1301),
.B(n_1284),
.C(n_1291),
.D(n_790),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1299),
.B(n_738),
.Y(n_1328)
);

NOR3xp33_ASAP7_75t_L g1329 ( 
.A(n_1300),
.B(n_765),
.C(n_757),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1319),
.Y(n_1330)
);

AOI221x1_ASAP7_75t_L g1331 ( 
.A1(n_1300),
.A2(n_751),
.B1(n_760),
.B2(n_757),
.C(n_790),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1297),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1317),
.B(n_741),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1304),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1305),
.B(n_790),
.Y(n_1335)
);

OAI322xp33_ASAP7_75t_L g1336 ( 
.A1(n_1320),
.A2(n_787),
.A3(n_751),
.B1(n_768),
.B2(n_769),
.C1(n_773),
.C2(n_758),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1306),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1307),
.A2(n_776),
.B1(n_743),
.B2(n_781),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1303),
.B(n_787),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_R g1340 ( 
.A(n_1298),
.B(n_781),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1310),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1318),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1302),
.B(n_729),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1308),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_R g1345 ( 
.A(n_1321),
.B(n_743),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1312),
.Y(n_1346)
);

AOI221xp5_ASAP7_75t_L g1347 ( 
.A1(n_1314),
.A2(n_751),
.B1(n_773),
.B2(n_769),
.C(n_768),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1313),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1326),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1332),
.B(n_1325),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1344),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1348),
.B(n_1323),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_L g1353 ( 
.A(n_1337),
.B(n_1342),
.C(n_1327),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1330),
.B(n_1322),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1334),
.A2(n_1315),
.B1(n_1309),
.B2(n_1311),
.Y(n_1355)
);

NOR3xp33_ASAP7_75t_SL g1356 ( 
.A(n_1341),
.B(n_1339),
.C(n_1333),
.Y(n_1356)
);

NOR2x1_ASAP7_75t_L g1357 ( 
.A(n_1335),
.B(n_1324),
.Y(n_1357)
);

NOR2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1328),
.B(n_730),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1346),
.A2(n_1329),
.B1(n_1339),
.B2(n_1338),
.C(n_1343),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1340),
.B(n_730),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1331),
.B(n_781),
.C(n_743),
.Y(n_1361)
);

NAND4xp25_ASAP7_75t_L g1362 ( 
.A(n_1353),
.B(n_1340),
.C(n_1347),
.D(n_1336),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1351),
.B(n_1345),
.C(n_773),
.Y(n_1363)
);

NOR2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1349),
.B(n_1345),
.Y(n_1364)
);

OAI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1357),
.A2(n_1359),
.B1(n_1354),
.B2(n_1352),
.C(n_1355),
.Y(n_1365)
);

NAND4xp25_ASAP7_75t_L g1366 ( 
.A(n_1350),
.B(n_730),
.C(n_734),
.D(n_737),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1360),
.A2(n_776),
.B1(n_769),
.B2(n_733),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1356),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_SL g1369 ( 
.A(n_1361),
.B(n_758),
.C(n_759),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1358),
.B(n_758),
.Y(n_1370)
);

AND3x2_ASAP7_75t_L g1371 ( 
.A(n_1353),
.B(n_770),
.C(n_738),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1350),
.A2(n_730),
.B(n_734),
.Y(n_1372)
);

NOR3xp33_ASAP7_75t_L g1373 ( 
.A(n_1353),
.B(n_759),
.C(n_733),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1349),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1365),
.A2(n_734),
.B(n_770),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1374),
.B(n_734),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1363),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1368),
.Y(n_1378)
);

OAI211xp5_ASAP7_75t_L g1379 ( 
.A1(n_1362),
.A2(n_759),
.B(n_733),
.C(n_746),
.Y(n_1379)
);

NAND4xp25_ASAP7_75t_L g1380 ( 
.A(n_1373),
.B(n_770),
.C(n_733),
.D(n_746),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1371),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1364),
.Y(n_1382)
);

XOR2x2_ASAP7_75t_L g1383 ( 
.A(n_1369),
.B(n_862),
.Y(n_1383)
);

NOR3xp33_ASAP7_75t_L g1384 ( 
.A(n_1370),
.B(n_746),
.C(n_758),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1372),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1366),
.B(n_746),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1376),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1381),
.B(n_1367),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1381),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1385),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1379),
.A2(n_776),
.B1(n_770),
.B2(n_758),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1378),
.A2(n_776),
.B1(n_770),
.B2(n_759),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1382),
.A2(n_746),
.B(n_759),
.Y(n_1393)
);

OAI222xp33_ASAP7_75t_L g1394 ( 
.A1(n_1377),
.A2(n_732),
.B1(n_776),
.B2(n_789),
.C1(n_1375),
.C2(n_1386),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1380),
.B(n_789),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1390),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1389),
.A2(n_1383),
.B(n_1384),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1387),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1398),
.Y(n_1399)
);

XNOR2xp5_ASAP7_75t_L g1400 ( 
.A(n_1396),
.B(n_1388),
.Y(n_1400)
);

OA22x2_ASAP7_75t_L g1401 ( 
.A1(n_1399),
.A2(n_1397),
.B1(n_1392),
.B2(n_1391),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1401),
.B(n_1400),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1402),
.A2(n_1395),
.B1(n_1393),
.B2(n_1394),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_R g1404 ( 
.A1(n_1403),
.A2(n_1393),
.B1(n_776),
.B2(n_732),
.C(n_789),
.Y(n_1404)
);

AOI211xp5_ASAP7_75t_L g1405 ( 
.A1(n_1404),
.A2(n_732),
.B(n_776),
.C(n_1390),
.Y(n_1405)
);


endmodule