module fake_ibex_1774_n_4927 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4927);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4927;

wire n_4557;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_962;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_3208;
wire n_4569;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_2253;
wire n_4479;
wire n_3858;
wire n_4173;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_3060;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_3293;
wire n_2550;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_3951;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_4757;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_3119;
wire n_2590;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_1471;
wire n_3441;
wire n_4559;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_4851;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_1127;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_2422;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_2223;
wire n_3876;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_1607;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_3096;
wire n_2059;
wire n_1278;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_985;
wire n_4611;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_4895;
wire n_3354;
wire n_4069;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_2574;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_4686;
wire n_4682;
wire n_2914;
wire n_1833;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_4733;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_960;
wire n_4412;
wire n_4266;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_3857;
wire n_2357;
wire n_4354;
wire n_2937;
wire n_3728;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_4539;
wire n_1205;
wire n_2969;
wire n_3550;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_3502;
wire n_3935;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_4926;
wire n_4688;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_1930;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_3484;
wire n_2485;
wire n_4477;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_3726;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_4491;
wire n_4672;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_4433;
wire n_3030;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4393;
wire n_3777;
wire n_4553;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_3633;
wire n_1731;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_2829;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_965;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_3787;
wire n_3445;
wire n_2080;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_2142;
wire n_3703;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_998;
wire n_1729;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_4579;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_4636;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_2442;
wire n_1067;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_1662;
wire n_3443;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_1660;
wire n_4000;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_3712;
wire n_2143;
wire n_4637;
wire n_4021;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_3327;
wire n_1114;
wire n_3647;
wire n_3928;
wire n_3619;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_1885;
wire n_1989;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_1221;
wire n_3875;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_4565;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_4574;
wire n_4242;
wire n_4748;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_4562;
wire n_1584;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_3050;
wire n_2666;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_4196;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_3036;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_3332;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_3861;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_1640;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_4590;
wire n_4602;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_1743;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_4159;
wire n_4372;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_3819;
wire n_3334;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_4360;
wire n_3653;
wire n_4897;
wire n_963;
wire n_2139;
wire n_3693;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_3641;
wire n_4887;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_3722;
wire n_3802;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_4806;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_2859;
wire n_2564;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_2114;
wire n_1609;
wire n_3530;
wire n_1132;
wire n_4548;
wire n_1803;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_2660;
wire n_4604;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_3282;
wire n_1003;
wire n_2708;
wire n_2748;
wire n_2224;
wire n_2233;
wire n_2499;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_1553;
wire n_3542;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_1189;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_2852;
wire n_2132;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_3785;
wire n_3525;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_2481;
wire n_4409;
wire n_1264;
wire n_2808;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_4152;
wire n_1352;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4255;
wire n_2908;
wire n_4561;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_3328;
wire n_2763;
wire n_994;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_961;
wire n_3735;
wire n_2127;
wire n_3028;
wire n_3228;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_2086;
wire n_4832;
wire n_3666;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2108;
wire n_2535;
wire n_2945;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_3302;
wire n_1673;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_2894;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_2315;
wire n_3623;
wire n_2157;
wire n_3446;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_1105;
wire n_2898;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_4670;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_4053;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_1693;
wire n_2081;
wire n_2993;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_3989;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_967;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_3430;
wire n_1685;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_1398;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_4088;
wire n_2136;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_2202;
wire n_2262;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_1080;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4668;
wire n_2383;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_2230;
wire n_3033;
wire n_2151;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_1606;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_2826;
wire n_2112;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_4671;
wire n_1326;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_3618;
wire n_2727;
wire n_2719;
wire n_2213;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_3847;
wire n_2203;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_2646;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_4136;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1360;
wire n_2070;
wire n_4098;
wire n_3471;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_1452;
wire n_4570;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_2819;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4407;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_3680;
wire n_3624;
wire n_2467;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1566;
wire n_1464;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_1608;
wire n_3776;
wire n_1009;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_4427;
wire n_3505;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_2525;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4297;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4880;
wire n_3167;
wire n_2986;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4176;
wire n_4454;
wire n_964;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_3867;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_3588;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_2187;
wire n_2105;
wire n_2642;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_4048;
wire n_4084;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_2849;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_4860;
wire n_4438;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_2665;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_2581;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_3454;
wire n_4143;
wire n_4410;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_1433;
wire n_1907;
wire n_3994;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_4487;
wire n_1165;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_3042;
wire n_2561;
wire n_2491;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_4811;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_1419;
wire n_4738;
wire n_1193;
wire n_980;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_4086;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_966;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4468;
wire n_3421;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_1791;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_1164;
wire n_3749;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

INVx1_ASAP7_75t_L g960 ( 
.A(n_263),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_616),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_120),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_225),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_936),
.Y(n_964)
);

BUFx10_ASAP7_75t_L g965 ( 
.A(n_835),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_608),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_81),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_141),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_572),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_770),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_929),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_488),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_403),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_628),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_742),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_406),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_416),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_483),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_204),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_657),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_195),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_670),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_438),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_239),
.Y(n_984)
);

BUFx10_ASAP7_75t_L g985 ( 
.A(n_418),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_441),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_240),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_643),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_908),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_9),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_508),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_258),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_176),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_512),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_331),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_944),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_311),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_120),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_838),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_895),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_837),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_877),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_57),
.Y(n_1003)
);

CKINVDCx11_ASAP7_75t_R g1004 ( 
.A(n_123),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_187),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_870),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_846),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_880),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_774),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_171),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_369),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_430),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_474),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_890),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_933),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_219),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_356),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_204),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_940),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_745),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_711),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_654),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_851),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_296),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_865),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_237),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_335),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_361),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_583),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_196),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_114),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_872),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_393),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_545),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_861),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_823),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_447),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_235),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_565),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_539),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_620),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_256),
.Y(n_1042)
);

CKINVDCx16_ASAP7_75t_R g1043 ( 
.A(n_923),
.Y(n_1043)
);

BUFx10_ASAP7_75t_L g1044 ( 
.A(n_174),
.Y(n_1044)
);

BUFx2_ASAP7_75t_SL g1045 ( 
.A(n_744),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_232),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_869),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_832),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_444),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_705),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_887),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_844),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_921),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_682),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_197),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_496),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_170),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_698),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_616),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_30),
.Y(n_1060)
);

CKINVDCx16_ASAP7_75t_R g1061 ( 
.A(n_769),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_7),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_377),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_333),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_832),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_435),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_199),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_163),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_64),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_887),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_103),
.Y(n_1071)
);

BUFx2_ASAP7_75t_SL g1072 ( 
.A(n_721),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_367),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_336),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_125),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_723),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_758),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_785),
.Y(n_1078)
);

BUFx10_ASAP7_75t_L g1079 ( 
.A(n_373),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_173),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_351),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_923),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_333),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_146),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_421),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_287),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_38),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_846),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_638),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_759),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_538),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_949),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_572),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_28),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_421),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_355),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_876),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_869),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_201),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_609),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_263),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_446),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_485),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_918),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_713),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_392),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_51),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_794),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_288),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_849),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_76),
.Y(n_1111)
);

BUFx10_ASAP7_75t_L g1112 ( 
.A(n_0),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_156),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_54),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_733),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_397),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_130),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_200),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_956),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_446),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_499),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_139),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_606),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_859),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_652),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_684),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_297),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_797),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_532),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_905),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_920),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_894),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_879),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_368),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_889),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_188),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_497),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_795),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_864),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_106),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_54),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_718),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_911),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_909),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_187),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_585),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_839),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_96),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_947),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_902),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_742),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_914),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_880),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_138),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_893),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_353),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_927),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_525),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_44),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_305),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_721),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_324),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_563),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_772),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_895),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_866),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_116),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_322),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_168),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_584),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_927),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_876),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_422),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_23),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_42),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_925),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_426),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_765),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_918),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_425),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_179),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_268),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_653),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_843),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_781),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_718),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_507),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_915),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_59),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_77),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_782),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_196),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_44),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_109),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_836),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_815),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_783),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_565),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_805),
.Y(n_1200)
);

INVxp67_ASAP7_75t_SL g1201 ( 
.A(n_874),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_948),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_744),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_441),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_924),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_194),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_575),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_755),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_672),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_853),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_378),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_350),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_798),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_930),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_641),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_230),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_680),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_372),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_885),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_469),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_950),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_472),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_655),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_561),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_953),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_183),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_189),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_862),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_272),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_219),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_408),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_450),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_406),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_324),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_490),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_379),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_888),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_948),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_922),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_764),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_756),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_951),
.Y(n_1242)
);

BUFx10_ASAP7_75t_L g1243 ( 
.A(n_325),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_165),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_645),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_595),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_556),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_522),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_750),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_586),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_337),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_407),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_468),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_384),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_669),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_215),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_113),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_812),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_501),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_867),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_902),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_899),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_64),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_36),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_829),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_322),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_847),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_857),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_870),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_953),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_882),
.Y(n_1271)
);

BUFx10_ASAP7_75t_L g1272 ( 
.A(n_196),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_829),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_167),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_105),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_844),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_866),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_249),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_435),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_66),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_864),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_652),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_632),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_640),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_200),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_500),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_236),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_440),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_738),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_654),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_868),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_266),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_528),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_934),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_213),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_98),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_747),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_268),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_23),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_873),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_178),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_935),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_932),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_952),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_131),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_856),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_261),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_438),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_804),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_105),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_43),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_428),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_850),
.Y(n_1313)
);

CKINVDCx16_ASAP7_75t_R g1314 ( 
.A(n_209),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_624),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_633),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_73),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_871),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_641),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_937),
.Y(n_1320)
);

BUFx10_ASAP7_75t_L g1321 ( 
.A(n_802),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_472),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_669),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_154),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_57),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_695),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_453),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_618),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_23),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_388),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_841),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_906),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_211),
.Y(n_1333)
);

CKINVDCx14_ASAP7_75t_R g1334 ( 
.A(n_926),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_238),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_833),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_612),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_858),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_775),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_949),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_381),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_317),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_272),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_606),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_592),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_578),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_288),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_121),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_786),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_87),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_47),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_514),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_931),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_589),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_874),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_422),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_838),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_570),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_938),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_214),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_3),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_661),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_498),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_729),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_324),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_900),
.Y(n_1366)
);

BUFx10_ASAP7_75t_L g1367 ( 
.A(n_916),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_597),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_919),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_847),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_681),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_531),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_281),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_647),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_845),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_405),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_852),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_955),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_868),
.Y(n_1379)
);

BUFx8_ASAP7_75t_SL g1380 ( 
.A(n_600),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_334),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_528),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_455),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_120),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_303),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_711),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_519),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_199),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_801),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_836),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_707),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_598),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_349),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_942),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_695),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_722),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_605),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_225),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_629),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_646),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_840),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_287),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_241),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_716),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_806),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_947),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_572),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_939),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_529),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_465),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_764),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_863),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_891),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_954),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_896),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_308),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_178),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_103),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_627),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_892),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_465),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_163),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_816),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_803),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_787),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_31),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_906),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_277),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_685),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_276),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_883),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_300),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_330),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_828),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_68),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_524),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_164),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_786),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_907),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_166),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_202),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_833),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_485),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_399),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_600),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_789),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_580),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_622),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_779),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_156),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_740),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_20),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_246),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_862),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_878),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_831),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_46),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_843),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_582),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_503),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_941),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_364),
.Y(n_1462)
);

CKINVDCx11_ASAP7_75t_R g1463 ( 
.A(n_901),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_903),
.Y(n_1464)
);

BUFx10_ASAP7_75t_L g1465 ( 
.A(n_431),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_523),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_693),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_848),
.Y(n_1468)
);

CKINVDCx16_ASAP7_75t_R g1469 ( 
.A(n_541),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_344),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_688),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_478),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_865),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_585),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_389),
.Y(n_1475)
);

CKINVDCx16_ASAP7_75t_R g1476 ( 
.A(n_301),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_877),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_93),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_855),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_913),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_553),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_246),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_261),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_215),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_119),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_24),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_298),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_946),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_912),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_945),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_296),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_144),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_886),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_141),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_381),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_494),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_958),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_760),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_278),
.Y(n_1499)
);

BUFx10_ASAP7_75t_L g1500 ( 
.A(n_101),
.Y(n_1500)
);

CKINVDCx16_ASAP7_75t_R g1501 ( 
.A(n_565),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_197),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_528),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_353),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_854),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_842),
.Y(n_1506)
);

BUFx10_ASAP7_75t_L g1507 ( 
.A(n_396),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_529),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_904),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_933),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_825),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_334),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_362),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_645),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_750),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_612),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_220),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_910),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_58),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_311),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_119),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_696),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_30),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_260),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_684),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_830),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_875),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_897),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_898),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_834),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_881),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_928),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_884),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_731),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_592),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_330),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_119),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_860),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_335),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_689),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_853),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_386),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_75),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_701),
.Y(n_1544)
);

BUFx5_ASAP7_75t_L g1545 ( 
.A(n_943),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_472),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_172),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_87),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_636),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_145),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_777),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_291),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_183),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_917),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_361),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1499),
.B(n_0),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1004),
.Y(n_1557)
);

INVxp33_ASAP7_75t_SL g1558 ( 
.A(n_1067),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1004),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1334),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1011),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1093),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_969),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1334),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1380),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1380),
.Y(n_1566)
);

CKINVDCx16_ASAP7_75t_R g1567 ( 
.A(n_1314),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1463),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1156),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1463),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1469),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1476),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1233),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1501),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1351),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1537),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1365),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_969),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_962),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_972),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1416),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_973),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1027),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1418),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1450),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1053),
.B(n_0),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1520),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_963),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1333),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_976),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1027),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_977),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1034),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1435),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_960),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_967),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_981),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_968),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_979),
.Y(n_1599)
);

CKINVDCx16_ASAP7_75t_R g1600 ( 
.A(n_963),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_984),
.Y(n_1601)
);

CKINVDCx16_ASAP7_75t_R g1602 ( 
.A(n_963),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_986),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1158),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_983),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_990),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_987),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1149),
.B(n_1),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1018),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1015),
.B(n_1),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_991),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1158),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_1193),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1028),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_992),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1039),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1429),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_993),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_994),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_L g1620 ( 
.A(n_1098),
.B(n_2),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_1193),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_995),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_997),
.Y(n_1623)
);

INVxp33_ASAP7_75t_SL g1624 ( 
.A(n_998),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1040),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1225),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1055),
.Y(n_1627)
);

INVxp33_ASAP7_75t_SL g1628 ( 
.A(n_1003),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_1253),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1060),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1005),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1010),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_SL g1633 ( 
.A(n_985),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1253),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1013),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1063),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1064),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1016),
.Y(n_1638)
);

CKINVDCx16_ASAP7_75t_R g1639 ( 
.A(n_985),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1545),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1017),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_1301),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1301),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1307),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1024),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_1292),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1026),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1030),
.Y(n_1648)
);

INVxp33_ASAP7_75t_SL g1649 ( 
.A(n_1031),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1033),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1066),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1083),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1268),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1101),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1107),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1128),
.B(n_2),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1037),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1038),
.Y(n_1658)
);

INVxp67_ASAP7_75t_SL g1659 ( 
.A(n_1012),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1042),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1046),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1049),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1116),
.Y(n_1663)
);

NOR2xp67_ASAP7_75t_L g1664 ( 
.A(n_1210),
.B(n_2),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1057),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1120),
.Y(n_1666)
);

XNOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1062),
.B(n_3),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1121),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1129),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1068),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1069),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1073),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1136),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1141),
.Y(n_1674)
);

CKINVDCx20_ASAP7_75t_R g1675 ( 
.A(n_1292),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1160),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1163),
.Y(n_1677)
);

CKINVDCx16_ASAP7_75t_R g1678 ( 
.A(n_985),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1177),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1307),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1461),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1192),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1075),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1273),
.B(n_3),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1231),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1084),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1659),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1640),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1561),
.Y(n_1689)
);

XOR2xp5_ASAP7_75t_L g1690 ( 
.A(n_1563),
.B(n_1322),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1558),
.B(n_1085),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1589),
.B(n_1306),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1593),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1562),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1593),
.Y(n_1695)
);

INVx6_ASAP7_75t_L g1696 ( 
.A(n_1588),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1569),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1573),
.Y(n_1698)
);

INVx4_ASAP7_75t_L g1699 ( 
.A(n_1633),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1600),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1575),
.B(n_1086),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1594),
.B(n_1459),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1577),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1581),
.B(n_1480),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1584),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1602),
.B(n_1044),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1585),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1639),
.B(n_1044),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1587),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1624),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1633),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1678),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1681),
.B(n_1044),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1593),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1628),
.B(n_1087),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1579),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1593),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1684),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1649),
.B(n_1213),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1595),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1626),
.B(n_1091),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1596),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1598),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1599),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1617),
.B(n_1079),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1605),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1607),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1609),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1614),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1616),
.B(n_1625),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1627),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1630),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1636),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1557),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1637),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1651),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1652),
.Y(n_1737)
);

OR2x6_ASAP7_75t_L g1738 ( 
.A(n_1653),
.B(n_1045),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1654),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1655),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1663),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1666),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1567),
.B(n_1079),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1668),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1580),
.B(n_1079),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_L g1746 ( 
.A(n_1669),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1673),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1674),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1582),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1676),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1677),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1679),
.B(n_1682),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1685),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1610),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1610),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1590),
.Y(n_1756)
);

INVx6_ASAP7_75t_L g1757 ( 
.A(n_1620),
.Y(n_1757)
);

BUFx8_ASAP7_75t_L g1758 ( 
.A(n_1559),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1656),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1656),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_L g1761 ( 
.A(n_1556),
.B(n_1061),
.C(n_1043),
.Y(n_1761)
);

AND2x6_ASAP7_75t_L g1762 ( 
.A(n_1556),
.B(n_1012),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1592),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1597),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1664),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1601),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1578),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1586),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1603),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1608),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1606),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1611),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1615),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1618),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1619),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1622),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1623),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1631),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1632),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1635),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1560),
.B(n_1094),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1638),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1571),
.B(n_1572),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1641),
.Y(n_1784)
);

AND3x2_ASAP7_75t_L g1785 ( 
.A(n_1568),
.B(n_1201),
.C(n_1332),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1645),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1647),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1648),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1686),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1650),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1657),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1658),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1660),
.Y(n_1793)
);

OA21x2_ASAP7_75t_L g1794 ( 
.A1(n_1661),
.A2(n_1071),
.B(n_978),
.Y(n_1794)
);

NAND2xp33_ASAP7_75t_L g1795 ( 
.A(n_1564),
.B(n_1545),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1662),
.Y(n_1796)
);

INVxp33_ASAP7_75t_L g1797 ( 
.A(n_1667),
.Y(n_1797)
);

AND3x2_ASAP7_75t_L g1798 ( 
.A(n_1570),
.B(n_1437),
.C(n_1071),
.Y(n_1798)
);

BUFx8_ASAP7_75t_L g1799 ( 
.A(n_1565),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1665),
.B(n_1112),
.Y(n_1800)
);

OA21x2_ASAP7_75t_L g1801 ( 
.A1(n_1670),
.A2(n_1080),
.B(n_978),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1671),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1672),
.B(n_1535),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1683),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1574),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1576),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1566),
.B(n_989),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1583),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1591),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1604),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1612),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1613),
.Y(n_1812)
);

INVx4_ASAP7_75t_L g1813 ( 
.A(n_1621),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1629),
.Y(n_1814)
);

INVxp33_ASAP7_75t_L g1815 ( 
.A(n_1634),
.Y(n_1815)
);

BUFx8_ASAP7_75t_L g1816 ( 
.A(n_1642),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1643),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1644),
.B(n_1112),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1646),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1675),
.B(n_1112),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1680),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1659),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1588),
.B(n_1243),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1593),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1659),
.B(n_1096),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1588),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1640),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1640),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1588),
.B(n_1243),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1589),
.B(n_989),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1640),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1659),
.Y(n_1832)
);

AND2x6_ASAP7_75t_L g1833 ( 
.A(n_1589),
.B(n_1056),
.Y(n_1833)
);

OA21x2_ASAP7_75t_L g1834 ( 
.A1(n_1640),
.A2(n_1081),
.B(n_1080),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1659),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1659),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1593),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1640),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1659),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1659),
.B(n_1099),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1640),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_SL g1842 ( 
.A1(n_1563),
.A2(n_1356),
.B1(n_1363),
.B2(n_1322),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1588),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1659),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1659),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1640),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1659),
.B(n_1102),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1659),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1588),
.B(n_1243),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1588),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1640),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1589),
.B(n_1164),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1588),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1588),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1558),
.A2(n_1363),
.B1(n_1387),
.B2(n_1356),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1659),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1640),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1659),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1659),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1588),
.B(n_1272),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1659),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1659),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1659),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1593),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1640),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1593),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1588),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1659),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1640),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1659),
.B(n_1106),
.Y(n_1870)
);

AND2x2_ASAP7_75t_R g1871 ( 
.A(n_1563),
.B(n_1387),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1659),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1633),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1659),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1659),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1588),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1659),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1659),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1659),
.B(n_1109),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1567),
.A2(n_1114),
.B1(n_1117),
.B2(n_1111),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1640),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1659),
.B(n_1118),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1633),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1640),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1640),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1659),
.B(n_1122),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1659),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1659),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1588),
.B(n_1272),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1588),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1593),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1659),
.B(n_1127),
.Y(n_1892)
);

INVx4_ASAP7_75t_L g1893 ( 
.A(n_1633),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1640),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1593),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1659),
.Y(n_1896)
);

OA21x2_ASAP7_75t_L g1897 ( 
.A1(n_1640),
.A2(n_1103),
.B(n_1081),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1659),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1567),
.A2(n_1137),
.B1(n_1140),
.B2(n_1134),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1659),
.B(n_1145),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1834),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1697),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1718),
.B(n_1726),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1754),
.A2(n_1056),
.B1(n_1266),
.B2(n_1074),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1700),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1706),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1698),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1736),
.B(n_1148),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1755),
.B(n_1154),
.Y(n_1909)
);

INVxp33_ASAP7_75t_SL g1910 ( 
.A(n_1712),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1707),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1834),
.Y(n_1912)
);

INVx4_ASAP7_75t_L g1913 ( 
.A(n_1696),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1745),
.B(n_1272),
.Y(n_1914)
);

INVx5_ASAP7_75t_L g1915 ( 
.A(n_1833),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1897),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1739),
.B(n_1159),
.Y(n_1917)
);

INVx2_ASAP7_75t_SL g1918 ( 
.A(n_1708),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1897),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1731),
.Y(n_1920)
);

INVx5_ASAP7_75t_L g1921 ( 
.A(n_1833),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1829),
.B(n_1164),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1710),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1725),
.B(n_1465),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1853),
.Y(n_1925)
);

AOI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1688),
.A2(n_1248),
.B(n_1235),
.Y(n_1926)
);

AND3x2_ASAP7_75t_L g1927 ( 
.A(n_1853),
.B(n_1502),
.C(n_1440),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1747),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1715),
.B(n_1465),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1759),
.B(n_1162),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1731),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1826),
.B(n_1095),
.Y(n_1932)
);

NOR2x1p5_ASAP7_75t_L g1933 ( 
.A(n_1843),
.B(n_1167),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1689),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1825),
.B(n_1168),
.Y(n_1935)
);

OAI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1855),
.A2(n_1502),
.B1(n_1519),
.B2(n_1440),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1849),
.B(n_1465),
.Y(n_1937)
);

AND2x6_ASAP7_75t_L g1938 ( 
.A(n_1889),
.B(n_1074),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1770),
.A2(n_1794),
.B1(n_1801),
.B2(n_1760),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1768),
.B(n_1500),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1794),
.A2(n_1266),
.B1(n_1296),
.B2(n_1280),
.Y(n_1941)
);

NAND2xp33_ASAP7_75t_L g1942 ( 
.A(n_1833),
.B(n_1545),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1801),
.A2(n_1324),
.B1(n_1325),
.B2(n_1308),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1694),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1744),
.Y(n_1945)
);

INVx5_ASAP7_75t_L g1946 ( 
.A(n_1744),
.Y(n_1946)
);

BUFx3_ASAP7_75t_L g1947 ( 
.A(n_1696),
.Y(n_1947)
);

AND3x2_ASAP7_75t_L g1948 ( 
.A(n_1867),
.B(n_1547),
.C(n_1519),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1781),
.B(n_1169),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1703),
.Y(n_1950)
);

CKINVDCx6p67_ASAP7_75t_R g1951 ( 
.A(n_1738),
.Y(n_1951)
);

BUFx3_ASAP7_75t_L g1952 ( 
.A(n_1867),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1699),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1850),
.B(n_1343),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1746),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1746),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_SL g1957 ( 
.A1(n_1716),
.A2(n_1552),
.B1(n_1547),
.B2(n_966),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1687),
.B(n_1173),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1771),
.B(n_1500),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1705),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1709),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1822),
.B(n_1174),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1840),
.B(n_1847),
.Y(n_1963)
);

OR2x6_ASAP7_75t_L g1964 ( 
.A(n_1890),
.B(n_1072),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1832),
.B(n_1175),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1890),
.Y(n_1966)
);

NOR2x1p5_ASAP7_75t_L g1967 ( 
.A(n_1711),
.B(n_1180),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1753),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1835),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1836),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1839),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1883),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1844),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1845),
.B(n_1182),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1893),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1704),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1722),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1848),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1856),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1858),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1704),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1727),
.Y(n_1982)
);

INVxp67_ASAP7_75t_SL g1983 ( 
.A(n_1854),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1713),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1859),
.Y(n_1985)
);

AND2x2_ASAP7_75t_SL g1986 ( 
.A(n_1876),
.B(n_1103),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1728),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1861),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1870),
.B(n_1187),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1716),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_L g1991 ( 
.A(n_1762),
.B(n_1720),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1879),
.B(n_1189),
.Y(n_1992)
);

BUFx10_ASAP7_75t_L g1993 ( 
.A(n_1734),
.Y(n_1993)
);

OAI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1738),
.A2(n_1552),
.B1(n_971),
.B2(n_996),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1729),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1764),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1862),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1732),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1882),
.B(n_1190),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1737),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1863),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1868),
.Y(n_2002)
);

INVx3_ASAP7_75t_L g2003 ( 
.A(n_1830),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1766),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_R g2005 ( 
.A(n_1779),
.B(n_1194),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1743),
.B(n_1500),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1740),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1751),
.Y(n_2008)
);

BUFx10_ASAP7_75t_L g2009 ( 
.A(n_1719),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1789),
.B(n_1507),
.Y(n_2010)
);

BUFx10_ASAP7_75t_L g2011 ( 
.A(n_1766),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1886),
.B(n_1198),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1723),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1724),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1802),
.B(n_1507),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1769),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1733),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1735),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1741),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1742),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1872),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1892),
.B(n_1900),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1874),
.Y(n_2023)
);

INVx6_ASAP7_75t_L g2024 ( 
.A(n_1769),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1875),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1804),
.B(n_1507),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1830),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1877),
.Y(n_2028)
);

INVx4_ASAP7_75t_L g2029 ( 
.A(n_1764),
.Y(n_2029)
);

AND2x2_ASAP7_75t_SL g2030 ( 
.A(n_1818),
.B(n_1113),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1878),
.B(n_1199),
.Y(n_2031)
);

AO22x2_ASAP7_75t_L g2032 ( 
.A1(n_1690),
.A2(n_1444),
.B1(n_1495),
.B2(n_1417),
.Y(n_2032)
);

BUFx3_ASAP7_75t_L g2033 ( 
.A(n_1758),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1765),
.B(n_1113),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1852),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1887),
.B(n_1204),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1748),
.Y(n_2037)
);

NAND2xp33_ASAP7_75t_L g2038 ( 
.A(n_1762),
.B(n_1545),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1750),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1691),
.B(n_965),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1888),
.B(n_1206),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1827),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_1820),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1852),
.B(n_1209),
.Y(n_2044)
);

AND2x6_ASAP7_75t_L g2045 ( 
.A(n_1763),
.B(n_1181),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_1756),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1828),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1831),
.Y(n_2048)
);

AND2x6_ASAP7_75t_L g2049 ( 
.A(n_1777),
.B(n_1181),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1896),
.B(n_1207),
.Y(n_2050)
);

INVx2_ASAP7_75t_SL g2051 ( 
.A(n_1757),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1838),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1841),
.Y(n_2053)
);

BUFx10_ASAP7_75t_L g2054 ( 
.A(n_1803),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1898),
.B(n_1211),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1692),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1762),
.A2(n_1761),
.B1(n_1702),
.B2(n_1692),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_1758),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1730),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1702),
.B(n_1212),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1780),
.Y(n_2061)
);

AND2x6_ASAP7_75t_L g2062 ( 
.A(n_1792),
.B(n_1793),
.Y(n_2062)
);

INVx2_ASAP7_75t_SL g2063 ( 
.A(n_1757),
.Y(n_2063)
);

INVx2_ASAP7_75t_SL g2064 ( 
.A(n_1803),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1752),
.B(n_1216),
.Y(n_2065)
);

AND3x2_ASAP7_75t_L g2066 ( 
.A(n_1873),
.B(n_971),
.C(n_966),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1846),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1851),
.Y(n_2068)
);

NOR2x1p5_ASAP7_75t_L g2069 ( 
.A(n_1783),
.B(n_1218),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1857),
.Y(n_2070)
);

AND2x6_ASAP7_75t_L g2071 ( 
.A(n_1772),
.B(n_1773),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1721),
.B(n_1701),
.Y(n_2072)
);

INVxp67_ASAP7_75t_L g2073 ( 
.A(n_1774),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1823),
.B(n_1220),
.Y(n_2074)
);

OR2x6_ASAP7_75t_L g2075 ( 
.A(n_1813),
.B(n_996),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_1690),
.Y(n_2076)
);

OR2x6_ASAP7_75t_L g2077 ( 
.A(n_1809),
.B(n_1000),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1775),
.A2(n_1350),
.B1(n_1352),
.B2(n_1327),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_1776),
.A2(n_1372),
.B1(n_1376),
.B2(n_1360),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1778),
.B(n_1222),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1865),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1798),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1782),
.B(n_1244),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_1860),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1816),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1869),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1881),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1800),
.B(n_1224),
.Y(n_2088)
);

AND2x6_ASAP7_75t_L g2089 ( 
.A(n_1784),
.B(n_1244),
.Y(n_2089)
);

AND2x6_ASAP7_75t_L g2090 ( 
.A(n_1786),
.B(n_1264),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_1767),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1884),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1885),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1807),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1787),
.B(n_1264),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1790),
.B(n_1226),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1749),
.B(n_965),
.Y(n_2097)
);

BUFx4f_ASAP7_75t_L g2098 ( 
.A(n_1809),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_1791),
.B(n_1227),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1894),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1796),
.B(n_1279),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1799),
.Y(n_2102)
);

INVx4_ASAP7_75t_L g2103 ( 
.A(n_1807),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1816),
.Y(n_2104)
);

NOR2x1p5_ASAP7_75t_L g2105 ( 
.A(n_1805),
.B(n_1229),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1795),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1693),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1880),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1806),
.B(n_1230),
.Y(n_2109)
);

AO21x2_ASAP7_75t_L g2110 ( 
.A1(n_1899),
.A2(n_1383),
.B(n_1381),
.Y(n_2110)
);

INVx4_ASAP7_75t_L g2111 ( 
.A(n_1785),
.Y(n_2111)
);

NAND2x1p5_ASAP7_75t_L g2112 ( 
.A(n_1808),
.B(n_1503),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1799),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1788),
.Y(n_2114)
);

XNOR2xp5_ASAP7_75t_L g2115 ( 
.A(n_1842),
.B(n_1000),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1797),
.B(n_965),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1812),
.B(n_1279),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1819),
.B(n_1388),
.Y(n_2118)
);

BUFx6f_ASAP7_75t_L g2119 ( 
.A(n_1693),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1695),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1695),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1714),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_1810),
.Y(n_2123)
);

NAND2xp33_ASAP7_75t_L g2124 ( 
.A(n_1714),
.B(n_1545),
.Y(n_2124)
);

AOI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_1811),
.A2(n_1385),
.B1(n_1453),
.B2(n_1428),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1717),
.Y(n_2126)
);

INVx4_ASAP7_75t_L g2127 ( 
.A(n_1717),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1824),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1824),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1814),
.B(n_1543),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1837),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1837),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_1817),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_1821),
.Y(n_2134)
);

INVx4_ASAP7_75t_L g2135 ( 
.A(n_1864),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1864),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1866),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1866),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1891),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1871),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1891),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1895),
.Y(n_2142)
);

BUFx2_ASAP7_75t_L g2143 ( 
.A(n_1815),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_L g2144 ( 
.A(n_1895),
.B(n_1232),
.Y(n_2144)
);

NAND2xp33_ASAP7_75t_L g2145 ( 
.A(n_1833),
.B(n_1545),
.Y(n_2145)
);

INVx2_ASAP7_75t_SL g2146 ( 
.A(n_1706),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_1718),
.B(n_1234),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1834),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1706),
.B(n_1265),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1697),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1718),
.B(n_1553),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1697),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_1696),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1834),
.Y(n_2154)
);

INVx4_ASAP7_75t_L g2155 ( 
.A(n_1696),
.Y(n_2155)
);

INVxp67_ASAP7_75t_L g2156 ( 
.A(n_1853),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1697),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1834),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1697),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1834),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1697),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1834),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_1700),
.Y(n_2163)
);

INVx5_ASAP7_75t_L g2164 ( 
.A(n_1833),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1718),
.B(n_1548),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1706),
.B(n_1265),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1834),
.Y(n_2167)
);

BUFx3_ASAP7_75t_L g2168 ( 
.A(n_1696),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1834),
.Y(n_2169)
);

BUFx2_ASAP7_75t_L g2170 ( 
.A(n_1853),
.Y(n_2170)
);

BUFx3_ASAP7_75t_L g2171 ( 
.A(n_1696),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1834),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1718),
.B(n_1388),
.Y(n_2173)
);

OR2x6_ASAP7_75t_L g2174 ( 
.A(n_1696),
.B(n_1008),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1697),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_1700),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1834),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1834),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1718),
.B(n_1236),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_1718),
.A2(n_1251),
.B1(n_1252),
.B2(n_1247),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_1718),
.A2(n_1457),
.B1(n_1472),
.B2(n_1470),
.Y(n_2181)
);

INVxp67_ASAP7_75t_SL g2182 ( 
.A(n_1712),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1834),
.Y(n_2183)
);

INVx4_ASAP7_75t_SL g2184 ( 
.A(n_1833),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1718),
.B(n_1254),
.Y(n_2185)
);

INVx3_ASAP7_75t_L g2186 ( 
.A(n_1700),
.Y(n_2186)
);

BUFx2_ASAP7_75t_L g2187 ( 
.A(n_1853),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_1853),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_1853),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1718),
.B(n_1256),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1834),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1834),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1834),
.Y(n_2193)
);

INVx3_ASAP7_75t_L g2194 ( 
.A(n_1700),
.Y(n_2194)
);

NOR2x1p5_ASAP7_75t_L g2195 ( 
.A(n_1700),
.B(n_1257),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1718),
.B(n_1536),
.Y(n_2196)
);

OR2x6_ASAP7_75t_L g2197 ( 
.A(n_1696),
.B(n_1008),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1697),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2059),
.B(n_1539),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1903),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1919),
.Y(n_2201)
);

AOI22xp33_ASAP7_75t_L g2202 ( 
.A1(n_2108),
.A2(n_1209),
.B1(n_1446),
.B2(n_1338),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2013),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2059),
.B(n_1259),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2017),
.Y(n_2205)
);

BUFx3_ASAP7_75t_L g2206 ( 
.A(n_2033),
.Y(n_2206)
);

AO221x1_ASAP7_75t_L g2207 ( 
.A1(n_1994),
.A2(n_1034),
.B1(n_1445),
.B2(n_1349),
.C(n_1100),
.Y(n_2207)
);

OAI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_1990),
.A2(n_1131),
.B1(n_1151),
.B2(n_1100),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2029),
.B(n_2184),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2018),
.Y(n_2210)
);

INVxp67_ASAP7_75t_L g2211 ( 
.A(n_1990),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_2085),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1963),
.B(n_1263),
.Y(n_2213)
);

AOI22xp33_ASAP7_75t_L g2214 ( 
.A1(n_2110),
.A2(n_1446),
.B1(n_1338),
.B2(n_1274),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1937),
.B(n_1275),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_1915),
.B(n_1312),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_1952),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2022),
.B(n_2072),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1915),
.B(n_1347),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2147),
.B(n_1278),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2179),
.B(n_1285),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2019),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_2006),
.B(n_1906),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1996),
.B(n_2046),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2151),
.B(n_1286),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2020),
.Y(n_2226)
);

OAI21xp33_ASAP7_75t_L g2227 ( 
.A1(n_1909),
.A2(n_1288),
.B(n_1287),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2165),
.B(n_1293),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2014),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2037),
.Y(n_2230)
);

OAI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_1996),
.A2(n_1151),
.B1(n_1184),
.B2(n_1131),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2196),
.B(n_1295),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1915),
.B(n_1373),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2065),
.B(n_1298),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_1919),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2039),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1930),
.B(n_1299),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2014),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_1918),
.B(n_1305),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2181),
.B(n_1310),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1921),
.B(n_1393),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1935),
.B(n_1311),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_2104),
.Y(n_2243)
);

HB1xp67_ASAP7_75t_L g2244 ( 
.A(n_2188),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1901),
.Y(n_2245)
);

OR2x2_ASAP7_75t_L g2246 ( 
.A(n_1932),
.B(n_1542),
.Y(n_2246)
);

INVxp33_ASAP7_75t_L g2247 ( 
.A(n_1954),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2149),
.A2(n_1329),
.B1(n_1330),
.B2(n_1317),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1989),
.B(n_1335),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1910),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2177),
.A2(n_1483),
.B(n_1478),
.Y(n_2251)
);

INVx1_ASAP7_75t_SL g2252 ( 
.A(n_2170),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1969),
.Y(n_2253)
);

OAI22xp5_ASAP7_75t_L g2254 ( 
.A1(n_1939),
.A2(n_1255),
.B1(n_1328),
.B2(n_1184),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1992),
.B(n_1341),
.Y(n_2255)
);

BUFx12f_ASAP7_75t_L g2256 ( 
.A(n_1993),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_1921),
.B(n_1342),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_SL g2258 ( 
.A(n_2058),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_1912),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_L g2260 ( 
.A(n_1949),
.B(n_1358),
.C(n_1348),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1970),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_L g2262 ( 
.A(n_2045),
.B(n_1384),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1916),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1971),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1999),
.B(n_1361),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_SL g2266 ( 
.A(n_1951),
.B(n_1255),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2012),
.B(n_1382),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2148),
.Y(n_2268)
);

AOI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_2166),
.A2(n_1402),
.B1(n_1403),
.B2(n_1398),
.Y(n_2269)
);

OAI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_1936),
.A2(n_1337),
.B1(n_1345),
.B2(n_1328),
.Y(n_2270)
);

CKINVDCx16_ASAP7_75t_R g2271 ( 
.A(n_2174),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2154),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2158),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2160),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_2102),
.Y(n_2275)
);

INVx2_ASAP7_75t_SL g2276 ( 
.A(n_1966),
.Y(n_2276)
);

INVxp33_ASAP7_75t_L g2277 ( 
.A(n_2170),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1973),
.B(n_1407),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_L g2279 ( 
.A1(n_1958),
.A2(n_1409),
.B1(n_1421),
.B2(n_1410),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1978),
.B(n_1422),
.Y(n_2280)
);

BUFx3_ASAP7_75t_L g2281 ( 
.A(n_1923),
.Y(n_2281)
);

NAND2xp33_ASAP7_75t_R g2282 ( 
.A(n_1925),
.B(n_1426),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2146),
.B(n_1430),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1979),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2162),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2167),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2057),
.A2(n_1345),
.B1(n_1349),
.B2(n_1337),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1980),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_SL g2289 ( 
.A(n_2046),
.B(n_1368),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_1962),
.A2(n_1432),
.B1(n_1436),
.B2(n_1433),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_1921),
.B(n_1441),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_2005),
.Y(n_2292)
);

INVxp33_ASAP7_75t_L g2293 ( 
.A(n_2187),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2184),
.B(n_980),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1985),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2164),
.B(n_2073),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_1988),
.B(n_1443),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1997),
.B(n_1452),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2001),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2164),
.B(n_1485),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2103),
.B(n_1460),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2002),
.B(n_1462),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2021),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2164),
.B(n_1475),
.Y(n_2304)
);

AND2x6_ASAP7_75t_SL g2305 ( 
.A(n_2075),
.B(n_1368),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2169),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_2156),
.B(n_1523),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2180),
.B(n_1466),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2172),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_1984),
.B(n_1481),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2023),
.B(n_1482),
.Y(n_2311)
);

BUFx6f_ASAP7_75t_L g2312 ( 
.A(n_2183),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_L g2313 ( 
.A1(n_1965),
.A2(n_1484),
.B1(n_1492),
.B2(n_1486),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2191),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2025),
.B(n_1496),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2187),
.B(n_1390),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2192),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_1923),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2105),
.B(n_988),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2189),
.B(n_1512),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2028),
.B(n_1550),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2189),
.B(n_961),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1934),
.B(n_1546),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2193),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1944),
.B(n_1555),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1950),
.B(n_1487),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_1943),
.B(n_964),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_1960),
.B(n_1491),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_1974),
.A2(n_1494),
.B1(n_1508),
.B2(n_1504),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2114),
.B(n_970),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_1961),
.B(n_1513),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_1938),
.A2(n_975),
.B1(n_1001),
.B2(n_982),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2054),
.B(n_1002),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_1986),
.B(n_1390),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2041),
.B(n_1517),
.Y(n_2335)
);

INVx2_ASAP7_75t_SL g2336 ( 
.A(n_2054),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_SL g2337 ( 
.A(n_2043),
.B(n_1533),
.C(n_1493),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_SL g2338 ( 
.A1(n_2115),
.A2(n_1493),
.B1(n_1533),
.B2(n_1445),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2055),
.B(n_1521),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2119),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2040),
.B(n_1524),
.Y(n_2341)
);

AOI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_1938),
.A2(n_1021),
.B1(n_1023),
.B2(n_1020),
.Y(n_2342)
);

BUFx8_ASAP7_75t_L g2343 ( 
.A(n_2143),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2007),
.Y(n_2344)
);

INVx3_ASAP7_75t_L g2345 ( 
.A(n_1946),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2007),
.B(n_1025),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_1908),
.B(n_1029),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_1977),
.Y(n_2348)
);

CKINVDCx20_ASAP7_75t_R g2349 ( 
.A(n_1993),
.Y(n_2349)
);

BUFx8_ASAP7_75t_L g2350 ( 
.A(n_2143),
.Y(n_2350)
);

NAND3xp33_ASAP7_75t_L g2351 ( 
.A(n_2109),
.B(n_1036),
.C(n_1032),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_1902),
.B(n_1041),
.Y(n_2352)
);

NAND2xp33_ASAP7_75t_L g2353 ( 
.A(n_2045),
.B(n_2049),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1982),
.Y(n_2354)
);

BUFx2_ASAP7_75t_L g2355 ( 
.A(n_2174),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1907),
.B(n_1048),
.Y(n_2356)
);

INVx2_ASAP7_75t_SL g2357 ( 
.A(n_1947),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1911),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2097),
.B(n_1050),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2150),
.B(n_1051),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2152),
.B(n_1054),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1917),
.B(n_1058),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_1946),
.B(n_1941),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_2197),
.B(n_2076),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_1946),
.B(n_1070),
.Y(n_2365)
);

INVx2_ASAP7_75t_SL g2366 ( 
.A(n_2153),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_2185),
.B(n_1006),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1987),
.Y(n_2368)
);

INVx2_ASAP7_75t_SL g2369 ( 
.A(n_2168),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2157),
.B(n_1076),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2030),
.B(n_1265),
.Y(n_2371)
);

INVxp67_ASAP7_75t_L g2372 ( 
.A(n_1983),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2159),
.B(n_1077),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_1938),
.A2(n_1088),
.B1(n_1089),
.B2(n_1078),
.Y(n_2374)
);

AND2x4_ASAP7_75t_L g2375 ( 
.A(n_2190),
.B(n_1007),
.Y(n_2375)
);

BUFx3_ASAP7_75t_L g2376 ( 
.A(n_2171),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2112),
.B(n_2182),
.Y(n_2377)
);

INVx4_ASAP7_75t_L g2378 ( 
.A(n_2004),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2161),
.B(n_1090),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2175),
.B(n_2198),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1995),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_1967),
.B(n_1009),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_2197),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2031),
.B(n_2036),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1998),
.Y(n_2385)
);

OR2x6_ASAP7_75t_L g2386 ( 
.A(n_2075),
.B(n_974),
.Y(n_2386)
);

NAND2xp33_ASAP7_75t_L g2387 ( 
.A(n_2045),
.B(n_1545),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_2064),
.B(n_1014),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2050),
.B(n_1092),
.Y(n_2389)
);

BUFx3_ASAP7_75t_L g2390 ( 
.A(n_2004),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2016),
.B(n_1097),
.Y(n_2391)
);

INVx3_ASAP7_75t_L g2392 ( 
.A(n_2000),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2078),
.B(n_1105),
.Y(n_2393)
);

INVxp67_ASAP7_75t_L g2394 ( 
.A(n_2077),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1976),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2060),
.A2(n_1110),
.B1(n_1115),
.B2(n_1108),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2079),
.B(n_1119),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_1922),
.A2(n_1126),
.B1(n_1135),
.B2(n_1124),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2077),
.B(n_999),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_1914),
.B(n_2009),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2008),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2067),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_2009),
.B(n_1138),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2177),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_1922),
.B(n_1142),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2173),
.B(n_1146),
.Y(n_2406)
);

AO22x2_ASAP7_75t_L g2407 ( 
.A1(n_2091),
.A2(n_1123),
.B1(n_1219),
.B2(n_1059),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2056),
.B(n_1147),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2089),
.B(n_1150),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_1957),
.B(n_1408),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_SL g2411 ( 
.A(n_2016),
.B(n_1152),
.Y(n_2411)
);

INVxp67_ASAP7_75t_L g2412 ( 
.A(n_2049),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2089),
.B(n_1153),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2178),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2178),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2090),
.B(n_1155),
.Y(n_2416)
);

INVxp67_ASAP7_75t_SL g2417 ( 
.A(n_2061),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1981),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_2084),
.B(n_1161),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_2080),
.B(n_2096),
.Y(n_2420)
);

NOR2xp33_ASAP7_75t_R g2421 ( 
.A(n_2140),
.B(n_1166),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2090),
.B(n_1171),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_1924),
.B(n_1178),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2116),
.B(n_1183),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2044),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2099),
.B(n_1186),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_1904),
.B(n_1188),
.Y(n_2427)
);

NOR3xp33_ASAP7_75t_L g2428 ( 
.A(n_2111),
.B(n_1551),
.C(n_1530),
.Y(n_2428)
);

INVxp67_ASAP7_75t_L g2429 ( 
.A(n_2049),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2044),
.B(n_1191),
.Y(n_2430)
);

AOI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2003),
.A2(n_1034),
.B1(n_1035),
.B2(n_1022),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2027),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_1928),
.B(n_2035),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2117),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_1926),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_1929),
.B(n_1195),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2125),
.B(n_1197),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2083),
.B(n_1200),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_1972),
.B(n_1203),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_1972),
.B(n_1208),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1926),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2094),
.B(n_1217),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2074),
.B(n_1221),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2095),
.B(n_1214),
.Y(n_2444)
);

NAND2xp33_ASAP7_75t_L g2445 ( 
.A(n_2062),
.B(n_1223),
.Y(n_2445)
);

NOR2xp67_ASAP7_75t_L g2446 ( 
.A(n_2106),
.B(n_5),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2101),
.B(n_1237),
.Y(n_2447)
);

INVx8_ASAP7_75t_L g2448 ( 
.A(n_2062),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2071),
.A2(n_1034),
.B1(n_1052),
.B2(n_1047),
.Y(n_2449)
);

NAND2xp33_ASAP7_75t_L g2450 ( 
.A(n_2062),
.B(n_1238),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2118),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2088),
.B(n_1239),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2130),
.B(n_1240),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2081),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_SL g2455 ( 
.A(n_2134),
.B(n_1241),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1940),
.B(n_1242),
.Y(n_2456)
);

INVx2_ASAP7_75t_SL g2457 ( 
.A(n_2011),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2071),
.B(n_1249),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_1905),
.B(n_1258),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2071),
.B(n_1260),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2144),
.B(n_1262),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2133),
.B(n_1269),
.Y(n_2462)
);

BUFx3_ASAP7_75t_L g2463 ( 
.A(n_2011),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_1959),
.B(n_1270),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2042),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2086),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2087),
.Y(n_2467)
);

NOR3xp33_ASAP7_75t_L g2468 ( 
.A(n_2123),
.B(n_1434),
.C(n_1413),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2113),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2034),
.B(n_1271),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2047),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2010),
.B(n_2015),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2026),
.B(n_1276),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2032),
.B(n_1313),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_1913),
.B(n_1281),
.Y(n_2475)
);

BUFx3_ASAP7_75t_L g2476 ( 
.A(n_2024),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2155),
.B(n_1282),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2093),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_SL g2479 ( 
.A(n_2163),
.B(n_2194),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2048),
.Y(n_2480)
);

NAND2xp33_ASAP7_75t_L g2481 ( 
.A(n_2100),
.B(n_1283),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2052),
.B(n_1290),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2053),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2068),
.B(n_1291),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2070),
.B(n_2092),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2176),
.B(n_1294),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_1953),
.B(n_1297),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2032),
.B(n_1313),
.Y(n_2488)
);

AOI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_1991),
.A2(n_1065),
.B1(n_1104),
.B2(n_1082),
.Y(n_2489)
);

INVx3_ASAP7_75t_L g2490 ( 
.A(n_1920),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_1975),
.B(n_1309),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_1964),
.B(n_1313),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2115),
.B(n_1464),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_SL g2494 ( 
.A(n_2082),
.B(n_1321),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_1942),
.B(n_1316),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_1931),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_1968),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2186),
.B(n_1319),
.Y(n_2498)
);

INVx2_ASAP7_75t_SL g2499 ( 
.A(n_2098),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2145),
.B(n_1326),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2082),
.B(n_1331),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_1964),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2069),
.B(n_1339),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_1933),
.B(n_1344),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_1945),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2195),
.B(n_1321),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2051),
.B(n_1346),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_1955),
.B(n_1956),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2024),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2063),
.B(n_1125),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2127),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2135),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_2119),
.B(n_1353),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2038),
.B(n_1357),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_1927),
.B(n_1359),
.Y(n_2515)
);

INVxp33_ASAP7_75t_L g2516 ( 
.A(n_1948),
.Y(n_2516)
);

NAND2xp33_ASAP7_75t_L g2517 ( 
.A(n_2132),
.B(n_1362),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2066),
.B(n_1366),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2132),
.B(n_1364),
.Y(n_2519)
);

O2A1O1Ixp33_ASAP7_75t_L g2520 ( 
.A1(n_2124),
.A2(n_1130),
.B(n_1133),
.C(n_1132),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2138),
.B(n_1369),
.Y(n_2521)
);

CKINVDCx11_ASAP7_75t_R g2522 ( 
.A(n_2107),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2121),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2122),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2128),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2136),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2142),
.B(n_1370),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2120),
.B(n_1371),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2126),
.B(n_1321),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_2129),
.B(n_1379),
.Y(n_2530)
);

BUFx2_ASAP7_75t_L g2531 ( 
.A(n_2131),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2137),
.B(n_1386),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_2139),
.B(n_1391),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2141),
.B(n_1392),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_1903),
.Y(n_2535)
);

INVxp67_ASAP7_75t_L g2536 ( 
.A(n_1990),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_1915),
.B(n_1395),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_R g2538 ( 
.A(n_2085),
.B(n_1399),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_1915),
.B(n_1401),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2013),
.Y(n_2540)
);

INVxp67_ASAP7_75t_R g2541 ( 
.A(n_1937),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2059),
.B(n_1404),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_1915),
.B(n_1411),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_1903),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_1915),
.B(n_1412),
.Y(n_2545)
);

BUFx12f_ASAP7_75t_SL g2546 ( 
.A(n_2075),
.Y(n_2546)
);

NAND2xp33_ASAP7_75t_L g2547 ( 
.A(n_2045),
.B(n_1414),
.Y(n_2547)
);

BUFx3_ASAP7_75t_L g2548 ( 
.A(n_2033),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_1990),
.B(n_1367),
.Y(n_2549)
);

AOI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2108),
.A2(n_1143),
.B1(n_1144),
.B2(n_1139),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2013),
.Y(n_2551)
);

AOI221xp5_ASAP7_75t_L g2552 ( 
.A1(n_1936),
.A2(n_1157),
.B1(n_1172),
.B2(n_1170),
.C(n_1165),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2059),
.B(n_1415),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2059),
.B(n_1419),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_1903),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_1903),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1903),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_1903),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2059),
.B(n_1420),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_1915),
.B(n_1424),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_1903),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2013),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_2059),
.B(n_1176),
.Y(n_2563)
);

NOR2xp67_ASAP7_75t_L g2564 ( 
.A(n_1915),
.B(n_5),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2188),
.B(n_1425),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2059),
.B(n_1431),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2059),
.B(n_1439),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2059),
.B(n_1442),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2059),
.B(n_1447),
.Y(n_2569)
);

INVx4_ASAP7_75t_L g2570 ( 
.A(n_2004),
.Y(n_2570)
);

NAND2xp33_ASAP7_75t_L g2571 ( 
.A(n_2045),
.B(n_1449),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2059),
.B(n_1451),
.Y(n_2572)
);

AO21x1_ASAP7_75t_L g2573 ( 
.A1(n_2435),
.A2(n_1185),
.B(n_1179),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2218),
.B(n_1454),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_L g2575 ( 
.A(n_2247),
.B(n_1455),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2277),
.B(n_1456),
.Y(n_2576)
);

INVx4_ASAP7_75t_L g2577 ( 
.A(n_2256),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_L g2578 ( 
.A(n_2293),
.B(n_1467),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2200),
.B(n_1471),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2535),
.B(n_1473),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2252),
.B(n_1479),
.Y(n_2581)
);

INVx4_ASAP7_75t_L g2582 ( 
.A(n_2448),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2544),
.B(n_1488),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2211),
.B(n_1489),
.Y(n_2584)
);

NAND2x1p5_ASAP7_75t_L g2585 ( 
.A(n_2463),
.B(n_1019),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2555),
.B(n_1490),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2536),
.B(n_1497),
.Y(n_2587)
);

OAI321xp33_ASAP7_75t_L g2588 ( 
.A1(n_2270),
.A2(n_1202),
.A3(n_1215),
.B1(n_1246),
.B2(n_1228),
.C(n_1205),
.Y(n_2588)
);

BUFx8_ASAP7_75t_L g2589 ( 
.A(n_2258),
.Y(n_2589)
);

OAI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_2251),
.A2(n_1267),
.B(n_1261),
.Y(n_2590)
);

AOI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2289),
.A2(n_1498),
.B1(n_1516),
.B2(n_1514),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2384),
.A2(n_1284),
.B(n_1277),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2224),
.B(n_1367),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2420),
.A2(n_1300),
.B(n_1289),
.Y(n_2594)
);

A2O1A1Ixp33_ASAP7_75t_L g2595 ( 
.A1(n_2446),
.A2(n_1303),
.B(n_1304),
.C(n_1302),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2556),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2557),
.B(n_1522),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2404),
.A2(n_1318),
.B(n_1315),
.Y(n_2598)
);

OAI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2441),
.A2(n_1336),
.B(n_1320),
.Y(n_2599)
);

OAI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2213),
.A2(n_1354),
.B(n_1340),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2246),
.B(n_1367),
.Y(n_2601)
);

NAND2x1_ASAP7_75t_L g2602 ( 
.A(n_2340),
.B(n_1019),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_SL g2603 ( 
.A(n_2244),
.B(n_1538),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2364),
.B(n_1525),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2316),
.B(n_1526),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2558),
.B(n_1532),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2561),
.B(n_1534),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_2414),
.A2(n_1375),
.B(n_1374),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2253),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2415),
.A2(n_1378),
.B(n_1377),
.Y(n_2610)
);

O2A1O1Ixp33_ASAP7_75t_SL g2611 ( 
.A1(n_2229),
.A2(n_1394),
.B(n_1396),
.C(n_1389),
.Y(n_2611)
);

INVx3_ASAP7_75t_L g2612 ( 
.A(n_2378),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2563),
.B(n_1540),
.Y(n_2613)
);

AOI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2199),
.A2(n_1400),
.B(n_1397),
.Y(n_2614)
);

O2A1O1Ixp33_ASAP7_75t_L g2615 ( 
.A1(n_2204),
.A2(n_1406),
.B(n_1423),
.C(n_1405),
.Y(n_2615)
);

O2A1O1Ixp33_ASAP7_75t_L g2616 ( 
.A1(n_2220),
.A2(n_1438),
.B(n_1458),
.C(n_1427),
.Y(n_2616)
);

INVx1_ASAP7_75t_SL g2617 ( 
.A(n_2250),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2377),
.B(n_1541),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2261),
.Y(n_2619)
);

AND2x6_ASAP7_75t_L g2620 ( 
.A(n_2238),
.B(n_974),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2264),
.Y(n_2621)
);

OAI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2563),
.A2(n_1549),
.B1(n_1554),
.B2(n_1544),
.Y(n_2622)
);

OAI21xp33_ASAP7_75t_L g2623 ( 
.A1(n_2215),
.A2(n_1505),
.B(n_1477),
.Y(n_2623)
);

OAI21xp33_ASAP7_75t_L g2624 ( 
.A1(n_2225),
.A2(n_1509),
.B(n_1506),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2284),
.B(n_1510),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2288),
.B(n_1515),
.Y(n_2626)
);

AOI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2337),
.A2(n_1527),
.B1(n_1528),
.B2(n_1518),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2245),
.A2(n_1531),
.B(n_1529),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2295),
.B(n_1245),
.Y(n_2629)
);

AOI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2268),
.A2(n_2273),
.B(n_2272),
.Y(n_2630)
);

OAI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2274),
.A2(n_1250),
.B(n_1245),
.Y(n_2631)
);

AOI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2285),
.A2(n_2306),
.B(n_2286),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2380),
.A2(n_1323),
.B1(n_1355),
.B2(n_1250),
.Y(n_2633)
);

NOR2xp67_ASAP7_75t_L g2634 ( 
.A(n_2372),
.B(n_4),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2217),
.B(n_1019),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2334),
.B(n_1323),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2276),
.B(n_1019),
.Y(n_2637)
);

A2O1A1Ixp33_ASAP7_75t_L g2638 ( 
.A1(n_2446),
.A2(n_1355),
.B(n_1468),
.C(n_1448),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2340),
.B(n_2266),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2254),
.A2(n_1448),
.B1(n_1511),
.B2(n_1468),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2299),
.B(n_1511),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2340),
.B(n_2332),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2303),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2321),
.B(n_4),
.Y(n_2644)
);

INVx3_ASAP7_75t_L g2645 ( 
.A(n_2378),
.Y(n_2645)
);

AOI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2309),
.A2(n_1474),
.B(n_1196),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2329),
.B(n_2341),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2314),
.A2(n_1474),
.B(n_1196),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2355),
.B(n_4),
.Y(n_2649)
);

O2A1O1Ixp33_ASAP7_75t_L g2650 ( 
.A1(n_2221),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_2650)
);

AOI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2367),
.A2(n_1474),
.B1(n_1196),
.B2(n_8),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2343),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2317),
.A2(n_1474),
.B(n_1196),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2541),
.B(n_6),
.Y(n_2654)
);

OAI21xp33_ASAP7_75t_L g2655 ( 
.A1(n_2228),
.A2(n_6),
.B(n_7),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2324),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2542),
.B(n_8),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_R g2658 ( 
.A(n_2546),
.B(n_8),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2201),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2208),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2342),
.B(n_10),
.Y(n_2661)
);

AND2x6_ASAP7_75t_L g2662 ( 
.A(n_2209),
.B(n_9),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2553),
.B(n_10),
.Y(n_2663)
);

INVx8_ASAP7_75t_L g2664 ( 
.A(n_2448),
.Y(n_2664)
);

OAI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2402),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2203),
.Y(n_2666)
);

OAI21xp5_ASAP7_75t_L g2667 ( 
.A1(n_2554),
.A2(n_11),
.B(n_12),
.Y(n_2667)
);

AND2x4_ASAP7_75t_L g2668 ( 
.A(n_2209),
.B(n_12),
.Y(n_2668)
);

OAI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2559),
.A2(n_13),
.B(n_14),
.Y(n_2669)
);

INVxp67_ASAP7_75t_L g2670 ( 
.A(n_2282),
.Y(n_2670)
);

AOI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2232),
.A2(n_13),
.B(n_14),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2374),
.B(n_15),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2549),
.B(n_14),
.Y(n_2673)
);

AOI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2566),
.A2(n_15),
.B(n_16),
.Y(n_2674)
);

BUFx2_ASAP7_75t_L g2675 ( 
.A(n_2343),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2567),
.B(n_15),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2568),
.B(n_16),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2569),
.B(n_16),
.Y(n_2678)
);

BUFx3_ASAP7_75t_L g2679 ( 
.A(n_2349),
.Y(n_2679)
);

OAI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2572),
.A2(n_17),
.B(n_18),
.Y(n_2680)
);

INVx3_ASAP7_75t_L g2681 ( 
.A(n_2570),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2223),
.B(n_17),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2335),
.B(n_17),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_2485),
.A2(n_18),
.B(n_19),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2205),
.Y(n_2685)
);

OAI321xp33_ASAP7_75t_L g2686 ( 
.A1(n_2474),
.A2(n_20),
.A3(n_22),
.B1(n_18),
.B2(n_19),
.C(n_21),
.Y(n_2686)
);

OAI21xp5_ASAP7_75t_L g2687 ( 
.A1(n_2234),
.A2(n_19),
.B(n_20),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2339),
.B(n_21),
.Y(n_2688)
);

AOI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2242),
.A2(n_21),
.B(n_22),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2249),
.B(n_2255),
.Y(n_2690)
);

OAI21xp5_ASAP7_75t_L g2691 ( 
.A1(n_2265),
.A2(n_2267),
.B(n_2344),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2278),
.B(n_22),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2280),
.B(n_24),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2297),
.B(n_24),
.Y(n_2694)
);

BUFx6f_ASAP7_75t_L g2695 ( 
.A(n_2201),
.Y(n_2695)
);

OAI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2489),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2298),
.A2(n_25),
.B(n_26),
.Y(n_2697)
);

AOI21x1_ASAP7_75t_L g2698 ( 
.A1(n_2564),
.A2(n_25),
.B(n_26),
.Y(n_2698)
);

AOI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2302),
.A2(n_27),
.B(n_28),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2311),
.B(n_27),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2371),
.B(n_28),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2210),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2315),
.A2(n_29),
.B(n_30),
.Y(n_2703)
);

BUFx12f_ASAP7_75t_L g2704 ( 
.A(n_2305),
.Y(n_2704)
);

NAND2x1_ASAP7_75t_L g2705 ( 
.A(n_2570),
.B(n_29),
.Y(n_2705)
);

AOI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2389),
.A2(n_29),
.B(n_31),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2240),
.B(n_31),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2222),
.Y(n_2708)
);

BUFx2_ASAP7_75t_L g2709 ( 
.A(n_2350),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2231),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2226),
.Y(n_2711)
);

NAND3xp33_ASAP7_75t_L g2712 ( 
.A(n_2424),
.B(n_32),
.C(n_33),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2201),
.Y(n_2713)
);

NOR2xp67_ASAP7_75t_L g2714 ( 
.A(n_2260),
.B(n_32),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2230),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2338),
.B(n_33),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2390),
.Y(n_2717)
);

O2A1O1Ixp33_ASAP7_75t_L g2718 ( 
.A1(n_2237),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2367),
.B(n_2375),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2508),
.A2(n_34),
.B(n_35),
.Y(n_2720)
);

AO21x1_ASAP7_75t_L g2721 ( 
.A1(n_2387),
.A2(n_579),
.B(n_578),
.Y(n_2721)
);

O2A1O1Ixp33_ASAP7_75t_L g2722 ( 
.A1(n_2488),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2350),
.Y(n_2723)
);

O2A1O1Ixp33_ASAP7_75t_L g2724 ( 
.A1(n_2410),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2724)
);

AOI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2327),
.A2(n_37),
.B(n_38),
.Y(n_2725)
);

AOI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2346),
.A2(n_39),
.B(n_40),
.Y(n_2726)
);

AOI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2453),
.A2(n_39),
.B(n_40),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2320),
.B(n_40),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2375),
.B(n_41),
.Y(n_2729)
);

AOI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_2323),
.A2(n_41),
.B(n_42),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2248),
.B(n_41),
.Y(n_2731)
);

A2O1A1Ixp33_ASAP7_75t_L g2732 ( 
.A1(n_2520),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2550),
.B(n_43),
.Y(n_2733)
);

AOI21xp5_ASAP7_75t_L g2734 ( 
.A1(n_2325),
.A2(n_45),
.B(n_46),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2489),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2235),
.Y(n_2736)
);

AO21x1_ASAP7_75t_L g2737 ( 
.A1(n_2353),
.A2(n_580),
.B(n_579),
.Y(n_2737)
);

NOR2xp67_ASAP7_75t_L g2738 ( 
.A(n_2564),
.B(n_45),
.Y(n_2738)
);

AOI21xp5_ASAP7_75t_L g2739 ( 
.A1(n_2326),
.A2(n_2331),
.B(n_2328),
.Y(n_2739)
);

NOR2xp33_ASAP7_75t_L g2740 ( 
.A(n_2394),
.B(n_47),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2358),
.B(n_48),
.Y(n_2741)
);

O2A1O1Ixp33_ASAP7_75t_L g2742 ( 
.A1(n_2308),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2236),
.Y(n_2743)
);

AOI21xp5_ASAP7_75t_L g2744 ( 
.A1(n_2259),
.A2(n_48),
.B(n_49),
.Y(n_2744)
);

AOI21xp33_ASAP7_75t_L g2745 ( 
.A1(n_2403),
.A2(n_49),
.B(n_50),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2540),
.Y(n_2746)
);

A2O1A1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_2227),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_2747)
);

OAI321xp33_ASAP7_75t_L g2748 ( 
.A1(n_2386),
.A2(n_53),
.A3(n_55),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2565),
.B(n_53),
.Y(n_2749)
);

BUFx4_ASAP7_75t_SL g2750 ( 
.A(n_2206),
.Y(n_2750)
);

A2O1A1Ixp33_ASAP7_75t_L g2751 ( 
.A1(n_2443),
.A2(n_55),
.B(n_52),
.C(n_53),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2269),
.B(n_55),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2388),
.B(n_56),
.Y(n_2753)
);

NOR2x1_ASAP7_75t_R g2754 ( 
.A(n_2383),
.B(n_56),
.Y(n_2754)
);

AOI21xp5_ASAP7_75t_L g2755 ( 
.A1(n_2259),
.A2(n_56),
.B(n_57),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2259),
.A2(n_58),
.B(n_59),
.Y(n_2756)
);

OR2x6_ASAP7_75t_L g2757 ( 
.A(n_2448),
.B(n_58),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2388),
.B(n_59),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2279),
.B(n_60),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2493),
.B(n_60),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2290),
.B(n_60),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2263),
.A2(n_61),
.B(n_62),
.Y(n_2762)
);

AOI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2263),
.A2(n_2312),
.B(n_2514),
.Y(n_2763)
);

BUFx8_ASAP7_75t_SL g2764 ( 
.A(n_2258),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2313),
.B(n_61),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2214),
.B(n_62),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2312),
.A2(n_2426),
.B(n_2362),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2407),
.B(n_63),
.Y(n_2768)
);

O2A1O1Ixp33_ASAP7_75t_L g2769 ( 
.A1(n_2437),
.A2(n_66),
.B(n_63),
.C(n_65),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2454),
.B(n_65),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2466),
.B(n_2467),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2235),
.Y(n_2772)
);

O2A1O1Ixp33_ASAP7_75t_L g2773 ( 
.A1(n_2399),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2551),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2347),
.A2(n_67),
.B(n_68),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2212),
.Y(n_2776)
);

BUFx6f_ASAP7_75t_L g2777 ( 
.A(n_2235),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_2322),
.B(n_67),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2562),
.Y(n_2779)
);

AOI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2352),
.A2(n_68),
.B(n_69),
.Y(n_2780)
);

AOI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2356),
.A2(n_2361),
.B(n_2360),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2478),
.B(n_69),
.Y(n_2782)
);

INVx3_ASAP7_75t_L g2783 ( 
.A(n_2345),
.Y(n_2783)
);

AOI21xp5_ASAP7_75t_L g2784 ( 
.A1(n_2370),
.A2(n_2379),
.B(n_2373),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2552),
.B(n_69),
.Y(n_2785)
);

AOI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2452),
.A2(n_70),
.B(n_71),
.Y(n_2786)
);

AOI21xp5_ASAP7_75t_L g2787 ( 
.A1(n_2472),
.A2(n_70),
.B(n_71),
.Y(n_2787)
);

AOI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2495),
.A2(n_72),
.B(n_73),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2345),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2393),
.B(n_72),
.Y(n_2790)
);

AO21x1_ASAP7_75t_L g2791 ( 
.A1(n_2363),
.A2(n_582),
.B(n_581),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2397),
.B(n_73),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2500),
.A2(n_74),
.B(n_75),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2359),
.B(n_74),
.Y(n_2794)
);

INVxp67_ASAP7_75t_L g2795 ( 
.A(n_2386),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2529),
.B(n_74),
.Y(n_2796)
);

AOI21xp33_ASAP7_75t_L g2797 ( 
.A1(n_2301),
.A2(n_75),
.B(n_76),
.Y(n_2797)
);

NAND2xp33_ASAP7_75t_L g2798 ( 
.A(n_2457),
.B(n_2336),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2348),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2468),
.B(n_76),
.Y(n_2800)
);

CKINVDCx5p33_ASAP7_75t_R g2801 ( 
.A(n_2243),
.Y(n_2801)
);

INVxp67_ASAP7_75t_L g2802 ( 
.A(n_2310),
.Y(n_2802)
);

O2A1O1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_2515),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_2803)
);

AOI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2482),
.A2(n_78),
.B(n_79),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2354),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2368),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2307),
.B(n_79),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2281),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2425),
.B(n_80),
.Y(n_2809)
);

OAI21xp5_ASAP7_75t_L g2810 ( 
.A1(n_2483),
.A2(n_80),
.B(n_81),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_2275),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_SL g2812 ( 
.A(n_2271),
.B(n_81),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2510),
.B(n_80),
.Y(n_2813)
);

INVx2_ASAP7_75t_SL g2814 ( 
.A(n_2548),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2484),
.A2(n_82),
.B(n_83),
.Y(n_2815)
);

BUFx6f_ASAP7_75t_L g2816 ( 
.A(n_2318),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2524),
.A2(n_82),
.B(n_83),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2526),
.A2(n_82),
.B(n_83),
.Y(n_2818)
);

AOI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2465),
.A2(n_84),
.B(n_85),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2471),
.A2(n_84),
.B(n_85),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_SL g2821 ( 
.A(n_2494),
.B(n_85),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2480),
.A2(n_84),
.B(n_86),
.Y(n_2822)
);

AOI21xp33_ASAP7_75t_L g2823 ( 
.A1(n_2239),
.A2(n_86),
.B(n_87),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2381),
.A2(n_86),
.B(n_88),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2385),
.Y(n_2825)
);

BUFx2_ASAP7_75t_L g2826 ( 
.A(n_2538),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2401),
.A2(n_88),
.B(n_89),
.Y(n_2827)
);

AOI21xp5_ASAP7_75t_L g2828 ( 
.A1(n_2497),
.A2(n_88),
.B(n_89),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2433),
.A2(n_90),
.B(n_91),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2510),
.B(n_90),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2407),
.B(n_91),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2496),
.A2(n_91),
.B(n_92),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2505),
.A2(n_92),
.B(n_93),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2523),
.A2(n_92),
.B(n_93),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2392),
.Y(n_2835)
);

OAI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2351),
.A2(n_94),
.B(n_95),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2525),
.A2(n_94),
.B(n_95),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2528),
.A2(n_94),
.B(n_95),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2319),
.B(n_2283),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2427),
.A2(n_96),
.B(n_97),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2395),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2319),
.B(n_96),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2287),
.B(n_97),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2434),
.B(n_2451),
.Y(n_2844)
);

OAI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2392),
.A2(n_97),
.B(n_98),
.Y(n_2845)
);

AO21x1_ASAP7_75t_L g2846 ( 
.A1(n_2262),
.A2(n_583),
.B(n_581),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2506),
.B(n_2418),
.Y(n_2847)
);

BUFx6f_ASAP7_75t_L g2848 ( 
.A(n_2522),
.Y(n_2848)
);

AOI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2330),
.A2(n_98),
.B(n_99),
.Y(n_2849)
);

AOI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2461),
.A2(n_99),
.B(n_100),
.Y(n_2850)
);

AOI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2406),
.A2(n_99),
.B(n_100),
.Y(n_2851)
);

OAI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2202),
.A2(n_100),
.B(n_101),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2481),
.B(n_101),
.Y(n_2853)
);

AOI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2207),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2432),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2408),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2398),
.B(n_102),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2456),
.A2(n_102),
.B(n_104),
.Y(n_2858)
);

BUFx3_ASAP7_75t_L g2859 ( 
.A(n_2376),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2503),
.B(n_104),
.Y(n_2860)
);

INVxp67_ASAP7_75t_L g2861 ( 
.A(n_2405),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2502),
.B(n_105),
.Y(n_2862)
);

AND2x4_ASAP7_75t_L g2863 ( 
.A(n_2417),
.B(n_106),
.Y(n_2863)
);

AOI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2487),
.A2(n_106),
.B(n_107),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2400),
.B(n_107),
.Y(n_2865)
);

AOI22xp33_ASAP7_75t_L g2866 ( 
.A1(n_2382),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2409),
.B(n_109),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2431),
.B(n_108),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2382),
.B(n_108),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2490),
.Y(n_2870)
);

NOR3xp33_ASAP7_75t_L g2871 ( 
.A(n_2428),
.B(n_112),
.C(n_111),
.Y(n_2871)
);

AOI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2491),
.A2(n_110),
.B(n_111),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2423),
.B(n_110),
.Y(n_2873)
);

INVx6_ASAP7_75t_L g2874 ( 
.A(n_2476),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2436),
.B(n_110),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2438),
.A2(n_111),
.B(n_112),
.Y(n_2876)
);

BUFx6f_ASAP7_75t_L g2877 ( 
.A(n_2531),
.Y(n_2877)
);

BUFx6f_ASAP7_75t_L g2878 ( 
.A(n_2511),
.Y(n_2878)
);

AO21x1_ASAP7_75t_L g2879 ( 
.A1(n_2547),
.A2(n_586),
.B(n_584),
.Y(n_2879)
);

AND2x4_ASAP7_75t_L g2880 ( 
.A(n_2412),
.B(n_112),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2430),
.B(n_2492),
.Y(n_2881)
);

BUFx4f_ASAP7_75t_L g2882 ( 
.A(n_2499),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2504),
.B(n_113),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2490),
.Y(n_2884)
);

BUFx6f_ASAP7_75t_L g2885 ( 
.A(n_2512),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2294),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2419),
.B(n_113),
.Y(n_2887)
);

OAI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2444),
.A2(n_114),
.B(n_115),
.Y(n_2888)
);

O2A1O1Ixp33_ASAP7_75t_L g2889 ( 
.A1(n_2571),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2889)
);

OR2x2_ASAP7_75t_L g2890 ( 
.A(n_2396),
.B(n_115),
.Y(n_2890)
);

AND2x2_ASAP7_75t_SL g2891 ( 
.A(n_2445),
.B(n_116),
.Y(n_2891)
);

A2O1A1Ixp33_ASAP7_75t_L g2892 ( 
.A1(n_2449),
.A2(n_121),
.B(n_117),
.C(n_118),
.Y(n_2892)
);

AND2x6_ASAP7_75t_L g2893 ( 
.A(n_2294),
.B(n_117),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2442),
.B(n_117),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_L g2895 ( 
.A(n_2462),
.B(n_118),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_SL g2896 ( 
.A(n_2413),
.B(n_121),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2459),
.B(n_118),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2509),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_SL g2899 ( 
.A(n_2292),
.B(n_122),
.Y(n_2899)
);

AOI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_2447),
.A2(n_122),
.B(n_123),
.Y(n_2900)
);

AND2x4_ASAP7_75t_L g2901 ( 
.A(n_2429),
.B(n_122),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2473),
.A2(n_123),
.B(n_124),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2521),
.Y(n_2903)
);

OAI321xp33_ASAP7_75t_L g2904 ( 
.A1(n_2518),
.A2(n_126),
.A3(n_128),
.B1(n_124),
.B2(n_125),
.C(n_127),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2455),
.A2(n_124),
.B(n_125),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_2333),
.B(n_2498),
.Y(n_2906)
);

HB1xp67_ASAP7_75t_L g2907 ( 
.A(n_2357),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2216),
.Y(n_2908)
);

OAI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2470),
.A2(n_126),
.B(n_127),
.Y(n_2909)
);

AO21x1_ASAP7_75t_L g2910 ( 
.A1(n_2458),
.A2(n_588),
.B(n_587),
.Y(n_2910)
);

AOI21x1_ASAP7_75t_L g2911 ( 
.A1(n_2219),
.A2(n_126),
.B(n_127),
.Y(n_2911)
);

BUFx2_ASAP7_75t_L g2912 ( 
.A(n_2469),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2416),
.B(n_128),
.Y(n_2913)
);

INVx2_ASAP7_75t_SL g2914 ( 
.A(n_2366),
.Y(n_2914)
);

BUFx4f_ASAP7_75t_L g2915 ( 
.A(n_2369),
.Y(n_2915)
);

AOI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2460),
.A2(n_128),
.B(n_129),
.Y(n_2916)
);

INVx3_ASAP7_75t_L g2917 ( 
.A(n_2422),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2421),
.B(n_130),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2464),
.B(n_129),
.Y(n_2919)
);

INVxp67_ASAP7_75t_L g2920 ( 
.A(n_2450),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2527),
.B(n_129),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2296),
.A2(n_130),
.B(n_131),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_SL g2923 ( 
.A(n_2516),
.B(n_132),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2530),
.Y(n_2924)
);

OAI21xp33_ASAP7_75t_L g2925 ( 
.A1(n_2507),
.A2(n_131),
.B(n_132),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2486),
.B(n_132),
.Y(n_2926)
);

AOI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2233),
.A2(n_133),
.B(n_134),
.Y(n_2927)
);

INVx1_ASAP7_75t_SL g2928 ( 
.A(n_2517),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2241),
.A2(n_133),
.B(n_134),
.Y(n_2929)
);

AOI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2257),
.A2(n_133),
.B(n_134),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2475),
.B(n_135),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_R g2932 ( 
.A(n_2532),
.B(n_135),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2477),
.B(n_135),
.Y(n_2933)
);

AOI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2291),
.A2(n_136),
.B(n_137),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_SL g2935 ( 
.A(n_2533),
.B(n_137),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2534),
.B(n_136),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2391),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2439),
.B(n_138),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2300),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2411),
.B(n_139),
.Y(n_2940)
);

O2A1O1Ixp33_ASAP7_75t_L g2941 ( 
.A1(n_2501),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_2941)
);

AOI22xp33_ASAP7_75t_L g2942 ( 
.A1(n_2440),
.A2(n_2304),
.B1(n_2365),
.B2(n_2479),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2513),
.Y(n_2943)
);

AOI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2537),
.A2(n_140),
.B(n_142),
.Y(n_2944)
);

INVx3_ASAP7_75t_L g2945 ( 
.A(n_2539),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2543),
.A2(n_140),
.B(n_142),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2519),
.B(n_142),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2545),
.B(n_143),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2560),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2218),
.B(n_144),
.Y(n_2950)
);

BUFx6f_ASAP7_75t_L g2951 ( 
.A(n_2340),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2218),
.A2(n_143),
.B(n_144),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2247),
.B(n_143),
.Y(n_2953)
);

AOI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2218),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2218),
.B(n_145),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2218),
.B(n_146),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2218),
.B(n_147),
.Y(n_2957)
);

AOI21x1_ASAP7_75t_L g2958 ( 
.A1(n_2435),
.A2(n_147),
.B(n_148),
.Y(n_2958)
);

OAI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2218),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2218),
.B(n_148),
.Y(n_2960)
);

BUFx6f_ASAP7_75t_L g2961 ( 
.A(n_2340),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2247),
.B(n_149),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2218),
.A2(n_149),
.B(n_150),
.Y(n_2963)
);

OAI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2218),
.A2(n_150),
.B(n_151),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2218),
.B(n_151),
.Y(n_2965)
);

OAI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2218),
.A2(n_151),
.B(n_152),
.Y(n_2966)
);

AOI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2218),
.A2(n_152),
.B(n_153),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_2218),
.B(n_153),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2218),
.A2(n_152),
.B(n_153),
.Y(n_2969)
);

NOR2xp33_ASAP7_75t_L g2970 ( 
.A(n_2247),
.B(n_154),
.Y(n_2970)
);

AOI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2289),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2971)
);

OAI21xp5_ASAP7_75t_L g2972 ( 
.A1(n_2218),
.A2(n_155),
.B(n_157),
.Y(n_2972)
);

AOI21xp5_ASAP7_75t_L g2973 ( 
.A1(n_2218),
.A2(n_155),
.B(n_157),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2200),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2200),
.Y(n_2975)
);

BUFx3_ASAP7_75t_L g2976 ( 
.A(n_2256),
.Y(n_2976)
);

BUFx4f_ASAP7_75t_L g2977 ( 
.A(n_2256),
.Y(n_2977)
);

HB1xp67_ASAP7_75t_L g2978 ( 
.A(n_2244),
.Y(n_2978)
);

O2A1O1Ixp5_ASAP7_75t_L g2979 ( 
.A1(n_2420),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2218),
.B(n_158),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2247),
.B(n_158),
.Y(n_2981)
);

O2A1O1Ixp33_ASAP7_75t_L g2982 ( 
.A1(n_2218),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2982)
);

BUFx3_ASAP7_75t_L g2983 ( 
.A(n_2256),
.Y(n_2983)
);

AOI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2218),
.A2(n_159),
.B(n_160),
.Y(n_2984)
);

O2A1O1Ixp33_ASAP7_75t_L g2985 ( 
.A1(n_2218),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2218),
.B(n_163),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2218),
.B(n_162),
.Y(n_2987)
);

O2A1O1Ixp33_ASAP7_75t_L g2988 ( 
.A1(n_2218),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2218),
.B(n_165),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2218),
.B(n_167),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2218),
.A2(n_167),
.B(n_168),
.Y(n_2991)
);

AOI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_2289),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2218),
.B(n_170),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_2200),
.B(n_169),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2247),
.B(n_169),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_SL g2996 ( 
.A(n_2218),
.B(n_172),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2404),
.Y(n_2997)
);

AOI21xp5_ASAP7_75t_L g2998 ( 
.A1(n_2218),
.A2(n_171),
.B(n_172),
.Y(n_2998)
);

AOI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2218),
.A2(n_171),
.B(n_173),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2200),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2218),
.B(n_173),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2218),
.B(n_174),
.Y(n_3002)
);

O2A1O1Ixp33_ASAP7_75t_L g3003 ( 
.A1(n_2218),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_3003)
);

OAI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2218),
.A2(n_175),
.B(n_176),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2218),
.A2(n_175),
.B(n_177),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2218),
.B(n_177),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2218),
.B(n_177),
.Y(n_3007)
);

O2A1O1Ixp5_ASAP7_75t_L g3008 ( 
.A1(n_2420),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_3008)
);

AND2x4_ASAP7_75t_L g3009 ( 
.A(n_2200),
.B(n_179),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2218),
.B(n_181),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2404),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2218),
.B(n_181),
.Y(n_3012)
);

NOR2x1_ASAP7_75t_L g3013 ( 
.A(n_2349),
.B(n_180),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2218),
.B(n_180),
.Y(n_3014)
);

O2A1O1Ixp5_ASAP7_75t_SL g3015 ( 
.A1(n_2391),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2247),
.B(n_182),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2218),
.B(n_182),
.Y(n_3017)
);

AOI21x1_ASAP7_75t_L g3018 ( 
.A1(n_2435),
.A2(n_184),
.B(n_185),
.Y(n_3018)
);

AOI21xp5_ASAP7_75t_L g3019 ( 
.A1(n_2218),
.A2(n_184),
.B(n_185),
.Y(n_3019)
);

AOI21xp5_ASAP7_75t_L g3020 ( 
.A1(n_2218),
.A2(n_184),
.B(n_185),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2200),
.Y(n_3021)
);

AOI21xp5_ASAP7_75t_L g3022 ( 
.A1(n_2218),
.A2(n_186),
.B(n_187),
.Y(n_3022)
);

NOR2xp67_ASAP7_75t_L g3023 ( 
.A(n_2218),
.B(n_186),
.Y(n_3023)
);

OAI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2218),
.A2(n_189),
.B1(n_186),
.B2(n_188),
.Y(n_3024)
);

OAI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2218),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2404),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2200),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2200),
.Y(n_3028)
);

OAI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2218),
.A2(n_190),
.B(n_191),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2247),
.B(n_190),
.Y(n_3030)
);

AND2x4_ASAP7_75t_L g3031 ( 
.A(n_2200),
.B(n_191),
.Y(n_3031)
);

AOI33xp33_ASAP7_75t_L g3032 ( 
.A1(n_2550),
.A2(n_193),
.A3(n_195),
.B1(n_191),
.B2(n_192),
.B3(n_194),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2218),
.B(n_192),
.Y(n_3033)
);

NOR2xp33_ASAP7_75t_L g3034 ( 
.A(n_2247),
.B(n_192),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2218),
.B(n_193),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2218),
.A2(n_193),
.B(n_194),
.Y(n_3036)
);

INVx4_ASAP7_75t_L g3037 ( 
.A(n_2256),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2218),
.B(n_195),
.Y(n_3038)
);

BUFx2_ASAP7_75t_SL g3039 ( 
.A(n_2349),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2404),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2218),
.B(n_197),
.Y(n_3041)
);

AOI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2218),
.A2(n_198),
.B(n_199),
.Y(n_3042)
);

OAI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2218),
.A2(n_198),
.B(n_200),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2218),
.A2(n_198),
.B(n_201),
.Y(n_3044)
);

HB1xp67_ASAP7_75t_L g3045 ( 
.A(n_2244),
.Y(n_3045)
);

AOI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2218),
.A2(n_201),
.B(n_202),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2218),
.B(n_202),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2200),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2218),
.B(n_203),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_SL g3050 ( 
.A(n_2546),
.B(n_203),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2200),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2218),
.A2(n_203),
.B(n_204),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2218),
.B(n_205),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2218),
.B(n_205),
.Y(n_3054)
);

OAI21xp33_ASAP7_75t_L g3055 ( 
.A1(n_2218),
.A2(n_205),
.B(n_206),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2218),
.B(n_206),
.Y(n_3056)
);

OAI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2218),
.A2(n_206),
.B(n_207),
.Y(n_3057)
);

INVx5_ASAP7_75t_L g3058 ( 
.A(n_2340),
.Y(n_3058)
);

INVxp67_ASAP7_75t_SL g3059 ( 
.A(n_2218),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2200),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2200),
.Y(n_3061)
);

OAI21xp33_ASAP7_75t_L g3062 ( 
.A1(n_2218),
.A2(n_207),
.B(n_208),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2218),
.A2(n_207),
.B(n_208),
.Y(n_3063)
);

AOI21xp5_ASAP7_75t_L g3064 ( 
.A1(n_2218),
.A2(n_208),
.B(n_209),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2200),
.Y(n_3065)
);

OAI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2218),
.A2(n_209),
.B(n_210),
.Y(n_3066)
);

NAND3xp33_ASAP7_75t_L g3067 ( 
.A(n_2424),
.B(n_210),
.C(n_211),
.Y(n_3067)
);

OAI21xp5_ASAP7_75t_L g3068 ( 
.A1(n_2218),
.A2(n_210),
.B(n_211),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2218),
.A2(n_212),
.B(n_213),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2404),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2218),
.B(n_213),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2218),
.B(n_212),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2218),
.B(n_212),
.Y(n_3073)
);

AOI22xp33_ASAP7_75t_L g3074 ( 
.A1(n_2207),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_3074)
);

BUFx8_ASAP7_75t_SL g3075 ( 
.A(n_2258),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2218),
.A2(n_214),
.B(n_216),
.Y(n_3076)
);

OR2x2_ASAP7_75t_L g3077 ( 
.A(n_2218),
.B(n_216),
.Y(n_3077)
);

NOR2xp33_ASAP7_75t_L g3078 ( 
.A(n_2247),
.B(n_217),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2218),
.A2(n_217),
.B(n_218),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2200),
.Y(n_3080)
);

AOI22xp5_ASAP7_75t_L g3081 ( 
.A1(n_2289),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2404),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2218),
.A2(n_218),
.B(n_220),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2218),
.B(n_220),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2218),
.B(n_221),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2200),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2218),
.A2(n_221),
.B(n_222),
.Y(n_3087)
);

INVx1_ASAP7_75t_SL g3088 ( 
.A(n_2244),
.Y(n_3088)
);

BUFx6f_ASAP7_75t_L g3089 ( 
.A(n_2340),
.Y(n_3089)
);

INVx1_ASAP7_75t_SL g3090 ( 
.A(n_2244),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2218),
.B(n_221),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2218),
.A2(n_222),
.B(n_223),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2200),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2218),
.A2(n_222),
.B(n_223),
.Y(n_3094)
);

OAI21x1_ASAP7_75t_L g3095 ( 
.A1(n_2435),
.A2(n_588),
.B(n_587),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2200),
.Y(n_3096)
);

AND2x2_ASAP7_75t_L g3097 ( 
.A(n_2218),
.B(n_223),
.Y(n_3097)
);

AND2x4_ASAP7_75t_L g3098 ( 
.A(n_2200),
.B(n_224),
.Y(n_3098)
);

OAI21xp33_ASAP7_75t_L g3099 ( 
.A1(n_2218),
.A2(n_224),
.B(n_225),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2218),
.B(n_224),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2218),
.B(n_226),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2247),
.B(n_226),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2218),
.B(n_226),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_2218),
.B(n_227),
.Y(n_3104)
);

HB1xp67_ASAP7_75t_L g3105 ( 
.A(n_2244),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2200),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2218),
.B(n_227),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2218),
.A2(n_227),
.B(n_228),
.Y(n_3108)
);

INVx1_ASAP7_75t_SL g3109 ( 
.A(n_2244),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2218),
.A2(n_228),
.B(n_229),
.Y(n_3110)
);

BUFx3_ASAP7_75t_L g3111 ( 
.A(n_2256),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2218),
.B(n_228),
.Y(n_3112)
);

AOI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2218),
.A2(n_229),
.B(n_230),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2200),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2218),
.B(n_229),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2218),
.B(n_230),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2218),
.A2(n_231),
.B(n_232),
.Y(n_3117)
);

BUFx12f_ASAP7_75t_L g3118 ( 
.A(n_2256),
.Y(n_3118)
);

INVxp67_ASAP7_75t_SL g3119 ( 
.A(n_2218),
.Y(n_3119)
);

CKINVDCx5p33_ASAP7_75t_R g3120 ( 
.A(n_2256),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2247),
.B(n_231),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2218),
.B(n_231),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2218),
.B(n_233),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2218),
.A2(n_232),
.B(n_233),
.Y(n_3124)
);

AOI21x1_ASAP7_75t_L g3125 ( 
.A1(n_2435),
.A2(n_233),
.B(n_234),
.Y(n_3125)
);

AOI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2218),
.A2(n_234),
.B(n_235),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2340),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2218),
.B(n_234),
.Y(n_3128)
);

A2O1A1Ixp33_ASAP7_75t_L g3129 ( 
.A1(n_2218),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_2218),
.A2(n_236),
.B(n_237),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2218),
.A2(n_238),
.B(n_239),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2200),
.Y(n_3132)
);

INVx5_ASAP7_75t_L g3133 ( 
.A(n_2340),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2218),
.B(n_238),
.Y(n_3134)
);

AOI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_2218),
.A2(n_239),
.B(n_240),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2404),
.Y(n_3136)
);

AOI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_2218),
.A2(n_240),
.B(n_241),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_2218),
.B(n_242),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2404),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2218),
.B(n_241),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2218),
.A2(n_242),
.B(n_243),
.Y(n_3141)
);

HB1xp67_ASAP7_75t_L g3142 ( 
.A(n_2244),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2200),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2200),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2218),
.B(n_242),
.Y(n_3145)
);

OAI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_2218),
.A2(n_243),
.B(n_244),
.Y(n_3146)
);

AOI21xp5_ASAP7_75t_L g3147 ( 
.A1(n_2218),
.A2(n_243),
.B(n_244),
.Y(n_3147)
);

AND2x2_ASAP7_75t_L g3148 ( 
.A(n_2218),
.B(n_244),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2218),
.B(n_245),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2218),
.B(n_245),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_2218),
.B(n_246),
.Y(n_3151)
);

AOI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_2218),
.A2(n_245),
.B(n_247),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_2218),
.A2(n_247),
.B(n_248),
.Y(n_3153)
);

HB1xp67_ASAP7_75t_L g3154 ( 
.A(n_2244),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_2200),
.B(n_247),
.Y(n_3155)
);

OAI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_2218),
.A2(n_248),
.B(n_249),
.Y(n_3156)
);

O2A1O1Ixp33_ASAP7_75t_L g3157 ( 
.A1(n_2218),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_3157)
);

AOI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_2289),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_3158)
);

OAI22xp5_ASAP7_75t_L g3159 ( 
.A1(n_2218),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_2247),
.B(n_251),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_2218),
.B(n_252),
.Y(n_3161)
);

INVx4_ASAP7_75t_L g3162 ( 
.A(n_2256),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2218),
.A2(n_253),
.B(n_254),
.Y(n_3163)
);

A2O1A1Ixp33_ASAP7_75t_L g3164 ( 
.A1(n_2218),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2200),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2218),
.B(n_253),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2200),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2218),
.B(n_255),
.Y(n_3168)
);

OAI21xp33_ASAP7_75t_L g3169 ( 
.A1(n_2218),
.A2(n_256),
.B(n_257),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2404),
.Y(n_3170)
);

A2O1A1Ixp33_ASAP7_75t_L g3171 ( 
.A1(n_2218),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_3171)
);

AOI21x1_ASAP7_75t_L g3172 ( 
.A1(n_2435),
.A2(n_257),
.B(n_258),
.Y(n_3172)
);

NAND2x1p5_ASAP7_75t_L g3173 ( 
.A(n_2463),
.B(n_259),
.Y(n_3173)
);

BUFx2_ASAP7_75t_L g3174 ( 
.A(n_2244),
.Y(n_3174)
);

AOI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_2218),
.A2(n_259),
.B(n_260),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2218),
.B(n_260),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_2218),
.A2(n_261),
.B(n_262),
.Y(n_3177)
);

O2A1O1Ixp33_ASAP7_75t_L g3178 ( 
.A1(n_2218),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_3178)
);

AOI21xp5_ASAP7_75t_L g3179 ( 
.A1(n_2218),
.A2(n_262),
.B(n_264),
.Y(n_3179)
);

AOI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2218),
.A2(n_264),
.B(n_265),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2218),
.B(n_265),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_SL g3182 ( 
.A(n_2218),
.B(n_266),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2218),
.B(n_265),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2218),
.B(n_266),
.Y(n_3184)
);

A2O1A1Ixp33_ASAP7_75t_L g3185 ( 
.A1(n_2218),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2218),
.B(n_267),
.Y(n_3186)
);

INVx2_ASAP7_75t_SL g3187 ( 
.A(n_2463),
.Y(n_3187)
);

AND2x2_ASAP7_75t_SL g3188 ( 
.A(n_2289),
.B(n_267),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2218),
.A2(n_269),
.B(n_270),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2218),
.A2(n_269),
.B(n_270),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2218),
.B(n_270),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2218),
.B(n_271),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2218),
.A2(n_271),
.B(n_272),
.Y(n_3193)
);

O2A1O1Ixp33_ASAP7_75t_SL g3194 ( 
.A1(n_2218),
.A2(n_274),
.B(n_271),
.C(n_273),
.Y(n_3194)
);

INVx2_ASAP7_75t_SL g3195 ( 
.A(n_2463),
.Y(n_3195)
);

OAI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_2218),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2218),
.B(n_273),
.Y(n_3197)
);

AOI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_2218),
.A2(n_274),
.B(n_275),
.Y(n_3198)
);

AOI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_2218),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_3199)
);

NAND2xp33_ASAP7_75t_L g3200 ( 
.A(n_2340),
.B(n_277),
.Y(n_3200)
);

O2A1O1Ixp33_ASAP7_75t_L g3201 ( 
.A1(n_2218),
.A2(n_279),
.B(n_276),
.C(n_278),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2218),
.B(n_278),
.Y(n_3202)
);

INVxp67_ASAP7_75t_L g3203 ( 
.A(n_2244),
.Y(n_3203)
);

HB1xp67_ASAP7_75t_L g3204 ( 
.A(n_3174),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3059),
.B(n_279),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_3119),
.B(n_279),
.Y(n_3206)
);

NAND2x1p5_ASAP7_75t_L g3207 ( 
.A(n_2977),
.B(n_2976),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_L g3208 ( 
.A(n_2802),
.B(n_280),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_SL g3209 ( 
.A1(n_3188),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3209)
);

A2O1A1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2739),
.A2(n_2781),
.B(n_2784),
.C(n_2691),
.Y(n_3210)
);

OR2x2_ASAP7_75t_L g3211 ( 
.A(n_3088),
.B(n_3090),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_2763),
.A2(n_280),
.B(n_281),
.Y(n_3212)
);

BUFx6f_ASAP7_75t_L g3213 ( 
.A(n_2659),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2647),
.B(n_282),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2891),
.B(n_589),
.Y(n_3215)
);

O2A1O1Ixp33_ASAP7_75t_SL g3216 ( 
.A1(n_2595),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2630),
.A2(n_283),
.B(n_284),
.Y(n_3217)
);

CKINVDCx5p33_ASAP7_75t_R g3218 ( 
.A(n_3118),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3192),
.B(n_283),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_3050),
.B(n_590),
.Y(n_3220)
);

O2A1O1Ixp33_ASAP7_75t_L g3221 ( 
.A1(n_2690),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_2596),
.Y(n_3222)
);

HB1xp67_ASAP7_75t_L g3223 ( 
.A(n_3109),
.Y(n_3223)
);

BUFx3_ASAP7_75t_L g3224 ( 
.A(n_2977),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_2632),
.A2(n_285),
.B(n_286),
.Y(n_3225)
);

OA22x2_ASAP7_75t_L g3226 ( 
.A1(n_2757),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_2659),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2974),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_3058),
.B(n_590),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2975),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3000),
.Y(n_3231)
);

OAI21x1_ASAP7_75t_L g3232 ( 
.A1(n_3095),
.A2(n_288),
.B(n_289),
.Y(n_3232)
);

AOI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_2994),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_3233)
);

A2O1A1Ixp33_ASAP7_75t_L g3234 ( 
.A1(n_3023),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3021),
.Y(n_3235)
);

AOI22xp5_ASAP7_75t_L g3236 ( 
.A1(n_2994),
.A2(n_293),
.B1(n_290),
.B2(n_292),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_2955),
.A2(n_292),
.B(n_293),
.Y(n_3237)
);

OAI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_2592),
.A2(n_292),
.B(n_293),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3007),
.B(n_294),
.Y(n_3239)
);

OAI22xp5_ASAP7_75t_SL g3240 ( 
.A1(n_2704),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3017),
.B(n_294),
.Y(n_3241)
);

AOI22xp5_ASAP7_75t_L g3242 ( 
.A1(n_3009),
.A2(n_3031),
.B1(n_3155),
.B2(n_3098),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3035),
.B(n_295),
.Y(n_3243)
);

INVx5_ASAP7_75t_L g3244 ( 
.A(n_2757),
.Y(n_3244)
);

AND2x2_ASAP7_75t_L g3245 ( 
.A(n_2716),
.B(n_2618),
.Y(n_3245)
);

BUFx2_ASAP7_75t_L g3246 ( 
.A(n_2757),
.Y(n_3246)
);

AND2x2_ASAP7_75t_L g3247 ( 
.A(n_3027),
.B(n_295),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3202),
.A2(n_297),
.B(n_298),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3028),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3048),
.Y(n_3250)
);

OAI21x1_ASAP7_75t_L g3251 ( 
.A1(n_2646),
.A2(n_297),
.B(n_298),
.Y(n_3251)
);

INVx5_ASAP7_75t_L g3252 ( 
.A(n_2664),
.Y(n_3252)
);

NOR3xp33_ASAP7_75t_SL g3253 ( 
.A(n_3120),
.B(n_299),
.C(n_300),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_2956),
.A2(n_299),
.B(n_300),
.Y(n_3254)
);

BUFx3_ASAP7_75t_L g3255 ( 
.A(n_2983),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_3097),
.B(n_299),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_2839),
.B(n_301),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_2795),
.B(n_301),
.Y(n_3258)
);

CKINVDCx20_ASAP7_75t_R g3259 ( 
.A(n_2764),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_3104),
.B(n_302),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3051),
.Y(n_3261)
);

AOI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_3197),
.A2(n_302),
.B(n_303),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_3060),
.Y(n_3263)
);

AOI21xp33_ASAP7_75t_L g3264 ( 
.A1(n_2616),
.A2(n_302),
.B(n_303),
.Y(n_3264)
);

CKINVDCx5p33_ASAP7_75t_R g3265 ( 
.A(n_3075),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_2957),
.A2(n_304),
.B(n_305),
.Y(n_3266)
);

OAI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3009),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_3267)
);

OAI22xp5_ASAP7_75t_L g3268 ( 
.A1(n_3031),
.A2(n_307),
.B1(n_304),
.B2(n_306),
.Y(n_3268)
);

HB1xp67_ASAP7_75t_L g3269 ( 
.A(n_2978),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3061),
.B(n_306),
.Y(n_3270)
);

AOI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_2960),
.A2(n_307),
.B(n_308),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_3111),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3065),
.B(n_307),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3080),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3115),
.B(n_308),
.Y(n_3275)
);

O2A1O1Ixp33_ASAP7_75t_L g3276 ( 
.A1(n_2745),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_3276)
);

AOI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_3191),
.A2(n_309),
.B(n_310),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3086),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3148),
.B(n_309),
.Y(n_3279)
);

NOR2xp67_ASAP7_75t_L g3280 ( 
.A(n_2577),
.B(n_310),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_2965),
.A2(n_312),
.B(n_313),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3093),
.Y(n_3282)
);

BUFx2_ASAP7_75t_L g3283 ( 
.A(n_2675),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_2980),
.A2(n_312),
.B(n_313),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3096),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3161),
.B(n_312),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_2987),
.A2(n_313),
.B(n_314),
.Y(n_3287)
);

A2O1A1Ixp33_ASAP7_75t_L g3288 ( 
.A1(n_3023),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3106),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3114),
.Y(n_3290)
);

OAI22xp5_ASAP7_75t_L g3291 ( 
.A1(n_3098),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_3291)
);

AOI21x1_ASAP7_75t_L g3292 ( 
.A1(n_2738),
.A2(n_315),
.B(n_316),
.Y(n_3292)
);

NAND2x1_ASAP7_75t_L g3293 ( 
.A(n_2951),
.B(n_317),
.Y(n_3293)
);

INVx4_ASAP7_75t_L g3294 ( 
.A(n_2664),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_L g3295 ( 
.A(n_2719),
.B(n_317),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3132),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_2990),
.A2(n_318),
.B(n_319),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3143),
.B(n_318),
.Y(n_3298)
);

BUFx8_ASAP7_75t_L g3299 ( 
.A(n_2709),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_3058),
.B(n_591),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_3001),
.A2(n_318),
.B(n_319),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3155),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3002),
.A2(n_320),
.B(n_321),
.Y(n_3303)
);

NOR2xp33_ASAP7_75t_L g3304 ( 
.A(n_2881),
.B(n_2861),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3144),
.Y(n_3305)
);

OAI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3077),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_SL g3307 ( 
.A(n_3058),
.B(n_591),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_2617),
.B(n_323),
.Y(n_3308)
);

BUFx2_ASAP7_75t_SL g3309 ( 
.A(n_2577),
.Y(n_3309)
);

NAND3xp33_ASAP7_75t_SL g3310 ( 
.A(n_2658),
.B(n_323),
.C(n_325),
.Y(n_3310)
);

A2O1A1Ixp33_ASAP7_75t_SL g3311 ( 
.A1(n_2682),
.A2(n_326),
.B(n_323),
.C(n_325),
.Y(n_3311)
);

A2O1A1Ixp33_ASAP7_75t_L g3312 ( 
.A1(n_2687),
.A2(n_2669),
.B(n_2680),
.C(n_2667),
.Y(n_3312)
);

HB1xp67_ASAP7_75t_L g3313 ( 
.A(n_3045),
.Y(n_3313)
);

NAND2xp33_ASAP7_75t_L g3314 ( 
.A(n_2620),
.B(n_326),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3165),
.Y(n_3315)
);

AOI22xp33_ASAP7_75t_L g3316 ( 
.A1(n_2760),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_3316)
);

O2A1O1Ixp33_ASAP7_75t_L g3317 ( 
.A1(n_2751),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_3317)
);

OAI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_2640),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3006),
.A2(n_329),
.B(n_330),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3167),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_2997),
.Y(n_3321)
);

O2A1O1Ixp33_ASAP7_75t_L g3322 ( 
.A1(n_2749),
.A2(n_333),
.B(n_331),
.C(n_332),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3186),
.A2(n_331),
.B(n_332),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3149),
.B(n_332),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3014),
.A2(n_334),
.B(n_335),
.Y(n_3325)
);

A2O1A1Ixp33_ASAP7_75t_L g3326 ( 
.A1(n_2889),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_3326)
);

AOI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_2605),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_3033),
.A2(n_338),
.B(n_339),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2609),
.B(n_339),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_2619),
.B(n_339),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2621),
.B(n_340),
.Y(n_3331)
);

INVxp67_ASAP7_75t_L g3332 ( 
.A(n_3105),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3011),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2636),
.B(n_340),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2643),
.Y(n_3335)
);

NOR2x1_ASAP7_75t_L g3336 ( 
.A(n_3037),
.B(n_340),
.Y(n_3336)
);

NOR3xp33_ASAP7_75t_L g3337 ( 
.A(n_2588),
.B(n_341),
.C(n_342),
.Y(n_3337)
);

AOI21xp5_ASAP7_75t_L g3338 ( 
.A1(n_3038),
.A2(n_341),
.B(n_342),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_3133),
.B(n_593),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2785),
.B(n_341),
.Y(n_3340)
);

OAI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_2651),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_3341)
);

A2O1A1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_2671),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_3342)
);

INVx2_ASAP7_75t_SL g3343 ( 
.A(n_2750),
.Y(n_3343)
);

AOI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_3041),
.A2(n_343),
.B(n_345),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_3037),
.Y(n_3345)
);

AOI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_3047),
.A2(n_345),
.B(n_346),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2856),
.B(n_346),
.Y(n_3347)
);

BUFx2_ASAP7_75t_L g3348 ( 
.A(n_2662),
.Y(n_3348)
);

NAND3xp33_ASAP7_75t_L g3349 ( 
.A(n_3015),
.B(n_346),
.C(n_347),
.Y(n_3349)
);

O2A1O1Ixp33_ASAP7_75t_SL g3350 ( 
.A1(n_2964),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_3350)
);

OAI22x1_ASAP7_75t_L g3351 ( 
.A1(n_2768),
.A2(n_2831),
.B1(n_3199),
.B2(n_2954),
.Y(n_3351)
);

BUFx2_ASAP7_75t_L g3352 ( 
.A(n_2662),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3049),
.A2(n_347),
.B(n_348),
.Y(n_3353)
);

NAND2x1_ASAP7_75t_L g3354 ( 
.A(n_2951),
.B(n_348),
.Y(n_3354)
);

AOI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_3053),
.A2(n_349),
.B(n_350),
.Y(n_3355)
);

A2O1A1Ixp33_ASAP7_75t_L g3356 ( 
.A1(n_2689),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_3356)
);

A2O1A1Ixp33_ASAP7_75t_L g3357 ( 
.A1(n_2706),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_3357)
);

AND3x1_ASAP7_75t_L g3358 ( 
.A(n_2899),
.B(n_352),
.C(n_354),
.Y(n_3358)
);

OAI21xp33_ASAP7_75t_L g3359 ( 
.A1(n_2623),
.A2(n_354),
.B(n_355),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_L g3360 ( 
.A(n_3203),
.B(n_354),
.Y(n_3360)
);

XNOR2xp5_ASAP7_75t_L g3361 ( 
.A(n_2652),
.B(n_355),
.Y(n_3361)
);

INVx3_ASAP7_75t_L g3362 ( 
.A(n_3162),
.Y(n_3362)
);

BUFx6f_ASAP7_75t_L g3363 ( 
.A(n_2659),
.Y(n_3363)
);

AOI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3054),
.A2(n_356),
.B(n_357),
.Y(n_3364)
);

BUFx3_ASAP7_75t_L g3365 ( 
.A(n_2589),
.Y(n_3365)
);

A2O1A1Ixp33_ASAP7_75t_L g3366 ( 
.A1(n_2650),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_SL g3367 ( 
.A(n_3133),
.B(n_593),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_2741),
.Y(n_3368)
);

NAND3xp33_ASAP7_75t_SL g3369 ( 
.A(n_2932),
.B(n_357),
.C(n_358),
.Y(n_3369)
);

AOI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_2581),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_3370)
);

CKINVDCx6p67_ASAP7_75t_R g3371 ( 
.A(n_3162),
.Y(n_3371)
);

BUFx2_ASAP7_75t_L g3372 ( 
.A(n_2662),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_SL g3373 ( 
.A(n_3133),
.B(n_594),
.Y(n_3373)
);

NOR2xp33_ASAP7_75t_L g3374 ( 
.A(n_2906),
.B(n_359),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_2770),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_3026),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_3040),
.Y(n_3377)
);

HB1xp67_ASAP7_75t_L g3378 ( 
.A(n_3142),
.Y(n_3378)
);

A2O1A1Ixp33_ASAP7_75t_L g3379 ( 
.A1(n_2718),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_3379)
);

INVx1_ASAP7_75t_SL g3380 ( 
.A(n_3154),
.Y(n_3380)
);

CKINVDCx5p33_ASAP7_75t_R g3381 ( 
.A(n_2589),
.Y(n_3381)
);

BUFx3_ASAP7_75t_L g3382 ( 
.A(n_2859),
.Y(n_3382)
);

NAND3xp33_ASAP7_75t_SL g3383 ( 
.A(n_2854),
.B(n_360),
.C(n_362),
.Y(n_3383)
);

OAI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_2651),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_2601),
.B(n_363),
.Y(n_3385)
);

OAI21xp33_ASAP7_75t_L g3386 ( 
.A1(n_2624),
.A2(n_363),
.B(n_364),
.Y(n_3386)
);

CKINVDCx20_ASAP7_75t_R g3387 ( 
.A(n_2679),
.Y(n_3387)
);

OR2x6_ASAP7_75t_L g3388 ( 
.A(n_2664),
.B(n_365),
.Y(n_3388)
);

OAI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_2954),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_3389)
);

OAI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3199),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_3390)
);

BUFx2_ASAP7_75t_L g3391 ( 
.A(n_2662),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3056),
.A2(n_366),
.B(n_368),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3070),
.Y(n_3393)
);

OAI22xp5_ASAP7_75t_L g3394 ( 
.A1(n_3072),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_2604),
.B(n_369),
.Y(n_3395)
);

AOI33xp33_ASAP7_75t_L g3396 ( 
.A1(n_2593),
.A2(n_372),
.A3(n_374),
.B1(n_370),
.B2(n_371),
.B3(n_373),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_R g3397 ( 
.A(n_2776),
.B(n_2801),
.Y(n_3397)
);

A2O1A1Ixp33_ASAP7_75t_L g3398 ( 
.A1(n_2615),
.A2(n_372),
.B(n_370),
.C(n_371),
.Y(n_3398)
);

AND2x2_ASAP7_75t_SL g3399 ( 
.A(n_2826),
.B(n_371),
.Y(n_3399)
);

OAI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3073),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3400)
);

CKINVDCx5p33_ASAP7_75t_R g3401 ( 
.A(n_3039),
.Y(n_3401)
);

BUFx2_ASAP7_75t_L g3402 ( 
.A(n_2723),
.Y(n_3402)
);

OAI22x1_ASAP7_75t_L g3403 ( 
.A1(n_3173),
.A2(n_2627),
.B1(n_3013),
.B2(n_2854),
.Y(n_3403)
);

INVx3_ASAP7_75t_L g3404 ( 
.A(n_2915),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2782),
.Y(n_3405)
);

INVx4_ASAP7_75t_L g3406 ( 
.A(n_2848),
.Y(n_3406)
);

INVx3_ASAP7_75t_SL g3407 ( 
.A(n_2848),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_2603),
.B(n_374),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3084),
.A2(n_375),
.B(n_376),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_2600),
.B(n_375),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_2903),
.B(n_376),
.Y(n_3411)
);

OA22x2_ASAP7_75t_L g3412 ( 
.A1(n_2660),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3085),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_3091),
.A2(n_379),
.B(n_380),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3082),
.Y(n_3415)
);

NOR3xp33_ASAP7_75t_L g3416 ( 
.A(n_2722),
.B(n_380),
.C(n_381),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_3100),
.A2(n_380),
.B(n_382),
.Y(n_3417)
);

OAI21x1_ASAP7_75t_L g3418 ( 
.A1(n_2648),
.A2(n_382),
.B(n_383),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3101),
.B(n_382),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2771),
.Y(n_3420)
);

A2O1A1Ixp33_ASAP7_75t_L g3421 ( 
.A1(n_2674),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_3136),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3032),
.Y(n_3423)
);

BUFx3_ASAP7_75t_L g3424 ( 
.A(n_2848),
.Y(n_3424)
);

AOI21xp5_ASAP7_75t_L g3425 ( 
.A1(n_3103),
.A2(n_383),
.B(n_384),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_SL g3426 ( 
.A(n_2877),
.B(n_594),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_2843),
.B(n_385),
.Y(n_3427)
);

A2O1A1Ixp33_ASAP7_75t_L g3428 ( 
.A1(n_2840),
.A2(n_387),
.B(n_385),
.C(n_386),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_2877),
.B(n_595),
.Y(n_3429)
);

INVxp67_ASAP7_75t_SL g3430 ( 
.A(n_2863),
.Y(n_3430)
);

OAI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_2614),
.A2(n_386),
.B(n_387),
.Y(n_3431)
);

BUFx5_ASAP7_75t_L g3432 ( 
.A(n_2620),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_2666),
.Y(n_3433)
);

OAI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3107),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_3434)
);

AOI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_3112),
.A2(n_388),
.B(n_389),
.Y(n_3435)
);

OR2x2_ASAP7_75t_L g3436 ( 
.A(n_2574),
.B(n_390),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_2582),
.B(n_390),
.Y(n_3437)
);

OAI22xp5_ASAP7_75t_L g3438 ( 
.A1(n_3116),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_3438)
);

AOI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_3122),
.A2(n_391),
.B(n_392),
.Y(n_3439)
);

AO21x1_ASAP7_75t_L g3440 ( 
.A1(n_2966),
.A2(n_3004),
.B(n_2972),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_2731),
.B(n_391),
.Y(n_3441)
);

AND2x4_ASAP7_75t_L g3442 ( 
.A(n_2582),
.B(n_393),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_2701),
.B(n_2673),
.Y(n_3443)
);

OR2x6_ASAP7_75t_SL g3444 ( 
.A(n_2754),
.B(n_393),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_2668),
.B(n_394),
.Y(n_3445)
);

AOI22xp33_ASAP7_75t_L g3446 ( 
.A1(n_2953),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3446)
);

OAI22x1_ASAP7_75t_L g3447 ( 
.A1(n_2971),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3447)
);

OAI22x1_ASAP7_75t_L g3448 ( 
.A1(n_2992),
.A2(n_3081),
.B1(n_3158),
.B2(n_2668),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3128),
.B(n_395),
.Y(n_3449)
);

OAI22xp5_ASAP7_75t_L g3450 ( 
.A1(n_3134),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_3450)
);

AOI21x1_ASAP7_75t_L g3451 ( 
.A1(n_2738),
.A2(n_397),
.B(n_398),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_2877),
.B(n_596),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3140),
.B(n_398),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_L g3454 ( 
.A(n_2847),
.B(n_399),
.Y(n_3454)
);

NAND3xp33_ASAP7_75t_L g3455 ( 
.A(n_3074),
.B(n_400),
.C(n_401),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_SL g3456 ( 
.A(n_2912),
.B(n_400),
.Y(n_3456)
);

INVx4_ASAP7_75t_L g3457 ( 
.A(n_2893),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3145),
.B(n_400),
.Y(n_3458)
);

A2O1A1Ixp33_ASAP7_75t_SL g3459 ( 
.A1(n_2860),
.A2(n_403),
.B(n_401),
.C(n_402),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3139),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_L g3461 ( 
.A(n_2670),
.B(n_2622),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2715),
.Y(n_3462)
);

O2A1O1Ixp5_ASAP7_75t_SL g3463 ( 
.A1(n_2639),
.A2(n_597),
.B(n_598),
.C(n_596),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_SL g3464 ( 
.A(n_2863),
.B(n_2634),
.Y(n_3464)
);

NOR3xp33_ASAP7_75t_SL g3465 ( 
.A(n_2918),
.B(n_401),
.C(n_402),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3150),
.B(n_402),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_2774),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3166),
.B(n_3168),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_SL g3469 ( 
.A(n_2915),
.B(n_2893),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_2620),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3176),
.A2(n_403),
.B(n_404),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3181),
.A2(n_404),
.B(n_405),
.Y(n_3472)
);

INVxp67_ASAP7_75t_L g3473 ( 
.A(n_2962),
.Y(n_3473)
);

BUFx6f_ASAP7_75t_L g3474 ( 
.A(n_2695),
.Y(n_3474)
);

BUFx4f_ASAP7_75t_L g3475 ( 
.A(n_2893),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_3183),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_2654),
.B(n_407),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3184),
.B(n_407),
.Y(n_3478)
);

A2O1A1Ixp33_ASAP7_75t_L g3479 ( 
.A1(n_2726),
.A2(n_410),
.B(n_408),
.C(n_409),
.Y(n_3479)
);

INVx1_ASAP7_75t_SL g3480 ( 
.A(n_2874),
.Y(n_3480)
);

AOI21x1_ASAP7_75t_L g3481 ( 
.A1(n_2698),
.A2(n_2573),
.B(n_2958),
.Y(n_3481)
);

BUFx12f_ASAP7_75t_L g3482 ( 
.A(n_2811),
.Y(n_3482)
);

A2O1A1Ixp33_ASAP7_75t_L g3483 ( 
.A1(n_2852),
.A2(n_410),
.B(n_408),
.C(n_409),
.Y(n_3483)
);

INVx4_ASAP7_75t_L g3484 ( 
.A(n_2893),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_2924),
.B(n_409),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_2644),
.A2(n_410),
.B(n_411),
.Y(n_3486)
);

BUFx2_ASAP7_75t_L g3487 ( 
.A(n_2620),
.Y(n_3487)
);

CKINVDCx5p33_ASAP7_75t_R g3488 ( 
.A(n_2882),
.Y(n_3488)
);

OAI22x1_ASAP7_75t_L g3489 ( 
.A1(n_2710),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2752),
.B(n_411),
.Y(n_3490)
);

AOI21xp5_ASAP7_75t_L g3491 ( 
.A1(n_2767),
.A2(n_412),
.B(n_413),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_2683),
.B(n_412),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_2688),
.B(n_413),
.Y(n_3493)
);

AND2x4_ASAP7_75t_L g3494 ( 
.A(n_2917),
.B(n_414),
.Y(n_3494)
);

AOI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_2657),
.A2(n_414),
.B(n_415),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_L g3496 ( 
.A(n_2613),
.B(n_414),
.Y(n_3496)
);

CKINVDCx5p33_ASAP7_75t_R g3497 ( 
.A(n_2882),
.Y(n_3497)
);

INVx4_ASAP7_75t_L g3498 ( 
.A(n_2816),
.Y(n_3498)
);

BUFx6f_ASAP7_75t_L g3499 ( 
.A(n_2695),
.Y(n_3499)
);

O2A1O1Ixp33_ASAP7_75t_L g3500 ( 
.A1(n_2800),
.A2(n_2794),
.B(n_2887),
.C(n_2773),
.Y(n_3500)
);

CKINVDCx5p33_ASAP7_75t_R g3501 ( 
.A(n_3187),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_2809),
.Y(n_3502)
);

BUFx2_ASAP7_75t_L g3503 ( 
.A(n_3195),
.Y(n_3503)
);

A2O1A1Ixp33_ASAP7_75t_L g3504 ( 
.A1(n_2742),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_3504)
);

O2A1O1Ixp33_ASAP7_75t_L g3505 ( 
.A1(n_2823),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_2575),
.B(n_417),
.Y(n_3506)
);

O2A1O1Ixp33_ASAP7_75t_L g3507 ( 
.A1(n_2894),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_3507)
);

BUFx2_ASAP7_75t_L g3508 ( 
.A(n_2814),
.Y(n_3508)
);

O2A1O1Ixp33_ASAP7_75t_L g3509 ( 
.A1(n_2797),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_3509)
);

INVx2_ASAP7_75t_SL g3510 ( 
.A(n_2874),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3170),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_2663),
.A2(n_419),
.B(n_420),
.Y(n_3512)
);

O2A1O1Ixp33_ASAP7_75t_L g3513 ( 
.A1(n_2875),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_2871),
.B(n_423),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_2890),
.B(n_2865),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_2676),
.A2(n_423),
.B(n_424),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_2677),
.A2(n_2678),
.B(n_2692),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_2733),
.B(n_424),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_2857),
.B(n_424),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_2970),
.B(n_2981),
.Y(n_3520)
);

NOR3xp33_ASAP7_75t_L g3521 ( 
.A(n_2724),
.B(n_425),
.C(n_426),
.Y(n_3521)
);

AOI21xp5_ASAP7_75t_L g3522 ( 
.A1(n_2693),
.A2(n_2700),
.B(n_2694),
.Y(n_3522)
);

AOI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_2653),
.A2(n_425),
.B(n_426),
.Y(n_3523)
);

OAI21xp33_ASAP7_75t_L g3524 ( 
.A1(n_2655),
.A2(n_427),
.B(n_428),
.Y(n_3524)
);

OAI21xp33_ASAP7_75t_L g3525 ( 
.A1(n_3055),
.A2(n_427),
.B(n_428),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_2995),
.A2(n_3030),
.B1(n_3034),
.B2(n_3016),
.Y(n_3526)
);

OAI221xp5_ASAP7_75t_L g3527 ( 
.A1(n_3078),
.A2(n_3102),
.B1(n_3160),
.B2(n_3121),
.C(n_2649),
.Y(n_3527)
);

OAI22xp5_ASAP7_75t_L g3528 ( 
.A1(n_2634),
.A2(n_430),
.B1(n_427),
.B2(n_429),
.Y(n_3528)
);

HB1xp67_ASAP7_75t_L g3529 ( 
.A(n_2880),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_2576),
.B(n_429),
.Y(n_3530)
);

INVx4_ASAP7_75t_L g3531 ( 
.A(n_2816),
.Y(n_3531)
);

INVx2_ASAP7_75t_SL g3532 ( 
.A(n_2816),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_SL g3533 ( 
.A(n_2591),
.B(n_599),
.Y(n_3533)
);

AND2x4_ASAP7_75t_L g3534 ( 
.A(n_2917),
.B(n_429),
.Y(n_3534)
);

O2A1O1Ixp33_ASAP7_75t_L g3535 ( 
.A1(n_2611),
.A2(n_432),
.B(n_430),
.C(n_431),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_2813),
.Y(n_3536)
);

CKINVDCx5p33_ASAP7_75t_R g3537 ( 
.A(n_2862),
.Y(n_3537)
);

BUFx8_ASAP7_75t_L g3538 ( 
.A(n_2938),
.Y(n_3538)
);

BUFx6f_ASAP7_75t_L g3539 ( 
.A(n_2695),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_2579),
.B(n_431),
.Y(n_3540)
);

AO21x2_ASAP7_75t_L g3541 ( 
.A1(n_2599),
.A2(n_432),
.B(n_433),
.Y(n_3541)
);

OAI21xp33_ASAP7_75t_L g3542 ( 
.A1(n_3062),
.A2(n_432),
.B(n_433),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_2656),
.Y(n_3543)
);

A2O1A1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_3029),
.A2(n_435),
.B(n_433),
.C(n_434),
.Y(n_3544)
);

CKINVDCx20_ASAP7_75t_R g3545 ( 
.A(n_2808),
.Y(n_3545)
);

AOI22xp33_ASAP7_75t_L g3546 ( 
.A1(n_2661),
.A2(n_437),
.B1(n_434),
.B2(n_436),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_2580),
.B(n_434),
.Y(n_3547)
);

BUFx12f_ASAP7_75t_L g3548 ( 
.A(n_2914),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_L g3549 ( 
.A(n_2578),
.B(n_436),
.Y(n_3549)
);

A2O1A1Ixp33_ASAP7_75t_SL g3550 ( 
.A1(n_2883),
.A2(n_438),
.B(n_436),
.C(n_437),
.Y(n_3550)
);

BUFx6f_ASAP7_75t_L g3551 ( 
.A(n_2713),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_2830),
.Y(n_3552)
);

AOI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_2642),
.A2(n_2707),
.B(n_2790),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_2729),
.Y(n_3554)
);

BUFx2_ASAP7_75t_L g3555 ( 
.A(n_2585),
.Y(n_3555)
);

AND2x4_ASAP7_75t_L g3556 ( 
.A(n_2886),
.B(n_437),
.Y(n_3556)
);

BUFx3_ASAP7_75t_L g3557 ( 
.A(n_2907),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_2951),
.B(n_2961),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_2792),
.A2(n_439),
.B(n_440),
.Y(n_3559)
);

BUFx2_ASAP7_75t_SL g3560 ( 
.A(n_2880),
.Y(n_3560)
);

BUFx3_ASAP7_75t_L g3561 ( 
.A(n_2717),
.Y(n_3561)
);

OAI21x1_ASAP7_75t_SL g3562 ( 
.A1(n_2845),
.A2(n_439),
.B(n_440),
.Y(n_3562)
);

BUFx3_ASAP7_75t_L g3563 ( 
.A(n_2717),
.Y(n_3563)
);

O2A1O1Ixp33_ASAP7_75t_L g3564 ( 
.A1(n_2873),
.A2(n_442),
.B(n_439),
.C(n_441),
.Y(n_3564)
);

A2O1A1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_3043),
.A2(n_444),
.B(n_442),
.C(n_443),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_2753),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_2584),
.B(n_442),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_SL g3568 ( 
.A(n_2961),
.B(n_599),
.Y(n_3568)
);

AO21x1_ASAP7_75t_L g3569 ( 
.A1(n_3057),
.A2(n_602),
.B(n_601),
.Y(n_3569)
);

BUFx2_ASAP7_75t_L g3570 ( 
.A(n_2901),
.Y(n_3570)
);

CKINVDCx20_ASAP7_75t_R g3571 ( 
.A(n_2812),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_L g3572 ( 
.A1(n_3018),
.A2(n_443),
.B(n_444),
.Y(n_3572)
);

AOI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_2672),
.A2(n_2728),
.B1(n_2778),
.B2(n_2807),
.Y(n_3573)
);

AOI22xp5_ASAP7_75t_L g3574 ( 
.A1(n_2587),
.A2(n_446),
.B1(n_443),
.B2(n_445),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_2713),
.A2(n_445),
.B(n_447),
.Y(n_3575)
);

HB1xp67_ASAP7_75t_L g3576 ( 
.A(n_2901),
.Y(n_3576)
);

INVx1_ASAP7_75t_SL g3577 ( 
.A(n_2798),
.Y(n_3577)
);

BUFx6f_ASAP7_75t_L g3578 ( 
.A(n_2713),
.Y(n_3578)
);

INVx5_ASAP7_75t_L g3579 ( 
.A(n_2961),
.Y(n_3579)
);

INVx3_ASAP7_75t_L g3580 ( 
.A(n_2789),
.Y(n_3580)
);

INVx5_ASAP7_75t_L g3581 ( 
.A(n_3089),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_SL g3582 ( 
.A1(n_3066),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_2736),
.A2(n_448),
.B(n_449),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_2583),
.B(n_448),
.Y(n_3584)
);

NOR3xp33_ASAP7_75t_SL g3585 ( 
.A(n_2923),
.B(n_449),
.C(n_450),
.Y(n_3585)
);

AOI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_2736),
.A2(n_449),
.B(n_450),
.Y(n_3586)
);

INVx1_ASAP7_75t_SL g3587 ( 
.A(n_2928),
.Y(n_3587)
);

OAI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_2590),
.A2(n_451),
.B(n_452),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_2758),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_2685),
.Y(n_3590)
);

INVx3_ASAP7_75t_L g3591 ( 
.A(n_2789),
.Y(n_3591)
);

OAI22xp5_ASAP7_75t_L g3592 ( 
.A1(n_2712),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_3592)
);

OAI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_2921),
.A2(n_451),
.B(n_452),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_2895),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_2586),
.B(n_2597),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_2789),
.Y(n_3596)
);

INVxp67_ASAP7_75t_L g3597 ( 
.A(n_2740),
.Y(n_3597)
);

A2O1A1Ixp33_ASAP7_75t_L g3598 ( 
.A1(n_3068),
.A2(n_456),
.B(n_454),
.C(n_455),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_2606),
.B(n_454),
.Y(n_3599)
);

NOR2xp33_ASAP7_75t_L g3600 ( 
.A(n_2607),
.B(n_456),
.Y(n_3600)
);

INVx3_ASAP7_75t_L g3601 ( 
.A(n_3089),
.Y(n_3601)
);

INVx6_ASAP7_75t_L g3602 ( 
.A(n_2878),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_2897),
.B(n_2759),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_2866),
.B(n_456),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2736),
.A2(n_457),
.B(n_458),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_SL g3606 ( 
.A(n_3089),
.B(n_601),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_2772),
.A2(n_457),
.B(n_458),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_2772),
.A2(n_457),
.B(n_458),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_2772),
.A2(n_459),
.B(n_460),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_2777),
.A2(n_2844),
.B(n_2936),
.Y(n_3610)
);

AND2x4_ASAP7_75t_L g3611 ( 
.A(n_2908),
.B(n_459),
.Y(n_3611)
);

NOR3xp33_ASAP7_75t_L g3612 ( 
.A(n_2748),
.B(n_459),
.C(n_460),
.Y(n_3612)
);

AOI222xp33_ASAP7_75t_L g3613 ( 
.A1(n_2696),
.A2(n_462),
.B1(n_464),
.B2(n_460),
.C1(n_461),
.C2(n_463),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2702),
.Y(n_3614)
);

CKINVDCx20_ASAP7_75t_R g3615 ( 
.A(n_2869),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_L g3616 ( 
.A1(n_3125),
.A2(n_461),
.B(n_462),
.Y(n_3616)
);

INVx4_ASAP7_75t_L g3617 ( 
.A(n_3127),
.Y(n_3617)
);

O2A1O1Ixp33_ASAP7_75t_L g3618 ( 
.A1(n_2935),
.A2(n_463),
.B(n_461),
.C(n_462),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_3127),
.B(n_602),
.Y(n_3619)
);

AOI22xp5_ASAP7_75t_L g3620 ( 
.A1(n_2931),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_3620)
);

NOR2xp67_ASAP7_75t_L g3621 ( 
.A(n_2945),
.B(n_464),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_2708),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2777),
.A2(n_466),
.B(n_467),
.Y(n_3623)
);

BUFx6f_ASAP7_75t_L g3624 ( 
.A(n_2777),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_2711),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_2950),
.A2(n_466),
.B(n_467),
.Y(n_3626)
);

O2A1O1Ixp33_ASAP7_75t_L g3627 ( 
.A1(n_2732),
.A2(n_468),
.B(n_466),
.C(n_467),
.Y(n_3627)
);

AOI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_2968),
.A2(n_468),
.B(n_469),
.Y(n_3628)
);

INVx3_ASAP7_75t_L g3629 ( 
.A(n_2612),
.Y(n_3629)
);

O2A1O1Ixp33_ASAP7_75t_L g3630 ( 
.A1(n_2761),
.A2(n_471),
.B(n_469),
.C(n_470),
.Y(n_3630)
);

AOI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_2933),
.A2(n_473),
.B1(n_470),
.B2(n_471),
.Y(n_3631)
);

CKINVDCx20_ASAP7_75t_R g3632 ( 
.A(n_2842),
.Y(n_3632)
);

INVx1_ASAP7_75t_SL g3633 ( 
.A(n_2878),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_2765),
.B(n_470),
.Y(n_3634)
);

OR2x6_ASAP7_75t_L g3635 ( 
.A(n_2705),
.B(n_471),
.Y(n_3635)
);

AND2x4_ASAP7_75t_L g3636 ( 
.A(n_2939),
.B(n_473),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_2743),
.B(n_473),
.Y(n_3637)
);

NOR3xp33_ASAP7_75t_SL g3638 ( 
.A(n_2686),
.B(n_474),
.C(n_475),
.Y(n_3638)
);

O2A1O1Ixp33_ASAP7_75t_L g3639 ( 
.A1(n_2986),
.A2(n_476),
.B(n_474),
.C(n_475),
.Y(n_3639)
);

OAI22xp5_ASAP7_75t_L g3640 ( 
.A1(n_3067),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_3640)
);

OAI21xp33_ASAP7_75t_L g3641 ( 
.A1(n_3099),
.A2(n_476),
.B(n_477),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_2625),
.B(n_477),
.Y(n_3642)
);

OAI21xp33_ASAP7_75t_L g3643 ( 
.A1(n_3169),
.A2(n_478),
.B(n_479),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_SL g3644 ( 
.A(n_3127),
.B(n_603),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_2626),
.B(n_478),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_SL g3646 ( 
.A(n_2714),
.B(n_603),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_2746),
.Y(n_3647)
);

AND2x4_ASAP7_75t_L g3648 ( 
.A(n_2783),
.B(n_479),
.Y(n_3648)
);

AOI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3172),
.A2(n_479),
.B(n_480),
.Y(n_3649)
);

NOR2xp33_ASAP7_75t_L g3650 ( 
.A(n_2943),
.B(n_480),
.Y(n_3650)
);

OAI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_2598),
.A2(n_480),
.B(n_481),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_2779),
.B(n_481),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_2594),
.B(n_481),
.Y(n_3653)
);

AOI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_2989),
.A2(n_482),
.B(n_483),
.Y(n_3654)
);

AOI21x1_ASAP7_75t_L g3655 ( 
.A1(n_2635),
.A2(n_482),
.B(n_483),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_2949),
.B(n_482),
.Y(n_3656)
);

NOR2xp33_ASAP7_75t_L g3657 ( 
.A(n_2920),
.B(n_484),
.Y(n_3657)
);

HB1xp67_ASAP7_75t_L g3658 ( 
.A(n_2799),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_2993),
.A2(n_3010),
.B(n_2996),
.Y(n_3659)
);

NAND2x1_ASAP7_75t_L g3660 ( 
.A(n_2612),
.B(n_484),
.Y(n_3660)
);

HB1xp67_ASAP7_75t_L g3661 ( 
.A(n_2805),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3146),
.A2(n_3156),
.B(n_2714),
.C(n_2780),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_2937),
.Y(n_3663)
);

BUFx3_ASAP7_75t_L g3664 ( 
.A(n_2645),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_2841),
.B(n_484),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_2796),
.B(n_485),
.Y(n_3666)
);

O2A1O1Ixp33_ASAP7_75t_L g3667 ( 
.A1(n_3012),
.A2(n_3071),
.B(n_3138),
.C(n_3123),
.Y(n_3667)
);

INVx4_ASAP7_75t_SL g3668 ( 
.A(n_2878),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_2937),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_2629),
.Y(n_3670)
);

INVx3_ASAP7_75t_L g3671 ( 
.A(n_2645),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3151),
.A2(n_486),
.B(n_487),
.Y(n_3672)
);

O2A1O1Ixp33_ASAP7_75t_L g3673 ( 
.A1(n_3182),
.A2(n_2638),
.B(n_2896),
.C(n_2867),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_2641),
.A2(n_486),
.B(n_487),
.Y(n_3674)
);

INVx1_ASAP7_75t_SL g3675 ( 
.A(n_2885),
.Y(n_3675)
);

AND2x4_ASAP7_75t_L g3676 ( 
.A(n_2783),
.B(n_486),
.Y(n_3676)
);

OAI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_2631),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_2608),
.B(n_488),
.Y(n_3678)
);

NOR3xp33_ASAP7_75t_L g3679 ( 
.A(n_2821),
.B(n_489),
.C(n_490),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_2610),
.B(n_489),
.Y(n_3680)
);

BUFx6f_ASAP7_75t_L g3681 ( 
.A(n_2885),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3200),
.A2(n_490),
.B(n_491),
.Y(n_3682)
);

O2A1O1Ixp33_ASAP7_75t_L g3683 ( 
.A1(n_2735),
.A2(n_3129),
.B(n_3171),
.C(n_3164),
.Y(n_3683)
);

INVx11_ASAP7_75t_L g3684 ( 
.A(n_2942),
.Y(n_3684)
);

CKINVDCx6p67_ASAP7_75t_R g3685 ( 
.A(n_2885),
.Y(n_3685)
);

OAI22xp5_ASAP7_75t_L g3686 ( 
.A1(n_2766),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_3686)
);

AOI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_2913),
.A2(n_491),
.B(n_492),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_2633),
.B(n_492),
.Y(n_3688)
);

BUFx2_ASAP7_75t_L g3689 ( 
.A(n_2681),
.Y(n_3689)
);

INVx1_ASAP7_75t_SL g3690 ( 
.A(n_2681),
.Y(n_3690)
);

O2A1O1Ixp33_ASAP7_75t_SL g3691 ( 
.A1(n_2747),
.A2(n_495),
.B(n_493),
.C(n_494),
.Y(n_3691)
);

INVx5_ASAP7_75t_L g3692 ( 
.A(n_2835),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_2806),
.B(n_493),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_2855),
.B(n_2628),
.Y(n_3694)
);

INVx4_ASAP7_75t_L g3695 ( 
.A(n_2835),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_2825),
.A2(n_494),
.B(n_495),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_2665),
.Y(n_3697)
);

OAI22xp5_ASAP7_75t_L g3698 ( 
.A1(n_2853),
.A2(n_2909),
.B1(n_2888),
.B2(n_3185),
.Y(n_3698)
);

AND3x1_ASAP7_75t_SL g3699 ( 
.A(n_2904),
.B(n_495),
.C(n_496),
.Y(n_3699)
);

AOI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_2637),
.A2(n_496),
.B(n_497),
.Y(n_3700)
);

O2A1O1Ixp33_ASAP7_75t_L g3701 ( 
.A1(n_2941),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_2959),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_2810),
.B(n_498),
.Y(n_3703)
);

A2O1A1Ixp33_ASAP7_75t_L g3704 ( 
.A1(n_2804),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_3704)
);

INVx3_ASAP7_75t_L g3705 ( 
.A(n_2945),
.Y(n_3705)
);

INVx3_ASAP7_75t_L g3706 ( 
.A(n_2898),
.Y(n_3706)
);

NOR2xp33_ASAP7_75t_L g3707 ( 
.A(n_2898),
.B(n_500),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_2870),
.A2(n_501),
.B(n_502),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_2911),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3024),
.Y(n_3710)
);

BUFx4f_ASAP7_75t_L g3711 ( 
.A(n_2884),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3194),
.A2(n_502),
.B(n_503),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_2926),
.B(n_502),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_2697),
.B(n_2699),
.Y(n_3714)
);

NAND3xp33_ASAP7_75t_SL g3715 ( 
.A(n_2910),
.B(n_503),
.C(n_504),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3025),
.Y(n_3716)
);

INVx3_ASAP7_75t_L g3717 ( 
.A(n_2602),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_2703),
.B(n_504),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3159),
.B(n_504),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_2868),
.B(n_505),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_2979),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3008),
.Y(n_3722)
);

NAND2x1p5_ASAP7_75t_L g3723 ( 
.A(n_2829),
.B(n_505),
.Y(n_3723)
);

AOI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_2725),
.A2(n_505),
.B(n_506),
.Y(n_3724)
);

OAI21xp33_ASAP7_75t_SL g3725 ( 
.A1(n_2836),
.A2(n_2948),
.B(n_3196),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_2919),
.B(n_506),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_2730),
.B(n_506),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_SL g3728 ( 
.A(n_2846),
.B(n_604),
.Y(n_3728)
);

A2O1A1Ixp33_ASAP7_75t_SL g3729 ( 
.A1(n_2982),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_2940),
.Y(n_3730)
);

BUFx8_ASAP7_75t_L g3731 ( 
.A(n_2922),
.Y(n_3731)
);

O2A1O1Ixp33_ASAP7_75t_L g3732 ( 
.A1(n_2769),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_2727),
.B(n_2947),
.Y(n_3733)
);

AOI21x1_ASAP7_75t_L g3734 ( 
.A1(n_2791),
.A2(n_509),
.B(n_510),
.Y(n_3734)
);

OAI21xp33_ASAP7_75t_L g3735 ( 
.A1(n_2925),
.A2(n_510),
.B(n_511),
.Y(n_3735)
);

INVxp67_ASAP7_75t_SL g3736 ( 
.A(n_2985),
.Y(n_3736)
);

OAI21x1_ASAP7_75t_L g3737 ( 
.A1(n_3481),
.A2(n_2755),
.B(n_2744),
.Y(n_3737)
);

AO31x2_ASAP7_75t_L g3738 ( 
.A1(n_3210),
.A2(n_2737),
.A3(n_2721),
.B(n_2879),
.Y(n_3738)
);

INVx3_ASAP7_75t_L g3739 ( 
.A(n_3294),
.Y(n_3739)
);

BUFx2_ASAP7_75t_L g3740 ( 
.A(n_3545),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3610),
.A2(n_2762),
.B(n_2756),
.Y(n_3741)
);

NOR2x1_ASAP7_75t_SL g3742 ( 
.A(n_3457),
.B(n_3484),
.Y(n_3742)
);

HB1xp67_ASAP7_75t_L g3743 ( 
.A(n_3211),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3420),
.B(n_3304),
.Y(n_3744)
);

AND2x6_ASAP7_75t_L g3745 ( 
.A(n_3242),
.B(n_2988),
.Y(n_3745)
);

AOI21x1_ASAP7_75t_L g3746 ( 
.A1(n_3470),
.A2(n_2815),
.B(n_2832),
.Y(n_3746)
);

AOI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3517),
.A2(n_3157),
.B(n_3003),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_3218),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3522),
.A2(n_3201),
.B(n_3178),
.Y(n_3749)
);

AO31x2_ASAP7_75t_L g3750 ( 
.A1(n_3440),
.A2(n_2833),
.A3(n_2819),
.B(n_2822),
.Y(n_3750)
);

OAI21x1_ASAP7_75t_L g3751 ( 
.A1(n_3709),
.A2(n_2824),
.B(n_2820),
.Y(n_3751)
);

OAI21x1_ASAP7_75t_L g3752 ( 
.A1(n_3558),
.A2(n_2827),
.B(n_2834),
.Y(n_3752)
);

AOI21xp5_ASAP7_75t_L g3753 ( 
.A1(n_3553),
.A2(n_2838),
.B(n_2793),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3230),
.Y(n_3754)
);

A2O1A1Ixp33_ASAP7_75t_L g3755 ( 
.A1(n_3475),
.A2(n_3314),
.B(n_3500),
.C(n_3588),
.Y(n_3755)
);

HB1xp67_ASAP7_75t_L g3756 ( 
.A(n_3223),
.Y(n_3756)
);

AND2x4_ASAP7_75t_L g3757 ( 
.A(n_3252),
.B(n_2905),
.Y(n_3757)
);

BUFx10_ASAP7_75t_L g3758 ( 
.A(n_3343),
.Y(n_3758)
);

HB1xp67_ASAP7_75t_L g3759 ( 
.A(n_3204),
.Y(n_3759)
);

NAND3xp33_ASAP7_75t_L g3760 ( 
.A(n_3253),
.B(n_2803),
.C(n_2952),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3222),
.Y(n_3761)
);

OAI21x1_ASAP7_75t_L g3762 ( 
.A1(n_3232),
.A2(n_2837),
.B(n_2720),
.Y(n_3762)
);

O2A1O1Ixp33_ASAP7_75t_SL g3763 ( 
.A1(n_3215),
.A2(n_2892),
.B(n_2967),
.C(n_2963),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3228),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3312),
.A2(n_2788),
.B(n_2684),
.Y(n_3765)
);

OAI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3457),
.A2(n_2734),
.B1(n_2973),
.B2(n_2969),
.Y(n_3766)
);

AOI21xp33_ASAP7_75t_L g3767 ( 
.A1(n_3725),
.A2(n_2916),
.B(n_2984),
.Y(n_3767)
);

BUFx6f_ASAP7_75t_L g3768 ( 
.A(n_3252),
.Y(n_3768)
);

NAND3xp33_ASAP7_75t_L g3769 ( 
.A(n_3526),
.B(n_2998),
.C(n_2991),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3714),
.A2(n_3005),
.B(n_2999),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3245),
.B(n_510),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3662),
.A2(n_3698),
.B(n_3468),
.Y(n_3772)
);

OA22x2_ASAP7_75t_L g3773 ( 
.A1(n_3388),
.A2(n_3020),
.B1(n_3022),
.B2(n_3019),
.Y(n_3773)
);

AOI21x1_ASAP7_75t_L g3774 ( 
.A1(n_3487),
.A2(n_2872),
.B(n_2864),
.Y(n_3774)
);

BUFx10_ASAP7_75t_L g3775 ( 
.A(n_3381),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3235),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3250),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3423),
.B(n_2858),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3659),
.A2(n_3042),
.B(n_3036),
.Y(n_3779)
);

BUFx10_ASAP7_75t_L g3780 ( 
.A(n_3388),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3274),
.Y(n_3781)
);

OAI22xp33_ASAP7_75t_L g3782 ( 
.A1(n_3456),
.A2(n_3046),
.B1(n_3052),
.B2(n_3044),
.Y(n_3782)
);

BUFx12f_ASAP7_75t_L g3783 ( 
.A(n_3207),
.Y(n_3783)
);

NOR2xp67_ASAP7_75t_L g3784 ( 
.A(n_3244),
.B(n_2849),
.Y(n_3784)
);

AO32x2_ASAP7_75t_L g3785 ( 
.A1(n_3341),
.A2(n_3069),
.A3(n_3076),
.B1(n_3064),
.B2(n_3063),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3443),
.B(n_511),
.Y(n_3786)
);

AND2x4_ASAP7_75t_L g3787 ( 
.A(n_3252),
.B(n_2775),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_L g3788 ( 
.A1(n_3721),
.A2(n_3083),
.B(n_3079),
.Y(n_3788)
);

O2A1O1Ixp33_ASAP7_75t_SL g3789 ( 
.A1(n_3483),
.A2(n_3092),
.B(n_3094),
.C(n_3087),
.Y(n_3789)
);

AOI21xp5_ASAP7_75t_L g3790 ( 
.A1(n_3722),
.A2(n_3110),
.B(n_3108),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3667),
.A2(n_3464),
.B(n_3484),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3572),
.A2(n_2787),
.B(n_3113),
.Y(n_3792)
);

BUFx3_ASAP7_75t_L g3793 ( 
.A(n_3255),
.Y(n_3793)
);

NAND3xp33_ASAP7_75t_SL g3794 ( 
.A(n_3469),
.B(n_2786),
.C(n_2902),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_L g3795 ( 
.A1(n_3616),
.A2(n_3152),
.B(n_3147),
.Y(n_3795)
);

OR2x2_ASAP7_75t_L g3796 ( 
.A(n_3380),
.B(n_3117),
.Y(n_3796)
);

OAI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3601),
.A2(n_3175),
.B(n_3163),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3278),
.Y(n_3798)
);

OAI21x1_ASAP7_75t_L g3799 ( 
.A1(n_3601),
.A2(n_3179),
.B(n_3177),
.Y(n_3799)
);

OAI21x1_ASAP7_75t_L g3800 ( 
.A1(n_3649),
.A2(n_3189),
.B(n_3180),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3269),
.B(n_3124),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3515),
.B(n_2851),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_SL g3803 ( 
.A(n_3294),
.B(n_3371),
.Y(n_3803)
);

OAI21x1_ASAP7_75t_L g3804 ( 
.A1(n_3292),
.A2(n_3198),
.B(n_3130),
.Y(n_3804)
);

OAI21x1_ASAP7_75t_L g3805 ( 
.A1(n_3451),
.A2(n_3131),
.B(n_3126),
.Y(n_3805)
);

OR2x2_ASAP7_75t_L g3806 ( 
.A(n_3313),
.B(n_3135),
.Y(n_3806)
);

A2O1A1Ixp33_ASAP7_75t_L g3807 ( 
.A1(n_3683),
.A2(n_3141),
.B(n_3153),
.C(n_3137),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3736),
.A2(n_3193),
.B(n_3190),
.Y(n_3808)
);

AOI21xp5_ASAP7_75t_L g3809 ( 
.A1(n_3733),
.A2(n_2900),
.B(n_2876),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3282),
.Y(n_3810)
);

OAI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3455),
.A2(n_2850),
.B(n_2927),
.Y(n_3811)
);

O2A1O1Ixp33_ASAP7_75t_SL g3812 ( 
.A1(n_3544),
.A2(n_2818),
.B(n_2828),
.C(n_2817),
.Y(n_3812)
);

A2O1A1Ixp33_ASAP7_75t_L g3813 ( 
.A1(n_3732),
.A2(n_2930),
.B(n_2934),
.C(n_2929),
.Y(n_3813)
);

BUFx6f_ASAP7_75t_L g3814 ( 
.A(n_3272),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_3733),
.A2(n_2946),
.B(n_2944),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3673),
.A2(n_511),
.B(n_512),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3214),
.A2(n_512),
.B(n_513),
.Y(n_3817)
);

A2O1A1Ixp33_ASAP7_75t_L g3818 ( 
.A1(n_3701),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_3818)
);

NOR2xp33_ASAP7_75t_L g3819 ( 
.A(n_3684),
.B(n_513),
.Y(n_3819)
);

OAI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3374),
.A2(n_514),
.B(n_515),
.Y(n_3820)
);

OAI22x1_ASAP7_75t_L g3821 ( 
.A1(n_3361),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_3821)
);

AOI21xp33_ASAP7_75t_L g3822 ( 
.A1(n_3527),
.A2(n_516),
.B(n_517),
.Y(n_3822)
);

AO31x2_ASAP7_75t_L g3823 ( 
.A1(n_3569),
.A2(n_518),
.A3(n_516),
.B(n_517),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3285),
.B(n_518),
.Y(n_3824)
);

AO31x2_ASAP7_75t_L g3825 ( 
.A1(n_3351),
.A2(n_520),
.A3(n_518),
.B(n_519),
.Y(n_3825)
);

AOI21xp5_ASAP7_75t_L g3826 ( 
.A1(n_3694),
.A2(n_519),
.B(n_520),
.Y(n_3826)
);

OA21x2_ASAP7_75t_L g3827 ( 
.A1(n_3525),
.A2(n_520),
.B(n_521),
.Y(n_3827)
);

AO31x2_ASAP7_75t_L g3828 ( 
.A1(n_3663),
.A2(n_523),
.A3(n_521),
.B(n_522),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3702),
.A2(n_521),
.B(n_522),
.Y(n_3829)
);

NAND3x1_ASAP7_75t_L g3830 ( 
.A(n_3336),
.B(n_523),
.C(n_524),
.Y(n_3830)
);

A2O1A1Ixp33_ASAP7_75t_L g3831 ( 
.A1(n_3317),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3445),
.B(n_525),
.Y(n_3832)
);

OAI22xp5_ASAP7_75t_L g3833 ( 
.A1(n_3244),
.A2(n_3560),
.B1(n_3352),
.B2(n_3372),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3290),
.B(n_526),
.Y(n_3834)
);

BUFx3_ASAP7_75t_L g3835 ( 
.A(n_3299),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3231),
.Y(n_3836)
);

BUFx3_ASAP7_75t_L g3837 ( 
.A(n_3299),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3296),
.B(n_526),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3244),
.B(n_527),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3315),
.Y(n_3840)
);

AOI21x1_ASAP7_75t_L g3841 ( 
.A1(n_3348),
.A2(n_605),
.B(n_604),
.Y(n_3841)
);

O2A1O1Ixp33_ASAP7_75t_SL g3842 ( 
.A1(n_3565),
.A2(n_530),
.B(n_527),
.C(n_529),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3249),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3261),
.Y(n_3844)
);

AND2x4_ASAP7_75t_L g3845 ( 
.A(n_3224),
.B(n_527),
.Y(n_3845)
);

AOI21xp5_ASAP7_75t_L g3846 ( 
.A1(n_3710),
.A2(n_530),
.B(n_531),
.Y(n_3846)
);

OAI21x1_ASAP7_75t_L g3847 ( 
.A1(n_3734),
.A2(n_532),
.B(n_531),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3257),
.B(n_530),
.Y(n_3848)
);

OAI21x1_ASAP7_75t_L g3849 ( 
.A1(n_3717),
.A2(n_534),
.B(n_533),
.Y(n_3849)
);

AO31x2_ASAP7_75t_L g3850 ( 
.A1(n_3669),
.A2(n_534),
.A3(n_532),
.B(n_533),
.Y(n_3850)
);

OAI21x1_ASAP7_75t_L g3851 ( 
.A1(n_3717),
.A2(n_535),
.B(n_534),
.Y(n_3851)
);

OA21x2_ASAP7_75t_L g3852 ( 
.A1(n_3542),
.A2(n_533),
.B(n_535),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3441),
.B(n_3427),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3554),
.B(n_535),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3477),
.B(n_536),
.Y(n_3855)
);

NOR2xp67_ASAP7_75t_SL g3856 ( 
.A(n_3309),
.B(n_3365),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3716),
.A2(n_536),
.B(n_537),
.Y(n_3857)
);

INVxp67_ASAP7_75t_L g3858 ( 
.A(n_3378),
.Y(n_3858)
);

OAI22xp5_ASAP7_75t_L g3859 ( 
.A1(n_3391),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_3859)
);

OAI21x1_ASAP7_75t_L g3860 ( 
.A1(n_3251),
.A2(n_3418),
.B(n_3463),
.Y(n_3860)
);

CKINVDCx5p33_ASAP7_75t_R g3861 ( 
.A(n_3397),
.Y(n_3861)
);

OAI22xp5_ASAP7_75t_SL g3862 ( 
.A1(n_3399),
.A2(n_539),
.B1(n_537),
.B2(n_538),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3263),
.Y(n_3863)
);

OAI21x1_ASAP7_75t_L g3864 ( 
.A1(n_3655),
.A2(n_541),
.B(n_540),
.Y(n_3864)
);

AO31x2_ASAP7_75t_L g3865 ( 
.A1(n_3448),
.A2(n_541),
.A3(n_539),
.B(n_540),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3289),
.Y(n_3866)
);

AO31x2_ASAP7_75t_L g3867 ( 
.A1(n_3598),
.A2(n_543),
.A3(n_540),
.B(n_542),
.Y(n_3867)
);

A2O1A1Ixp33_ASAP7_75t_L g3868 ( 
.A1(n_3627),
.A2(n_3221),
.B(n_3238),
.C(n_3395),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3385),
.B(n_542),
.Y(n_3869)
);

OAI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3600),
.A2(n_542),
.B(n_543),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3603),
.A2(n_543),
.B(n_544),
.Y(n_3871)
);

OAI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3595),
.A2(n_3473),
.B(n_3506),
.Y(n_3872)
);

BUFx2_ASAP7_75t_L g3873 ( 
.A(n_3557),
.Y(n_3873)
);

AOI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3728),
.A2(n_544),
.B(n_545),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3350),
.A2(n_544),
.B(n_545),
.Y(n_3875)
);

AOI221x1_ASAP7_75t_L g3876 ( 
.A1(n_3403),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.C(n_549),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3368),
.A2(n_546),
.B(n_547),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_SL g3878 ( 
.A(n_3259),
.B(n_546),
.Y(n_3878)
);

AOI221x1_ASAP7_75t_L g3879 ( 
.A1(n_3715),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.C(n_550),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3520),
.B(n_548),
.Y(n_3880)
);

INVx2_ASAP7_75t_SL g3881 ( 
.A(n_3711),
.Y(n_3881)
);

AND2x4_ASAP7_75t_L g3882 ( 
.A(n_3382),
.B(n_549),
.Y(n_3882)
);

NAND3xp33_ASAP7_75t_SL g3883 ( 
.A(n_3209),
.B(n_550),
.C(n_551),
.Y(n_3883)
);

AOI221x1_ASAP7_75t_L g3884 ( 
.A1(n_3612),
.A2(n_552),
.B1(n_550),
.B2(n_551),
.C(n_553),
.Y(n_3884)
);

BUFx10_ASAP7_75t_L g3885 ( 
.A(n_3265),
.Y(n_3885)
);

NOR2xp67_ASAP7_75t_L g3886 ( 
.A(n_3404),
.B(n_551),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_SL g3887 ( 
.A1(n_3430),
.A2(n_552),
.B(n_553),
.Y(n_3887)
);

NAND2x1p5_ASAP7_75t_L g3888 ( 
.A(n_3345),
.B(n_552),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3375),
.A2(n_554),
.B(n_555),
.Y(n_3889)
);

O2A1O1Ixp5_ASAP7_75t_SL g3890 ( 
.A1(n_3646),
.A2(n_608),
.B(n_609),
.C(n_607),
.Y(n_3890)
);

OAI21x1_ASAP7_75t_L g3891 ( 
.A1(n_3580),
.A2(n_554),
.B(n_555),
.Y(n_3891)
);

CKINVDCx5p33_ASAP7_75t_R g3892 ( 
.A(n_3401),
.Y(n_3892)
);

INVx5_ASAP7_75t_L g3893 ( 
.A(n_3406),
.Y(n_3893)
);

AND2x4_ASAP7_75t_L g3894 ( 
.A(n_3246),
.B(n_554),
.Y(n_3894)
);

OAI21x1_ASAP7_75t_SL g3895 ( 
.A1(n_3562),
.A2(n_3651),
.B(n_3431),
.Y(n_3895)
);

OAI21x1_ASAP7_75t_L g3896 ( 
.A1(n_3580),
.A2(n_555),
.B(n_556),
.Y(n_3896)
);

AO32x2_ASAP7_75t_L g3897 ( 
.A1(n_3384),
.A2(n_558),
.A3(n_556),
.B1(n_557),
.B2(n_559),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3488),
.B(n_3497),
.Y(n_3898)
);

AOI22xp33_ASAP7_75t_SL g3899 ( 
.A1(n_3570),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_L g3900 ( 
.A(n_3571),
.B(n_557),
.Y(n_3900)
);

O2A1O1Ixp5_ASAP7_75t_L g3901 ( 
.A1(n_3533),
.A2(n_560),
.B(n_558),
.C(n_559),
.Y(n_3901)
);

INVxp67_ASAP7_75t_L g3902 ( 
.A(n_3503),
.Y(n_3902)
);

OAI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_3573),
.A2(n_560),
.B(n_561),
.Y(n_3903)
);

OAI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3349),
.A2(n_560),
.B(n_561),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3305),
.B(n_562),
.Y(n_3905)
);

NOR4xp25_ASAP7_75t_L g3906 ( 
.A(n_3369),
.B(n_564),
.C(n_562),
.D(n_563),
.Y(n_3906)
);

AO31x2_ASAP7_75t_L g3907 ( 
.A1(n_3712),
.A2(n_564),
.A3(n_562),
.B(n_563),
.Y(n_3907)
);

BUFx3_ASAP7_75t_L g3908 ( 
.A(n_3482),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3320),
.B(n_564),
.Y(n_3909)
);

A2O1A1Ixp33_ASAP7_75t_L g3910 ( 
.A1(n_3513),
.A2(n_568),
.B(n_566),
.C(n_567),
.Y(n_3910)
);

AOI21xp5_ASAP7_75t_L g3911 ( 
.A1(n_3405),
.A2(n_566),
.B(n_567),
.Y(n_3911)
);

AO21x2_ASAP7_75t_L g3912 ( 
.A1(n_3383),
.A2(n_566),
.B(n_567),
.Y(n_3912)
);

HB1xp67_ASAP7_75t_L g3913 ( 
.A(n_3658),
.Y(n_3913)
);

A2O1A1Ixp33_ASAP7_75t_L g3914 ( 
.A1(n_3564),
.A2(n_570),
.B(n_568),
.C(n_569),
.Y(n_3914)
);

AOI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_3691),
.A2(n_568),
.B(n_569),
.Y(n_3915)
);

AOI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_3697),
.A2(n_569),
.B(n_570),
.Y(n_3916)
);

AND2x6_ASAP7_75t_L g3917 ( 
.A(n_3494),
.B(n_571),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3454),
.B(n_571),
.Y(n_3918)
);

OAI21x1_ASAP7_75t_L g3919 ( 
.A1(n_3591),
.A2(n_571),
.B(n_573),
.Y(n_3919)
);

OAI21xp5_ASAP7_75t_SL g3920 ( 
.A1(n_3310),
.A2(n_573),
.B(n_574),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3335),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3729),
.A2(n_573),
.B(n_574),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3433),
.Y(n_3923)
);

OAI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3591),
.A2(n_574),
.B(n_575),
.Y(n_3924)
);

AOI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3311),
.A2(n_575),
.B(n_576),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3419),
.A2(n_576),
.B(n_577),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3462),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3536),
.B(n_576),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_3449),
.A2(n_577),
.B(n_607),
.Y(n_3929)
);

NOR2xp33_ASAP7_75t_L g3930 ( 
.A(n_3597),
.B(n_577),
.Y(n_3930)
);

NOR2xp67_ASAP7_75t_L g3931 ( 
.A(n_3362),
.B(n_610),
.Y(n_3931)
);

INVx3_ASAP7_75t_L g3932 ( 
.A(n_3548),
.Y(n_3932)
);

OAI21x1_ASAP7_75t_L g3933 ( 
.A1(n_3293),
.A2(n_610),
.B(n_611),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3321),
.Y(n_3934)
);

AND2x4_ASAP7_75t_L g3935 ( 
.A(n_3283),
.B(n_3501),
.Y(n_3935)
);

OAI21x1_ASAP7_75t_L g3936 ( 
.A1(n_3354),
.A2(n_611),
.B(n_613),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3467),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_SL g3938 ( 
.A1(n_3494),
.A2(n_613),
.B(n_614),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3453),
.A2(n_614),
.B(n_615),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3552),
.B(n_615),
.Y(n_3940)
);

BUFx3_ASAP7_75t_L g3941 ( 
.A(n_3387),
.Y(n_3941)
);

NAND3xp33_ASAP7_75t_L g3942 ( 
.A(n_3585),
.B(n_617),
.C(n_618),
.Y(n_3942)
);

CKINVDCx12_ASAP7_75t_R g3943 ( 
.A(n_3240),
.Y(n_3943)
);

OAI22xp33_ASAP7_75t_L g3944 ( 
.A1(n_3226),
.A2(n_3236),
.B1(n_3233),
.B2(n_3444),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3458),
.A2(n_617),
.B(n_619),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_SL g3946 ( 
.A(n_3432),
.B(n_619),
.Y(n_3946)
);

INVx3_ASAP7_75t_L g3947 ( 
.A(n_3664),
.Y(n_3947)
);

A2O1A1Ixp33_ASAP7_75t_L g3948 ( 
.A1(n_3639),
.A2(n_622),
.B(n_620),
.C(n_621),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3566),
.B(n_621),
.Y(n_3949)
);

NAND2x1p5_ASAP7_75t_L g3950 ( 
.A(n_3406),
.B(n_959),
.Y(n_3950)
);

AO31x2_ASAP7_75t_L g3951 ( 
.A1(n_3326),
.A2(n_625),
.A3(n_623),
.B(n_624),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3589),
.B(n_623),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3295),
.B(n_959),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3333),
.Y(n_3954)
);

AO31x2_ASAP7_75t_L g3955 ( 
.A1(n_3212),
.A2(n_627),
.A3(n_625),
.B(n_626),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_L g3956 ( 
.A(n_3537),
.B(n_626),
.Y(n_3956)
);

A2O1A1Ixp33_ASAP7_75t_L g3957 ( 
.A1(n_3507),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_3957)
);

A2O1A1Ixp33_ASAP7_75t_L g3958 ( 
.A1(n_3521),
.A2(n_632),
.B(n_630),
.C(n_631),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3466),
.A2(n_631),
.B(n_633),
.Y(n_3959)
);

A2O1A1Ixp33_ASAP7_75t_L g3960 ( 
.A1(n_3618),
.A2(n_636),
.B(n_634),
.C(n_635),
.Y(n_3960)
);

AO31x2_ASAP7_75t_L g3961 ( 
.A1(n_3504),
.A2(n_637),
.A3(n_634),
.B(n_635),
.Y(n_3961)
);

NOR2xp33_ASAP7_75t_L g3962 ( 
.A(n_3402),
.B(n_3615),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3478),
.A2(n_637),
.B(n_638),
.Y(n_3963)
);

AO31x2_ASAP7_75t_L g3964 ( 
.A1(n_3366),
.A2(n_642),
.A3(n_639),
.B(n_640),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3247),
.Y(n_3965)
);

OR2x6_ASAP7_75t_L g3966 ( 
.A(n_3635),
.B(n_639),
.Y(n_3966)
);

INVx3_ASAP7_75t_L g3967 ( 
.A(n_3555),
.Y(n_3967)
);

AOI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3459),
.A2(n_642),
.B(n_643),
.Y(n_3968)
);

OAI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3626),
.A2(n_644),
.B(n_646),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3514),
.B(n_644),
.Y(n_3970)
);

AO31x2_ASAP7_75t_L g3971 ( 
.A1(n_3379),
.A2(n_649),
.A3(n_647),
.B(n_648),
.Y(n_3971)
);

AOI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3550),
.A2(n_648),
.B(n_649),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3502),
.A2(n_650),
.B(n_651),
.Y(n_3973)
);

OAI21xp5_ASAP7_75t_SL g3974 ( 
.A1(n_3582),
.A2(n_650),
.B(n_651),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3270),
.Y(n_3975)
);

CKINVDCx9p33_ASAP7_75t_R g3976 ( 
.A(n_3508),
.Y(n_3976)
);

BUFx2_ASAP7_75t_L g3977 ( 
.A(n_3685),
.Y(n_3977)
);

OAI21x1_ASAP7_75t_L g3978 ( 
.A1(n_3706),
.A2(n_653),
.B(n_655),
.Y(n_3978)
);

OAI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_3358),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.Y(n_3979)
);

O2A1O1Ixp33_ASAP7_75t_L g3980 ( 
.A1(n_3398),
.A2(n_659),
.B(n_656),
.C(n_658),
.Y(n_3980)
);

BUFx2_ASAP7_75t_SL g3981 ( 
.A(n_3437),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3376),
.Y(n_3982)
);

AO21x2_ASAP7_75t_L g3983 ( 
.A1(n_3641),
.A2(n_3643),
.B(n_3524),
.Y(n_3983)
);

OAI21xp5_ASAP7_75t_L g3984 ( 
.A1(n_3628),
.A2(n_659),
.B(n_660),
.Y(n_3984)
);

OAI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3654),
.A2(n_660),
.B(n_661),
.Y(n_3985)
);

BUFx6f_ASAP7_75t_L g3986 ( 
.A(n_3579),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3377),
.Y(n_3987)
);

AND2x4_ASAP7_75t_L g3988 ( 
.A(n_3437),
.B(n_958),
.Y(n_3988)
);

OAI21x1_ASAP7_75t_L g3989 ( 
.A1(n_3706),
.A2(n_662),
.B(n_663),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_3632),
.B(n_662),
.Y(n_3990)
);

OAI21x1_ASAP7_75t_L g3991 ( 
.A1(n_3660),
.A2(n_663),
.B(n_664),
.Y(n_3991)
);

INVx1_ASAP7_75t_SL g3992 ( 
.A(n_3480),
.Y(n_3992)
);

AO31x2_ASAP7_75t_L g3993 ( 
.A1(n_3528),
.A2(n_666),
.A3(n_664),
.B(n_665),
.Y(n_3993)
);

INVx1_ASAP7_75t_SL g3994 ( 
.A(n_3587),
.Y(n_3994)
);

O2A1O1Ixp33_ASAP7_75t_SL g3995 ( 
.A1(n_3234),
.A2(n_667),
.B(n_665),
.C(n_666),
.Y(n_3995)
);

AOI21xp33_ASAP7_75t_L g3996 ( 
.A1(n_3461),
.A2(n_667),
.B(n_668),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3340),
.B(n_668),
.Y(n_3997)
);

INVx4_ASAP7_75t_L g3998 ( 
.A(n_3407),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_SL g3999 ( 
.A(n_3432),
.B(n_670),
.Y(n_3999)
);

NOR4xp25_ASAP7_75t_L g4000 ( 
.A(n_3396),
.B(n_673),
.C(n_671),
.D(n_672),
.Y(n_4000)
);

OR2x2_ASAP7_75t_L g4001 ( 
.A(n_3661),
.B(n_671),
.Y(n_4001)
);

BUFx2_ASAP7_75t_L g4002 ( 
.A(n_3498),
.Y(n_4002)
);

AOI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3492),
.A2(n_673),
.B(n_674),
.Y(n_4003)
);

BUFx3_ASAP7_75t_L g4004 ( 
.A(n_3424),
.Y(n_4004)
);

AOI22xp33_ASAP7_75t_L g4005 ( 
.A1(n_3416),
.A2(n_676),
.B1(n_674),
.B2(n_675),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3393),
.Y(n_4006)
);

AO31x2_ASAP7_75t_L g4007 ( 
.A1(n_3447),
.A2(n_677),
.A3(n_675),
.B(n_676),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3273),
.Y(n_4008)
);

OAI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3672),
.A2(n_677),
.B(n_678),
.Y(n_4009)
);

BUFx6f_ASAP7_75t_L g4010 ( 
.A(n_3579),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3298),
.B(n_678),
.Y(n_4011)
);

BUFx4f_ASAP7_75t_L g4012 ( 
.A(n_3442),
.Y(n_4012)
);

A2O1A1Ixp33_ASAP7_75t_L g4013 ( 
.A1(n_3535),
.A2(n_681),
.B(n_679),
.C(n_680),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3411),
.B(n_679),
.Y(n_4014)
);

BUFx6f_ASAP7_75t_L g4015 ( 
.A(n_3579),
.Y(n_4015)
);

NOR2xp33_ASAP7_75t_L g4016 ( 
.A(n_3529),
.B(n_682),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3432),
.B(n_3577),
.Y(n_4017)
);

AND2x4_ASAP7_75t_L g4018 ( 
.A(n_3442),
.B(n_683),
.Y(n_4018)
);

CKINVDCx8_ASAP7_75t_R g4019 ( 
.A(n_3534),
.Y(n_4019)
);

OAI21x1_ASAP7_75t_SL g4020 ( 
.A1(n_3486),
.A2(n_683),
.B(n_685),
.Y(n_4020)
);

INVxp67_ASAP7_75t_L g4021 ( 
.A(n_3360),
.Y(n_4021)
);

BUFx12f_ASAP7_75t_L g4022 ( 
.A(n_3510),
.Y(n_4022)
);

OAI21xp33_ASAP7_75t_L g4023 ( 
.A1(n_3530),
.A2(n_686),
.B(n_687),
.Y(n_4023)
);

BUFx6f_ASAP7_75t_L g4024 ( 
.A(n_3581),
.Y(n_4024)
);

A2O1A1Ixp33_ASAP7_75t_L g4025 ( 
.A1(n_3593),
.A2(n_688),
.B(n_686),
.C(n_687),
.Y(n_4025)
);

AND2x4_ASAP7_75t_L g4026 ( 
.A(n_3561),
.B(n_3563),
.Y(n_4026)
);

A2O1A1Ixp33_ASAP7_75t_L g4027 ( 
.A1(n_3630),
.A2(n_691),
.B(n_689),
.C(n_690),
.Y(n_4027)
);

NAND3xp33_ASAP7_75t_L g4028 ( 
.A(n_3465),
.B(n_690),
.C(n_691),
.Y(n_4028)
);

BUFx6f_ASAP7_75t_L g4029 ( 
.A(n_3581),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3665),
.Y(n_4030)
);

O2A1O1Ixp33_ASAP7_75t_SL g4031 ( 
.A1(n_3288),
.A2(n_694),
.B(n_692),
.C(n_693),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3496),
.B(n_957),
.Y(n_4032)
);

O2A1O1Ixp33_ASAP7_75t_SL g4033 ( 
.A1(n_3220),
.A2(n_696),
.B(n_692),
.C(n_694),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3410),
.B(n_697),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3415),
.Y(n_4035)
);

INVx1_ASAP7_75t_SL g4036 ( 
.A(n_3534),
.Y(n_4036)
);

AOI21xp33_ASAP7_75t_L g4037 ( 
.A1(n_3493),
.A2(n_697),
.B(n_698),
.Y(n_4037)
);

O2A1O1Ixp33_ASAP7_75t_L g4038 ( 
.A1(n_3264),
.A2(n_701),
.B(n_699),
.C(n_700),
.Y(n_4038)
);

A2O1A1Ixp33_ASAP7_75t_L g4039 ( 
.A1(n_3682),
.A2(n_702),
.B(n_699),
.C(n_700),
.Y(n_4039)
);

OAI21x1_ASAP7_75t_L g4040 ( 
.A1(n_3723),
.A2(n_702),
.B(n_703),
.Y(n_4040)
);

AO31x2_ASAP7_75t_L g4041 ( 
.A1(n_3489),
.A2(n_705),
.A3(n_703),
.B(n_704),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3567),
.B(n_704),
.Y(n_4042)
);

AO31x2_ASAP7_75t_L g4043 ( 
.A1(n_3617),
.A2(n_708),
.A3(n_706),
.B(n_707),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3590),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3208),
.B(n_706),
.Y(n_4045)
);

BUFx2_ASAP7_75t_L g4046 ( 
.A(n_3498),
.Y(n_4046)
);

NAND3xp33_ASAP7_75t_L g4047 ( 
.A(n_3549),
.B(n_708),
.C(n_709),
.Y(n_4047)
);

A2O1A1Ixp33_ASAP7_75t_L g4048 ( 
.A1(n_3322),
.A2(n_712),
.B(n_709),
.C(n_710),
.Y(n_4048)
);

O2A1O1Ixp5_ASAP7_75t_L g4049 ( 
.A1(n_3568),
.A2(n_713),
.B(n_710),
.C(n_712),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3422),
.Y(n_4050)
);

INVx3_ASAP7_75t_L g4051 ( 
.A(n_3531),
.Y(n_4051)
);

INVx3_ASAP7_75t_L g4052 ( 
.A(n_3531),
.Y(n_4052)
);

AO31x2_ASAP7_75t_L g4053 ( 
.A1(n_3617),
.A2(n_716),
.A3(n_714),
.B(n_715),
.Y(n_4053)
);

OAI21x1_ASAP7_75t_L g4054 ( 
.A1(n_3217),
.A2(n_714),
.B(n_715),
.Y(n_4054)
);

BUFx12f_ASAP7_75t_L g4055 ( 
.A(n_3538),
.Y(n_4055)
);

AOI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_3735),
.A2(n_3206),
.B(n_3205),
.Y(n_4056)
);

INVx1_ASAP7_75t_SL g4057 ( 
.A(n_3976),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3761),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3764),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3776),
.Y(n_4060)
);

BUFx2_ASAP7_75t_L g4061 ( 
.A(n_3873),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3777),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3781),
.Y(n_4063)
);

CKINVDCx11_ASAP7_75t_R g4064 ( 
.A(n_3775),
.Y(n_4064)
);

OAI21xp5_ASAP7_75t_SL g4065 ( 
.A1(n_3920),
.A2(n_3613),
.B(n_3390),
.Y(n_4065)
);

BUFx8_ASAP7_75t_L g4066 ( 
.A(n_4055),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3745),
.A2(n_3412),
.B1(n_3389),
.B2(n_3679),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3745),
.A2(n_3883),
.B1(n_3944),
.B2(n_3917),
.Y(n_4068)
);

BUFx2_ASAP7_75t_L g4069 ( 
.A(n_4002),
.Y(n_4069)
);

BUFx6f_ASAP7_75t_L g4070 ( 
.A(n_3783),
.Y(n_4070)
);

INVx2_ASAP7_75t_SL g4071 ( 
.A(n_3835),
.Y(n_4071)
);

BUFx6f_ASAP7_75t_L g4072 ( 
.A(n_3768),
.Y(n_4072)
);

CKINVDCx11_ASAP7_75t_R g4073 ( 
.A(n_3885),
.Y(n_4073)
);

CKINVDCx11_ASAP7_75t_R g4074 ( 
.A(n_3758),
.Y(n_4074)
);

AOI22xp33_ASAP7_75t_L g4075 ( 
.A1(n_3745),
.A2(n_3337),
.B1(n_3719),
.B2(n_3635),
.Y(n_4075)
);

AOI22xp33_ASAP7_75t_SL g4076 ( 
.A1(n_3981),
.A2(n_3432),
.B1(n_3576),
.B2(n_3703),
.Y(n_4076)
);

CKINVDCx20_ASAP7_75t_R g4077 ( 
.A(n_3748),
.Y(n_4077)
);

AOI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3917),
.A2(n_3604),
.B1(n_3731),
.B2(n_3267),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3934),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_4019),
.A2(n_3638),
.B1(n_3621),
.B2(n_3327),
.Y(n_4080)
);

BUFx2_ASAP7_75t_L g4081 ( 
.A(n_4046),
.Y(n_4081)
);

CKINVDCx5p33_ASAP7_75t_R g4082 ( 
.A(n_3837),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3954),
.Y(n_4083)
);

BUFx3_ASAP7_75t_L g4084 ( 
.A(n_3793),
.Y(n_4084)
);

BUFx2_ASAP7_75t_SL g4085 ( 
.A(n_3908),
.Y(n_4085)
);

BUFx2_ASAP7_75t_L g4086 ( 
.A(n_4012),
.Y(n_4086)
);

AOI22xp33_ASAP7_75t_L g4087 ( 
.A1(n_3917),
.A2(n_3731),
.B1(n_3268),
.B2(n_3302),
.Y(n_4087)
);

BUFx8_ASAP7_75t_L g4088 ( 
.A(n_3814),
.Y(n_4088)
);

OAI21xp5_ASAP7_75t_SL g4089 ( 
.A1(n_3974),
.A2(n_3291),
.B(n_3370),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3862),
.A2(n_3318),
.B1(n_3306),
.B2(n_3657),
.Y(n_4090)
);

BUFx2_ASAP7_75t_L g4091 ( 
.A(n_3768),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3798),
.Y(n_4092)
);

OAI22xp33_ASAP7_75t_L g4093 ( 
.A1(n_3966),
.A2(n_3280),
.B1(n_3574),
.B2(n_3620),
.Y(n_4093)
);

CKINVDCx20_ASAP7_75t_R g4094 ( 
.A(n_3861),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3810),
.Y(n_4095)
);

BUFx6f_ASAP7_75t_L g4096 ( 
.A(n_3814),
.Y(n_4096)
);

INVx4_ASAP7_75t_L g4097 ( 
.A(n_3893),
.Y(n_4097)
);

AOI22xp33_ASAP7_75t_SL g4098 ( 
.A1(n_3966),
.A2(n_3432),
.B1(n_3636),
.B2(n_3611),
.Y(n_4098)
);

INVx2_ASAP7_75t_SL g4099 ( 
.A(n_3893),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_3853),
.B(n_3648),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3840),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3923),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3786),
.B(n_3648),
.Y(n_4103)
);

INVx6_ASAP7_75t_L g4104 ( 
.A(n_3998),
.Y(n_4104)
);

BUFx6f_ASAP7_75t_L g4105 ( 
.A(n_3986),
.Y(n_4105)
);

INVx6_ASAP7_75t_L g4106 ( 
.A(n_3780),
.Y(n_4106)
);

BUFx4f_ASAP7_75t_SL g4107 ( 
.A(n_4022),
.Y(n_4107)
);

BUFx8_ASAP7_75t_L g4108 ( 
.A(n_3740),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_3982),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_3744),
.B(n_3332),
.Y(n_4110)
);

OAI22xp5_ASAP7_75t_L g4111 ( 
.A1(n_3755),
.A2(n_3631),
.B1(n_3594),
.B2(n_3556),
.Y(n_4111)
);

INVx6_ASAP7_75t_SL g4112 ( 
.A(n_3935),
.Y(n_4112)
);

AOI22xp33_ASAP7_75t_L g4113 ( 
.A1(n_3760),
.A2(n_3359),
.B1(n_3386),
.B2(n_3677),
.Y(n_4113)
);

INVx3_ASAP7_75t_L g4114 ( 
.A(n_3739),
.Y(n_4114)
);

INVx6_ASAP7_75t_L g4115 ( 
.A(n_4026),
.Y(n_4115)
);

AOI22xp33_ASAP7_75t_L g4116 ( 
.A1(n_3773),
.A2(n_3394),
.B1(n_3413),
.B2(n_3400),
.Y(n_4116)
);

CKINVDCx11_ASAP7_75t_R g4117 ( 
.A(n_3941),
.Y(n_4117)
);

OAI22xp5_ASAP7_75t_L g4118 ( 
.A1(n_4036),
.A2(n_3556),
.B1(n_3316),
.B2(n_3676),
.Y(n_4118)
);

HB1xp67_ASAP7_75t_L g4119 ( 
.A(n_3913),
.Y(n_4119)
);

BUFx12f_ASAP7_75t_L g4120 ( 
.A(n_3892),
.Y(n_4120)
);

INVx1_ASAP7_75t_SL g4121 ( 
.A(n_4004),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3927),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3937),
.Y(n_4123)
);

BUFx3_ASAP7_75t_L g4124 ( 
.A(n_3977),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3965),
.B(n_3656),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_SL g4126 ( 
.A1(n_3742),
.A2(n_3611),
.B1(n_3636),
.B2(n_3676),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3771),
.B(n_3637),
.Y(n_4127)
);

BUFx3_ASAP7_75t_L g4128 ( 
.A(n_3932),
.Y(n_4128)
);

AOI22xp33_ASAP7_75t_L g4129 ( 
.A1(n_3822),
.A2(n_3438),
.B1(n_3450),
.B2(n_3434),
.Y(n_4129)
);

INVx1_ASAP7_75t_SL g4130 ( 
.A(n_3803),
.Y(n_4130)
);

OAI22xp33_ASAP7_75t_L g4131 ( 
.A1(n_3878),
.A2(n_3476),
.B1(n_3688),
.B2(n_3670),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3855),
.B(n_3652),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3921),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_3987),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_4006),
.Y(n_4135)
);

OAI22xp5_ASAP7_75t_L g4136 ( 
.A1(n_3988),
.A2(n_3446),
.B1(n_3546),
.B2(n_3707),
.Y(n_4136)
);

INVxp67_ASAP7_75t_L g4137 ( 
.A(n_3962),
.Y(n_4137)
);

BUFx2_ASAP7_75t_L g4138 ( 
.A(n_3986),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3843),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3975),
.B(n_3730),
.Y(n_4140)
);

CKINVDCx11_ASAP7_75t_R g4141 ( 
.A(n_3898),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_4010),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3863),
.Y(n_4143)
);

INVx2_ASAP7_75t_SL g4144 ( 
.A(n_3881),
.Y(n_4144)
);

AOI22xp33_ASAP7_75t_L g4145 ( 
.A1(n_3895),
.A2(n_3408),
.B1(n_3429),
.B2(n_3426),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3866),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4044),
.Y(n_4147)
);

AOI22xp33_ASAP7_75t_L g4148 ( 
.A1(n_3820),
.A2(n_3452),
.B1(n_3686),
.B2(n_3718),
.Y(n_4148)
);

AOI21xp5_ASAP7_75t_L g4149 ( 
.A1(n_3772),
.A2(n_3578),
.B(n_3539),
.Y(n_4149)
);

CKINVDCx5p33_ASAP7_75t_R g4150 ( 
.A(n_3943),
.Y(n_4150)
);

BUFx8_ASAP7_75t_SL g4151 ( 
.A(n_3845),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_3832),
.B(n_3693),
.Y(n_4152)
);

CKINVDCx20_ASAP7_75t_R g4153 ( 
.A(n_3743),
.Y(n_4153)
);

AOI22xp33_ASAP7_75t_SL g4154 ( 
.A1(n_4018),
.A2(n_3689),
.B1(n_3538),
.B2(n_3541),
.Y(n_4154)
);

INVx8_ASAP7_75t_L g4155 ( 
.A(n_3882),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3754),
.Y(n_4156)
);

AOI22xp5_ASAP7_75t_L g4157 ( 
.A1(n_3819),
.A2(n_3308),
.B1(n_3258),
.B2(n_3650),
.Y(n_4157)
);

AOI22xp33_ASAP7_75t_L g4158 ( 
.A1(n_3903),
.A2(n_3592),
.B1(n_3640),
.B2(n_3727),
.Y(n_4158)
);

CKINVDCx20_ASAP7_75t_R g4159 ( 
.A(n_3759),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4008),
.B(n_3614),
.Y(n_4160)
);

BUFx3_ASAP7_75t_L g4161 ( 
.A(n_3947),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4030),
.B(n_3622),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3836),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3844),
.Y(n_4164)
);

CKINVDCx20_ASAP7_75t_R g4165 ( 
.A(n_3756),
.Y(n_4165)
);

INVx6_ASAP7_75t_L g4166 ( 
.A(n_4010),
.Y(n_4166)
);

CKINVDCx6p67_ASAP7_75t_R g4167 ( 
.A(n_3821),
.Y(n_4167)
);

BUFx6f_ASAP7_75t_L g4168 ( 
.A(n_4015),
.Y(n_4168)
);

AOI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3769),
.A2(n_3490),
.B1(n_3519),
.B2(n_3634),
.Y(n_4169)
);

INVx5_ASAP7_75t_L g4170 ( 
.A(n_4015),
.Y(n_4170)
);

CKINVDCx11_ASAP7_75t_R g4171 ( 
.A(n_3992),
.Y(n_4171)
);

AOI22xp33_ASAP7_75t_SL g4172 ( 
.A1(n_3833),
.A2(n_3695),
.B1(n_3690),
.B2(n_3671),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_4035),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_L g4174 ( 
.A1(n_3872),
.A2(n_3559),
.B1(n_3248),
.B2(n_3254),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4050),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_3849),
.Y(n_4176)
);

OAI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_3942),
.A2(n_3642),
.B1(n_3645),
.B2(n_3436),
.Y(n_4177)
);

OAI22xp5_ASAP7_75t_L g4178 ( 
.A1(n_3868),
.A2(n_3356),
.B1(n_3357),
.B2(n_3342),
.Y(n_4178)
);

HB1xp67_ASAP7_75t_L g4179 ( 
.A(n_3858),
.Y(n_4179)
);

OAI22xp33_ASAP7_75t_L g4180 ( 
.A1(n_3888),
.A2(n_4028),
.B1(n_3886),
.B2(n_3979),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4001),
.Y(n_4181)
);

OAI22xp5_ASAP7_75t_L g4182 ( 
.A1(n_4005),
.A2(n_3479),
.B1(n_3421),
.B2(n_3704),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_SL g4183 ( 
.A1(n_4020),
.A2(n_3695),
.B1(n_3629),
.B2(n_3705),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_3828),
.Y(n_4184)
);

AOI22xp33_ASAP7_75t_L g4185 ( 
.A1(n_4021),
.A2(n_3262),
.B1(n_3266),
.B2(n_3237),
.Y(n_4185)
);

OAI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_3950),
.A2(n_3428),
.B1(n_3219),
.B2(n_3241),
.Y(n_4186)
);

INVx4_ASAP7_75t_L g4187 ( 
.A(n_4024),
.Y(n_4187)
);

AOI22xp33_ASAP7_75t_L g4188 ( 
.A1(n_4023),
.A2(n_3277),
.B1(n_3281),
.B2(n_3271),
.Y(n_4188)
);

INVx4_ASAP7_75t_L g4189 ( 
.A(n_4024),
.Y(n_4189)
);

OAI22xp5_ASAP7_75t_L g4190 ( 
.A1(n_4025),
.A2(n_3239),
.B1(n_3256),
.B2(n_3243),
.Y(n_4190)
);

BUFx4f_ASAP7_75t_SL g4191 ( 
.A(n_3994),
.Y(n_4191)
);

AOI22xp33_ASAP7_75t_L g4192 ( 
.A1(n_3870),
.A2(n_3287),
.B1(n_3297),
.B2(n_3284),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3828),
.Y(n_4193)
);

AOI21xp33_ASAP7_75t_L g4194 ( 
.A1(n_3782),
.A2(n_3276),
.B(n_3509),
.Y(n_4194)
);

BUFx2_ASAP7_75t_L g4195 ( 
.A(n_4029),
.Y(n_4195)
);

BUFx3_ASAP7_75t_L g4196 ( 
.A(n_4029),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_3850),
.Y(n_4197)
);

CKINVDCx5p33_ASAP7_75t_R g4198 ( 
.A(n_3990),
.Y(n_4198)
);

CKINVDCx11_ASAP7_75t_R g4199 ( 
.A(n_3894),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3850),
.Y(n_4200)
);

NAND2x1p5_ASAP7_75t_L g4201 ( 
.A(n_3856),
.B(n_3581),
.Y(n_4201)
);

CKINVDCx20_ASAP7_75t_R g4202 ( 
.A(n_3900),
.Y(n_4202)
);

AOI22xp33_ASAP7_75t_L g4203 ( 
.A1(n_3802),
.A2(n_3303),
.B1(n_3319),
.B2(n_3301),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3824),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3834),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3838),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3869),
.B(n_3460),
.Y(n_4207)
);

INVx1_ASAP7_75t_SL g4208 ( 
.A(n_3967),
.Y(n_4208)
);

INVx3_ASAP7_75t_L g4209 ( 
.A(n_4051),
.Y(n_4209)
);

INVx1_ASAP7_75t_SL g4210 ( 
.A(n_4052),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_4000),
.B(n_3329),
.Y(n_4211)
);

CKINVDCx20_ASAP7_75t_R g4212 ( 
.A(n_3902),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_3796),
.B(n_3330),
.Y(n_4213)
);

BUFx2_ASAP7_75t_L g4214 ( 
.A(n_4011),
.Y(n_4214)
);

HB1xp67_ASAP7_75t_L g4215 ( 
.A(n_3801),
.Y(n_4215)
);

CKINVDCx11_ASAP7_75t_R g4216 ( 
.A(n_3757),
.Y(n_4216)
);

BUFx12f_ASAP7_75t_L g4217 ( 
.A(n_3787),
.Y(n_4217)
);

AOI22xp33_ASAP7_75t_SL g4218 ( 
.A1(n_3912),
.A2(n_3705),
.B1(n_3692),
.B2(n_3596),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_4042),
.B(n_3511),
.Y(n_4219)
);

OAI22xp5_ASAP7_75t_L g4220 ( 
.A1(n_3931),
.A2(n_3899),
.B1(n_3938),
.B2(n_3887),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3905),
.Y(n_4221)
);

OAI21xp33_ASAP7_75t_L g4222 ( 
.A1(n_3906),
.A2(n_3485),
.B(n_3275),
.Y(n_4222)
);

AOI22xp33_ASAP7_75t_L g4223 ( 
.A1(n_4047),
.A2(n_3325),
.B1(n_3328),
.B2(n_3323),
.Y(n_4223)
);

BUFx12f_ASAP7_75t_L g4224 ( 
.A(n_3806),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3909),
.Y(n_4225)
);

AOI22xp33_ASAP7_75t_L g4226 ( 
.A1(n_3930),
.A2(n_3344),
.B1(n_3346),
.B2(n_3338),
.Y(n_4226)
);

INVx6_ASAP7_75t_L g4227 ( 
.A(n_3970),
.Y(n_4227)
);

AOI22xp33_ASAP7_75t_SL g4228 ( 
.A1(n_3791),
.A2(n_3692),
.B1(n_3602),
.B2(n_3279),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3851),
.Y(n_4229)
);

INVx3_ASAP7_75t_L g4230 ( 
.A(n_3830),
.Y(n_4230)
);

AOI22xp33_ASAP7_75t_L g4231 ( 
.A1(n_3996),
.A2(n_3355),
.B1(n_3364),
.B2(n_3353),
.Y(n_4231)
);

AOI22xp33_ASAP7_75t_SL g4232 ( 
.A1(n_3956),
.A2(n_3692),
.B1(n_3602),
.B2(n_3286),
.Y(n_4232)
);

AOI22xp33_ASAP7_75t_L g4233 ( 
.A1(n_3918),
.A2(n_3409),
.B1(n_3414),
.B2(n_3392),
.Y(n_4233)
);

INVx6_ASAP7_75t_L g4234 ( 
.A(n_3839),
.Y(n_4234)
);

AOI22xp33_ASAP7_75t_SL g4235 ( 
.A1(n_3827),
.A2(n_3324),
.B1(n_3260),
.B2(n_3681),
.Y(n_4235)
);

BUFx2_ASAP7_75t_L g4236 ( 
.A(n_4040),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_3891),
.Y(n_4237)
);

INVx6_ASAP7_75t_L g4238 ( 
.A(n_3784),
.Y(n_4238)
);

BUFx4_ASAP7_75t_R g4239 ( 
.A(n_3897),
.Y(n_4239)
);

BUFx3_ASAP7_75t_L g4240 ( 
.A(n_3880),
.Y(n_4240)
);

BUFx12f_ASAP7_75t_L g4241 ( 
.A(n_3876),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4043),
.Y(n_4242)
);

BUFx8_ASAP7_75t_SL g4243 ( 
.A(n_3854),
.Y(n_4243)
);

BUFx2_ASAP7_75t_L g4244 ( 
.A(n_4043),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4053),
.Y(n_4245)
);

AOI22xp33_ASAP7_75t_SL g4246 ( 
.A1(n_3852),
.A2(n_3681),
.B1(n_3633),
.B2(n_3675),
.Y(n_4246)
);

BUFx4f_ASAP7_75t_SL g4247 ( 
.A(n_4017),
.Y(n_4247)
);

INVx6_ASAP7_75t_L g4248 ( 
.A(n_4016),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_4079),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4181),
.B(n_3928),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4184),
.Y(n_4251)
);

AO21x2_ASAP7_75t_L g4252 ( 
.A1(n_4242),
.A2(n_4245),
.B(n_4197),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_4083),
.Y(n_4253)
);

OAI21x1_ASAP7_75t_L g4254 ( 
.A1(n_4149),
.A2(n_3737),
.B(n_3751),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_4109),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_4134),
.Y(n_4256)
);

INVx2_ASAP7_75t_L g4257 ( 
.A(n_4135),
.Y(n_4257)
);

BUFx2_ASAP7_75t_L g4258 ( 
.A(n_4069),
.Y(n_4258)
);

BUFx2_ASAP7_75t_L g4259 ( 
.A(n_4081),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4058),
.Y(n_4260)
);

OR2x2_ASAP7_75t_L g4261 ( 
.A(n_4119),
.B(n_3865),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4100),
.B(n_3825),
.Y(n_4262)
);

AOI21x1_ASAP7_75t_L g4263 ( 
.A1(n_4244),
.A2(n_3841),
.B(n_4056),
.Y(n_4263)
);

OAI21x1_ASAP7_75t_L g4264 ( 
.A1(n_4237),
.A2(n_3741),
.B(n_3860),
.Y(n_4264)
);

BUFx3_ASAP7_75t_L g4265 ( 
.A(n_4070),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4059),
.Y(n_4266)
);

AO21x1_ASAP7_75t_L g4267 ( 
.A1(n_4093),
.A2(n_4180),
.B(n_4220),
.Y(n_4267)
);

INVx2_ASAP7_75t_SL g4268 ( 
.A(n_4104),
.Y(n_4268)
);

AND2x4_ASAP7_75t_L g4269 ( 
.A(n_4215),
.B(n_3825),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4173),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4060),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4062),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4063),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4156),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4092),
.Y(n_4275)
);

AO21x2_ASAP7_75t_L g4276 ( 
.A1(n_4193),
.A2(n_3972),
.B(n_3968),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4095),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4103),
.B(n_3865),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4163),
.Y(n_4279)
);

BUFx6f_ASAP7_75t_L g4280 ( 
.A(n_4072),
.Y(n_4280)
);

INVx3_ASAP7_75t_L g4281 ( 
.A(n_4097),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4207),
.B(n_4053),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4101),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_4164),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4175),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4214),
.B(n_4132),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4139),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4143),
.Y(n_4288)
);

BUFx2_ASAP7_75t_L g4289 ( 
.A(n_4112),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4102),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4122),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4123),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4133),
.Y(n_4293)
);

CKINVDCx14_ASAP7_75t_R g4294 ( 
.A(n_4070),
.Y(n_4294)
);

BUFx6f_ASAP7_75t_L g4295 ( 
.A(n_4072),
.Y(n_4295)
);

INVx3_ASAP7_75t_L g4296 ( 
.A(n_4217),
.Y(n_4296)
);

INVxp67_ASAP7_75t_L g4297 ( 
.A(n_4061),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_4152),
.B(n_4007),
.Y(n_4298)
);

INVx3_ASAP7_75t_L g4299 ( 
.A(n_4238),
.Y(n_4299)
);

AOI22xp33_ASAP7_75t_L g4300 ( 
.A1(n_4068),
.A2(n_3794),
.B1(n_3766),
.B2(n_3859),
.Y(n_4300)
);

INVxp67_ASAP7_75t_SL g4301 ( 
.A(n_4224),
.Y(n_4301)
);

AND2x2_ASAP7_75t_L g4302 ( 
.A(n_4127),
.B(n_4007),
.Y(n_4302)
);

HB1xp67_ASAP7_75t_L g4303 ( 
.A(n_4179),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4147),
.Y(n_4304)
);

OAI21x1_ASAP7_75t_L g4305 ( 
.A1(n_4176),
.A2(n_3809),
.B(n_3770),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4146),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4160),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4162),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4140),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4200),
.Y(n_4310)
);

OAI21x1_ASAP7_75t_L g4311 ( 
.A1(n_4229),
.A2(n_3805),
.B(n_3804),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4236),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4219),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4221),
.Y(n_4314)
);

NOR2xp33_ASAP7_75t_L g4315 ( 
.A(n_4243),
.B(n_4045),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4238),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4213),
.Y(n_4317)
);

AOI22xp33_ASAP7_75t_L g4318 ( 
.A1(n_4167),
.A2(n_3767),
.B1(n_3984),
.B2(n_3969),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4239),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4225),
.Y(n_4320)
);

AOI21x1_ASAP7_75t_L g4321 ( 
.A1(n_4211),
.A2(n_3999),
.B(n_3946),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4204),
.Y(n_4322)
);

BUFx2_ASAP7_75t_L g4323 ( 
.A(n_4112),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4205),
.Y(n_4324)
);

AOI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_4065),
.A2(n_3699),
.B1(n_4032),
.B2(n_3848),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4206),
.Y(n_4326)
);

AOI222xp33_ASAP7_75t_L g4327 ( 
.A1(n_4089),
.A2(n_4014),
.B1(n_3953),
.B2(n_3334),
.C1(n_3997),
.C2(n_4009),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4110),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_4125),
.B(n_3940),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4210),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4208),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4209),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4105),
.Y(n_4333)
);

AOI22xp5_ASAP7_75t_L g4334 ( 
.A1(n_4075),
.A2(n_3958),
.B1(n_4034),
.B2(n_3778),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4227),
.B(n_4041),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4227),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4114),
.Y(n_4337)
);

INVx3_ASAP7_75t_L g4338 ( 
.A(n_4201),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4099),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4091),
.Y(n_4340)
);

BUFx6f_ASAP7_75t_L g4341 ( 
.A(n_4105),
.Y(n_4341)
);

INVx2_ASAP7_75t_SL g4342 ( 
.A(n_4104),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4241),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4194),
.A2(n_3749),
.B(n_3747),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4138),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4142),
.Y(n_4346)
);

OA21x2_ASAP7_75t_L g4347 ( 
.A1(n_4169),
.A2(n_3847),
.B(n_3879),
.Y(n_4347)
);

BUFx3_ASAP7_75t_L g4348 ( 
.A(n_4088),
.Y(n_4348)
);

BUFx2_ASAP7_75t_L g4349 ( 
.A(n_4159),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4240),
.B(n_4041),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4168),
.Y(n_4351)
);

CKINVDCx20_ASAP7_75t_R g4352 ( 
.A(n_4066),
.Y(n_4352)
);

BUFx4f_ASAP7_75t_SL g4353 ( 
.A(n_4066),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4195),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4165),
.Y(n_4355)
);

OAI21x1_ASAP7_75t_L g4356 ( 
.A1(n_4145),
.A2(n_3815),
.B(n_3790),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_4137),
.B(n_3823),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4057),
.Y(n_4358)
);

NAND2xp33_ASAP7_75t_SL g4359 ( 
.A(n_4153),
.B(n_3983),
.Y(n_4359)
);

BUFx3_ASAP7_75t_L g4360 ( 
.A(n_4088),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4121),
.B(n_3823),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_4098),
.B(n_3949),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4168),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4130),
.Y(n_4364)
);

OAI21x1_ASAP7_75t_L g4365 ( 
.A1(n_4113),
.A2(n_3788),
.B(n_3800),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4161),
.Y(n_4366)
);

INVxp33_ASAP7_75t_L g4367 ( 
.A(n_4151),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4218),
.Y(n_4368)
);

BUFx8_ASAP7_75t_SL g4369 ( 
.A(n_4077),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4246),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4196),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4235),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4155),
.B(n_3952),
.Y(n_4373)
);

HB1xp67_ASAP7_75t_L g4374 ( 
.A(n_4170),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4166),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4247),
.Y(n_4376)
);

HB1xp67_ASAP7_75t_L g4377 ( 
.A(n_4170),
.Y(n_4377)
);

INVx2_ASAP7_75t_SL g4378 ( 
.A(n_4084),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4166),
.Y(n_4379)
);

AO32x2_ASAP7_75t_L g4380 ( 
.A1(n_4378),
.A2(n_4071),
.A3(n_4118),
.B1(n_4080),
.B2(n_4111),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4317),
.B(n_4222),
.Y(n_4381)
);

OR2x2_ASAP7_75t_L g4382 ( 
.A(n_4313),
.B(n_4317),
.Y(n_4382)
);

AND2x2_ASAP7_75t_L g4383 ( 
.A(n_4286),
.B(n_4096),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4357),
.B(n_4067),
.Y(n_4384)
);

A2O1A1Ixp33_ASAP7_75t_L g4385 ( 
.A1(n_4338),
.A2(n_4230),
.B(n_4155),
.C(n_4086),
.Y(n_4385)
);

OR2x6_ASAP7_75t_L g4386 ( 
.A(n_4348),
.B(n_4085),
.Y(n_4386)
);

OAI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_4344),
.A2(n_4154),
.B(n_4131),
.Y(n_4387)
);

AOI221xp5_ASAP7_75t_L g4388 ( 
.A1(n_4267),
.A2(n_4177),
.B1(n_4325),
.B2(n_4303),
.C(n_4372),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4258),
.B(n_4096),
.Y(n_4389)
);

O2A1O1Ixp33_ASAP7_75t_L g4390 ( 
.A1(n_4327),
.A2(n_4186),
.B(n_4190),
.C(n_4136),
.Y(n_4390)
);

OA21x2_ASAP7_75t_L g4391 ( 
.A1(n_4343),
.A2(n_3884),
.B(n_3978),
.Y(n_4391)
);

A2O1A1Ixp33_ASAP7_75t_L g4392 ( 
.A1(n_4338),
.A2(n_4124),
.B(n_4087),
.C(n_4126),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4298),
.B(n_4157),
.Y(n_4393)
);

AOI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4334),
.A2(n_4078),
.B1(n_4234),
.B2(n_4248),
.Y(n_4394)
);

AOI221xp5_ASAP7_75t_L g4395 ( 
.A1(n_4372),
.A2(n_4178),
.B1(n_4037),
.B2(n_4174),
.C(n_4226),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_4302),
.B(n_4076),
.Y(n_4396)
);

AND2x4_ASAP7_75t_L g4397 ( 
.A(n_4259),
.B(n_4187),
.Y(n_4397)
);

AND2x2_ASAP7_75t_L g4398 ( 
.A(n_4319),
.B(n_4115),
.Y(n_4398)
);

AO32x1_ASAP7_75t_L g4399 ( 
.A1(n_4343),
.A2(n_4189),
.A3(n_4144),
.B1(n_4182),
.B2(n_3532),
.Y(n_4399)
);

BUFx2_ASAP7_75t_L g4400 ( 
.A(n_4281),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4319),
.B(n_4331),
.Y(n_4401)
);

AOI221xp5_ASAP7_75t_L g4402 ( 
.A1(n_4328),
.A2(n_4185),
.B1(n_3926),
.B2(n_4090),
.C(n_3871),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4364),
.B(n_4115),
.Y(n_4403)
);

NAND2x1p5_ASAP7_75t_L g4404 ( 
.A(n_4360),
.B(n_4170),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4330),
.B(n_4216),
.Y(n_4405)
);

OR2x2_ASAP7_75t_L g4406 ( 
.A(n_4324),
.B(n_4128),
.Y(n_4406)
);

OAI21xp5_ASAP7_75t_L g4407 ( 
.A1(n_4318),
.A2(n_3991),
.B(n_3875),
.Y(n_4407)
);

CKINVDCx5p33_ASAP7_75t_R g4408 ( 
.A(n_4353),
.Y(n_4408)
);

BUFx2_ASAP7_75t_L g4409 ( 
.A(n_4281),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_4249),
.Y(n_4410)
);

A2O1A1Ixp33_ASAP7_75t_L g4411 ( 
.A1(n_4268),
.A2(n_4232),
.B(n_4150),
.C(n_4172),
.Y(n_4411)
);

OR2x2_ASAP7_75t_L g4412 ( 
.A(n_4324),
.B(n_3993),
.Y(n_4412)
);

AOI22xp5_ASAP7_75t_L g4413 ( 
.A1(n_4362),
.A2(n_4234),
.B1(n_4248),
.B2(n_4202),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4340),
.B(n_4171),
.Y(n_4414)
);

CKINVDCx10_ASAP7_75t_R g4415 ( 
.A(n_4352),
.Y(n_4415)
);

AND2x6_ASAP7_75t_L g4416 ( 
.A(n_4368),
.B(n_3681),
.Y(n_4416)
);

O2A1O1Ixp33_ASAP7_75t_L g4417 ( 
.A1(n_4329),
.A2(n_3910),
.B(n_3914),
.C(n_3818),
.Y(n_4417)
);

AO21x2_ASAP7_75t_L g4418 ( 
.A1(n_4263),
.A2(n_3904),
.B(n_3925),
.Y(n_4418)
);

AND2x6_ASAP7_75t_L g4419 ( 
.A(n_4368),
.B(n_4199),
.Y(n_4419)
);

OA21x2_ASAP7_75t_L g4420 ( 
.A1(n_4370),
.A2(n_3989),
.B(n_3919),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4309),
.B(n_4307),
.Y(n_4421)
);

AND2x2_ASAP7_75t_L g4422 ( 
.A(n_4345),
.B(n_4106),
.Y(n_4422)
);

OAI21x1_ASAP7_75t_L g4423 ( 
.A1(n_4365),
.A2(n_3924),
.B(n_3896),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4260),
.Y(n_4424)
);

BUFx2_ASAP7_75t_L g4425 ( 
.A(n_4374),
.Y(n_4425)
);

OR2x2_ASAP7_75t_L g4426 ( 
.A(n_4287),
.B(n_3993),
.Y(n_4426)
);

NOR2xp33_ASAP7_75t_SL g4427 ( 
.A(n_4265),
.B(n_4107),
.Y(n_4427)
);

OR2x2_ASAP7_75t_L g4428 ( 
.A(n_4288),
.B(n_3955),
.Y(n_4428)
);

HB1xp67_ASAP7_75t_L g4429 ( 
.A(n_4297),
.Y(n_4429)
);

NOR2xp33_ASAP7_75t_L g4430 ( 
.A(n_4342),
.B(n_4367),
.Y(n_4430)
);

AOI211xp5_ASAP7_75t_L g4431 ( 
.A1(n_4370),
.A2(n_4359),
.B(n_4278),
.C(n_4262),
.Y(n_4431)
);

OAI22xp5_ASAP7_75t_L g4432 ( 
.A1(n_4349),
.A2(n_4116),
.B1(n_4212),
.B2(n_4191),
.Y(n_4432)
);

AND2x2_ASAP7_75t_L g4433 ( 
.A(n_4346),
.B(n_4106),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4266),
.Y(n_4434)
);

INVx5_ASAP7_75t_L g4435 ( 
.A(n_4296),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4354),
.B(n_4228),
.Y(n_4436)
);

AND4x1_ASAP7_75t_L g4437 ( 
.A(n_4315),
.B(n_4064),
.C(n_4074),
.D(n_4073),
.Y(n_4437)
);

AND2x4_ASAP7_75t_L g4438 ( 
.A(n_4358),
.B(n_4082),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4308),
.B(n_3867),
.Y(n_4439)
);

INVx3_ASAP7_75t_L g4440 ( 
.A(n_4296),
.Y(n_4440)
);

AOI211xp5_ASAP7_75t_L g4441 ( 
.A1(n_4350),
.A2(n_3842),
.B(n_3985),
.C(n_3980),
.Y(n_4441)
);

AO32x2_ASAP7_75t_L g4442 ( 
.A1(n_4261),
.A2(n_4269),
.A3(n_4361),
.B1(n_4271),
.B2(n_4273),
.Y(n_4442)
);

OR2x6_ASAP7_75t_L g4443 ( 
.A(n_4289),
.B(n_4120),
.Y(n_4443)
);

AND2x4_ASAP7_75t_L g4444 ( 
.A(n_4336),
.B(n_3668),
.Y(n_4444)
);

INVx3_ASAP7_75t_L g4445 ( 
.A(n_4280),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4282),
.B(n_4183),
.Y(n_4446)
);

OAI21x1_ASAP7_75t_L g4447 ( 
.A1(n_4356),
.A2(n_3936),
.B(n_3933),
.Y(n_4447)
);

INVx4_ASAP7_75t_L g4448 ( 
.A(n_4323),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4314),
.B(n_4117),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4320),
.B(n_3867),
.Y(n_4450)
);

NOR2x1_ASAP7_75t_SL g4451 ( 
.A(n_4376),
.B(n_3229),
.Y(n_4451)
);

AO21x1_ASAP7_75t_SL g4452 ( 
.A1(n_4377),
.A2(n_4188),
.B(n_4192),
.Y(n_4452)
);

A2O1A1Ixp33_ASAP7_75t_L g4453 ( 
.A1(n_4301),
.A2(n_3889),
.B(n_3911),
.C(n_3877),
.Y(n_4453)
);

AOI22xp33_ASAP7_75t_L g4454 ( 
.A1(n_4300),
.A2(n_4223),
.B1(n_4203),
.B2(n_4231),
.Y(n_4454)
);

NOR2x1_ASAP7_75t_SL g4455 ( 
.A(n_4376),
.B(n_4280),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4335),
.B(n_4198),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4322),
.B(n_3897),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4253),
.Y(n_4458)
);

AOI22xp33_ASAP7_75t_L g4459 ( 
.A1(n_4388),
.A2(n_4355),
.B1(n_4269),
.B2(n_4347),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4424),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4456),
.B(n_4316),
.Y(n_4461)
);

NOR2x1p5_ASAP7_75t_L g4462 ( 
.A(n_4448),
.B(n_4299),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_SL g4463 ( 
.A(n_4400),
.B(n_4299),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_4401),
.B(n_4316),
.Y(n_4464)
);

INVx3_ASAP7_75t_L g4465 ( 
.A(n_4386),
.Y(n_4465)
);

AND2x2_ASAP7_75t_L g4466 ( 
.A(n_4383),
.B(n_4339),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4434),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4389),
.B(n_4366),
.Y(n_4468)
);

HB1xp67_ASAP7_75t_L g4469 ( 
.A(n_4425),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4403),
.B(n_4272),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4429),
.B(n_4275),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4398),
.B(n_4277),
.Y(n_4472)
);

HB1xp67_ASAP7_75t_L g4473 ( 
.A(n_4409),
.Y(n_4473)
);

INVx4_ASAP7_75t_L g4474 ( 
.A(n_4386),
.Y(n_4474)
);

AND2x2_ASAP7_75t_L g4475 ( 
.A(n_4422),
.B(n_4283),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4457),
.B(n_4306),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4433),
.B(n_4290),
.Y(n_4477)
);

NOR2x1_ASAP7_75t_L g4478 ( 
.A(n_4440),
.B(n_4371),
.Y(n_4478)
);

AND2x4_ASAP7_75t_L g4479 ( 
.A(n_4446),
.B(n_4312),
.Y(n_4479)
);

NOR2xp33_ASAP7_75t_L g4480 ( 
.A(n_4435),
.B(n_4294),
.Y(n_4480)
);

HB1xp67_ASAP7_75t_L g4481 ( 
.A(n_4406),
.Y(n_4481)
);

OR2x6_ASAP7_75t_L g4482 ( 
.A(n_4387),
.B(n_4312),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4382),
.Y(n_4483)
);

AND2x2_ASAP7_75t_L g4484 ( 
.A(n_4449),
.B(n_4291),
.Y(n_4484)
);

INVx1_ASAP7_75t_SL g4485 ( 
.A(n_4397),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4421),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4414),
.B(n_4292),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4436),
.B(n_4293),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4410),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4381),
.B(n_4304),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4458),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4393),
.B(n_4326),
.Y(n_4492)
);

OR2x2_ASAP7_75t_L g4493 ( 
.A(n_4384),
.B(n_4274),
.Y(n_4493)
);

OR2x2_ASAP7_75t_L g4494 ( 
.A(n_4396),
.B(n_4279),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4412),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4442),
.Y(n_4496)
);

BUFx2_ASAP7_75t_L g4497 ( 
.A(n_4435),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_4405),
.B(n_4332),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4442),
.B(n_4337),
.Y(n_4499)
);

OR2x2_ASAP7_75t_L g4500 ( 
.A(n_4426),
.B(n_4284),
.Y(n_4500)
);

INVx2_ASAP7_75t_L g4501 ( 
.A(n_4428),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4450),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4439),
.Y(n_4503)
);

BUFx2_ASAP7_75t_L g4504 ( 
.A(n_4404),
.Y(n_4504)
);

AND2x4_ASAP7_75t_L g4505 ( 
.A(n_4455),
.B(n_4252),
.Y(n_4505)
);

HB1xp67_ASAP7_75t_L g4506 ( 
.A(n_4445),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4438),
.B(n_4285),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4413),
.B(n_4255),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4431),
.B(n_4251),
.Y(n_4509)
);

NOR2xp33_ASAP7_75t_L g4510 ( 
.A(n_4427),
.B(n_4108),
.Y(n_4510)
);

NOR2xp67_ASAP7_75t_L g4511 ( 
.A(n_4394),
.B(n_4333),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4395),
.B(n_4251),
.Y(n_4512)
);

INVx3_ASAP7_75t_L g4513 ( 
.A(n_4416),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4420),
.Y(n_4514)
);

HB1xp67_ASAP7_75t_L g4515 ( 
.A(n_4447),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4430),
.B(n_4256),
.Y(n_4516)
);

HB1xp67_ASAP7_75t_L g4517 ( 
.A(n_4391),
.Y(n_4517)
);

AOI22xp33_ASAP7_75t_SL g4518 ( 
.A1(n_4419),
.A2(n_4108),
.B1(n_4341),
.B2(n_4295),
.Y(n_4518)
);

AOI22xp33_ASAP7_75t_L g4519 ( 
.A1(n_4419),
.A2(n_4347),
.B1(n_4233),
.B2(n_4373),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4454),
.B(n_4257),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_4423),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4390),
.B(n_4270),
.Y(n_4522)
);

AND2x4_ASAP7_75t_L g4523 ( 
.A(n_4416),
.B(n_4310),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4419),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4416),
.B(n_4250),
.Y(n_4525)
);

OR2x6_ASAP7_75t_L g4526 ( 
.A(n_4474),
.B(n_4443),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_4482),
.A2(n_4411),
.B(n_4399),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4520),
.B(n_4441),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4495),
.Y(n_4529)
);

AOI22xp33_ASAP7_75t_SL g4530 ( 
.A1(n_4474),
.A2(n_4432),
.B1(n_4451),
.B2(n_4380),
.Y(n_4530)
);

AOI33xp33_ASAP7_75t_L g4531 ( 
.A1(n_4459),
.A2(n_4402),
.A3(n_4417),
.B1(n_4129),
.B2(n_4148),
.B3(n_4158),
.Y(n_4531)
);

OR2x2_ASAP7_75t_L g4532 ( 
.A(n_4493),
.B(n_4305),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_4460),
.Y(n_4533)
);

AND2x2_ASAP7_75t_L g4534 ( 
.A(n_4479),
.B(n_4452),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4479),
.B(n_4443),
.Y(n_4535)
);

INVx3_ASAP7_75t_L g4536 ( 
.A(n_4505),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4467),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_4520),
.B(n_4407),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4481),
.B(n_4380),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4512),
.B(n_4392),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4471),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4512),
.B(n_4418),
.Y(n_4542)
);

NAND4xp25_ASAP7_75t_L g4543 ( 
.A(n_4519),
.B(n_4385),
.C(n_4453),
.D(n_3929),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_4473),
.Y(n_4544)
);

BUFx2_ASAP7_75t_L g4545 ( 
.A(n_4497),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4485),
.B(n_4351),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4485),
.B(n_4363),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4503),
.B(n_4502),
.Y(n_4548)
);

AND2x4_ASAP7_75t_L g4549 ( 
.A(n_4462),
.B(n_4375),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4461),
.B(n_4379),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_4469),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4486),
.Y(n_4552)
);

INVx2_ASAP7_75t_L g4553 ( 
.A(n_4501),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4500),
.Y(n_4554)
);

INVx3_ASAP7_75t_L g4555 ( 
.A(n_4505),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4517),
.Y(n_4556)
);

AOI33xp33_ASAP7_75t_L g4557 ( 
.A1(n_4518),
.A2(n_4524),
.A3(n_4492),
.B1(n_4496),
.B2(n_4488),
.B3(n_4484),
.Y(n_4557)
);

AND2x4_ASAP7_75t_SL g4558 ( 
.A(n_4480),
.B(n_4280),
.Y(n_4558)
);

INVx2_ASAP7_75t_SL g4559 ( 
.A(n_4465),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4476),
.Y(n_4560)
);

AOI22xp33_ASAP7_75t_SL g4561 ( 
.A1(n_4465),
.A2(n_4444),
.B1(n_4408),
.B2(n_4295),
.Y(n_4561)
);

AO21x2_ASAP7_75t_L g4562 ( 
.A1(n_4514),
.A2(n_4264),
.B(n_4311),
.Y(n_4562)
);

AND2x4_ASAP7_75t_SL g4563 ( 
.A(n_4510),
.B(n_4295),
.Y(n_4563)
);

AO21x2_ASAP7_75t_L g4564 ( 
.A1(n_4515),
.A2(n_4321),
.B(n_4254),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_4464),
.B(n_4341),
.Y(n_4565)
);

AND2x2_ASAP7_75t_L g4566 ( 
.A(n_4468),
.B(n_4341),
.Y(n_4566)
);

INVxp67_ASAP7_75t_L g4567 ( 
.A(n_4478),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4489),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4470),
.B(n_4472),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4491),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_4509),
.B(n_3738),
.Y(n_4571)
);

AND2x2_ASAP7_75t_L g4572 ( 
.A(n_4475),
.B(n_4437),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4477),
.B(n_4276),
.Y(n_4573)
);

AOI22xp33_ASAP7_75t_L g4574 ( 
.A1(n_4482),
.A2(n_3922),
.B1(n_3826),
.B2(n_3874),
.Y(n_4574)
);

AOI221xp5_ASAP7_75t_L g4575 ( 
.A1(n_4522),
.A2(n_3216),
.B1(n_4033),
.B2(n_4031),
.C(n_3995),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4483),
.Y(n_4576)
);

AOI22xp33_ASAP7_75t_L g4577 ( 
.A1(n_4482),
.A2(n_3816),
.B1(n_3765),
.B2(n_3307),
.Y(n_4577)
);

AOI221x1_ASAP7_75t_L g4578 ( 
.A1(n_4522),
.A2(n_3753),
.B1(n_3808),
.B2(n_3779),
.C(n_4399),
.Y(n_4578)
);

INVx4_ASAP7_75t_L g4579 ( 
.A(n_4504),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4476),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4490),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4506),
.Y(n_4582)
);

OR2x2_ASAP7_75t_L g4583 ( 
.A(n_4494),
.B(n_3738),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4534),
.B(n_4499),
.Y(n_4584)
);

OR2x2_ASAP7_75t_L g4585 ( 
.A(n_4580),
.B(n_4490),
.Y(n_4585)
);

AND2x4_ASAP7_75t_SL g4586 ( 
.A(n_4526),
.B(n_4507),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4545),
.B(n_4516),
.Y(n_4587)
);

AND2x2_ASAP7_75t_L g4588 ( 
.A(n_4559),
.B(n_4466),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4581),
.B(n_4542),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_4579),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4538),
.B(n_4509),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4548),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4568),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4579),
.B(n_4487),
.Y(n_4594)
);

NOR2x1_ASAP7_75t_R g4595 ( 
.A(n_4572),
.B(n_4141),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_4580),
.B(n_4511),
.Y(n_4596)
);

OR2x2_ASAP7_75t_L g4597 ( 
.A(n_4560),
.B(n_4554),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4573),
.B(n_4498),
.Y(n_4598)
);

OR2x2_ASAP7_75t_L g4599 ( 
.A(n_4583),
.B(n_4529),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4529),
.B(n_4511),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4546),
.B(n_4508),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4568),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_4582),
.Y(n_4603)
);

INVx1_ASAP7_75t_SL g4604 ( 
.A(n_4547),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4566),
.B(n_4463),
.Y(n_4605)
);

HB1xp67_ASAP7_75t_L g4606 ( 
.A(n_4556),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4535),
.B(n_4565),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4571),
.B(n_4521),
.Y(n_4608)
);

INVx2_ASAP7_75t_L g4609 ( 
.A(n_4570),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4549),
.B(n_4513),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4570),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4552),
.Y(n_4612)
);

NOR2xp67_ASAP7_75t_L g4613 ( 
.A(n_4536),
.B(n_4513),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4533),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4528),
.B(n_4537),
.Y(n_4615)
);

NOR2x1_ASAP7_75t_L g4616 ( 
.A(n_4526),
.B(n_4523),
.Y(n_4616)
);

INVx1_ASAP7_75t_SL g4617 ( 
.A(n_4590),
.Y(n_4617)
);

AOI32xp33_ASAP7_75t_SL g4618 ( 
.A1(n_4615),
.A2(n_4540),
.A3(n_4556),
.B1(n_4541),
.B2(n_4557),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4585),
.Y(n_4619)
);

OR2x2_ASAP7_75t_L g4620 ( 
.A(n_4615),
.B(n_4532),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4612),
.Y(n_4621)
);

INVx2_ASAP7_75t_L g4622 ( 
.A(n_4603),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4616),
.B(n_4539),
.Y(n_4623)
);

AND2x2_ASAP7_75t_L g4624 ( 
.A(n_4610),
.B(n_4536),
.Y(n_4624)
);

HB1xp67_ASAP7_75t_L g4625 ( 
.A(n_4606),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4586),
.B(n_4555),
.Y(n_4626)
);

OR2x2_ASAP7_75t_L g4627 ( 
.A(n_4589),
.B(n_4551),
.Y(n_4627)
);

OR2x6_ASAP7_75t_L g4628 ( 
.A(n_4613),
.B(n_4527),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4614),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4604),
.B(n_4555),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4591),
.B(n_4592),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4591),
.B(n_4530),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4604),
.B(n_4567),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4584),
.B(n_4549),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4597),
.Y(n_4635)
);

INVxp67_ASAP7_75t_L g4636 ( 
.A(n_4595),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4593),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4602),
.Y(n_4638)
);

AOI211xp5_ASAP7_75t_L g4639 ( 
.A1(n_4594),
.A2(n_4543),
.B(n_4575),
.C(n_4523),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4609),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4611),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4589),
.B(n_4531),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4599),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4608),
.B(n_4576),
.Y(n_4644)
);

OR2x2_ASAP7_75t_L g4645 ( 
.A(n_4608),
.B(n_4544),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4598),
.B(n_4569),
.Y(n_4646)
);

INVx2_ASAP7_75t_L g4647 ( 
.A(n_4587),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4600),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4605),
.Y(n_4649)
);

INVx1_ASAP7_75t_SL g4650 ( 
.A(n_4588),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4596),
.B(n_4553),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_SL g4652 ( 
.A(n_4600),
.B(n_4561),
.Y(n_4652)
);

OR2x2_ASAP7_75t_L g4653 ( 
.A(n_4596),
.B(n_4525),
.Y(n_4653)
);

INVxp67_ASAP7_75t_L g4654 ( 
.A(n_4607),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_4601),
.B(n_4550),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4585),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4585),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4590),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4591),
.B(n_4564),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_L g4660 ( 
.A(n_4642),
.B(n_4525),
.Y(n_4660)
);

OR2x2_ASAP7_75t_L g4661 ( 
.A(n_4631),
.B(n_4564),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4625),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4617),
.B(n_4578),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4617),
.B(n_4574),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4626),
.B(n_4563),
.Y(n_4665)
);

NAND2x1_ASAP7_75t_SL g4666 ( 
.A(n_4633),
.B(n_4415),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4634),
.B(n_4558),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4624),
.B(n_4562),
.Y(n_4668)
);

BUFx2_ASAP7_75t_L g4669 ( 
.A(n_4636),
.Y(n_4669)
);

INVx3_ASAP7_75t_SL g4670 ( 
.A(n_4628),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4630),
.B(n_4562),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4648),
.B(n_4577),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4619),
.B(n_4656),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4657),
.B(n_3955),
.Y(n_4674)
);

NOR2x1_ASAP7_75t_L g4675 ( 
.A(n_4628),
.B(n_4094),
.Y(n_4675)
);

NOR2x1_ASAP7_75t_L g4676 ( 
.A(n_4628),
.B(n_4652),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4639),
.B(n_3951),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4639),
.B(n_3951),
.Y(n_4678)
);

NAND3xp33_ASAP7_75t_L g4679 ( 
.A(n_4632),
.B(n_3957),
.C(n_4027),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_L g4680 ( 
.A(n_4650),
.B(n_3964),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4627),
.Y(n_4681)
);

INVx2_ASAP7_75t_L g4682 ( 
.A(n_4658),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4650),
.B(n_3964),
.Y(n_4683)
);

INVx2_ASAP7_75t_L g4684 ( 
.A(n_4647),
.Y(n_4684)
);

OR2x2_ASAP7_75t_L g4685 ( 
.A(n_4620),
.B(n_4622),
.Y(n_4685)
);

AND2x2_ASAP7_75t_L g4686 ( 
.A(n_4623),
.B(n_3961),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4635),
.B(n_3971),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4643),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4654),
.B(n_3971),
.Y(n_4689)
);

INVxp67_ASAP7_75t_SL g4690 ( 
.A(n_4659),
.Y(n_4690)
);

OR2x2_ASAP7_75t_L g4691 ( 
.A(n_4645),
.B(n_3961),
.Y(n_4691)
);

INVx1_ASAP7_75t_SL g4692 ( 
.A(n_4653),
.Y(n_4692)
);

AND2x2_ASAP7_75t_L g4693 ( 
.A(n_4649),
.B(n_4646),
.Y(n_4693)
);

OR2x2_ASAP7_75t_L g4694 ( 
.A(n_4644),
.B(n_3907),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4621),
.B(n_3907),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4629),
.Y(n_4696)
);

OR2x2_ASAP7_75t_L g4697 ( 
.A(n_4651),
.B(n_3750),
.Y(n_4697)
);

NAND4xp25_ASAP7_75t_L g4698 ( 
.A(n_4659),
.B(n_3945),
.C(n_3959),
.D(n_3939),
.Y(n_4698)
);

AND2x2_ASAP7_75t_SL g4699 ( 
.A(n_4618),
.B(n_4369),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4637),
.B(n_3807),
.Y(n_4700)
);

AO21x1_ASAP7_75t_L g4701 ( 
.A1(n_4690),
.A2(n_4641),
.B(n_4638),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4662),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4682),
.Y(n_4703)
);

HB1xp67_ASAP7_75t_L g4704 ( 
.A(n_4692),
.Y(n_4704)
);

O2A1O1Ixp33_ASAP7_75t_L g4705 ( 
.A1(n_4669),
.A2(n_4039),
.B(n_3831),
.C(n_4048),
.Y(n_4705)
);

NAND2xp33_ASAP7_75t_SL g4706 ( 
.A(n_4666),
.B(n_4640),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4665),
.B(n_4655),
.Y(n_4707)
);

NAND3xp33_ASAP7_75t_SL g4708 ( 
.A(n_4677),
.B(n_3505),
.C(n_4038),
.Y(n_4708)
);

INVx3_ASAP7_75t_L g4709 ( 
.A(n_4670),
.Y(n_4709)
);

INVx1_ASAP7_75t_SL g4710 ( 
.A(n_4664),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4681),
.B(n_3817),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4699),
.B(n_3785),
.Y(n_4712)
);

HB1xp67_ASAP7_75t_L g4713 ( 
.A(n_4688),
.Y(n_4713)
);

AOI21xp33_ASAP7_75t_L g4714 ( 
.A1(n_4676),
.A2(n_717),
.B(n_719),
.Y(n_4714)
);

INVx1_ASAP7_75t_SL g4715 ( 
.A(n_4675),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4685),
.Y(n_4716)
);

NOR2xp33_ASAP7_75t_L g4717 ( 
.A(n_4675),
.B(n_4660),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4673),
.B(n_717),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4693),
.B(n_3785),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4684),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4672),
.B(n_3963),
.Y(n_4721)
);

OR2x2_ASAP7_75t_L g4722 ( 
.A(n_4694),
.B(n_719),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4678),
.B(n_4003),
.Y(n_4723)
);

BUFx2_ASAP7_75t_L g4724 ( 
.A(n_4676),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4696),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4697),
.Y(n_4726)
);

NAND4xp25_ASAP7_75t_L g4727 ( 
.A(n_4679),
.B(n_3846),
.C(n_3857),
.D(n_3829),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4700),
.Y(n_4728)
);

OAI22xp5_ASAP7_75t_L g4729 ( 
.A1(n_4663),
.A2(n_4686),
.B1(n_4689),
.B2(n_4661),
.Y(n_4729)
);

OAI22xp33_ASAP7_75t_L g4730 ( 
.A1(n_4691),
.A2(n_3915),
.B1(n_3916),
.B2(n_3774),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4674),
.B(n_4687),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4695),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4680),
.B(n_3973),
.Y(n_4733)
);

OR2x2_ASAP7_75t_L g4734 ( 
.A(n_4683),
.B(n_720),
.Y(n_4734)
);

NAND3xp33_ASAP7_75t_L g4735 ( 
.A(n_4709),
.B(n_4679),
.C(n_4671),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4704),
.B(n_4668),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4716),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4720),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4713),
.Y(n_4739)
);

OAI211xp5_ASAP7_75t_L g4740 ( 
.A1(n_4709),
.A2(n_4698),
.B(n_4667),
.C(n_3960),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4703),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4702),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4711),
.Y(n_4743)
);

INVxp67_ASAP7_75t_L g4744 ( 
.A(n_4724),
.Y(n_4744)
);

AOI21xp5_ASAP7_75t_L g4745 ( 
.A1(n_4706),
.A2(n_3763),
.B(n_3339),
.Y(n_4745)
);

OR2x2_ASAP7_75t_L g4746 ( 
.A(n_4710),
.B(n_720),
.Y(n_4746)
);

AOI31xp33_ASAP7_75t_L g4747 ( 
.A1(n_4714),
.A2(n_3547),
.A3(n_3584),
.B(n_3540),
.Y(n_4747)
);

OAI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_4715),
.A2(n_4717),
.B(n_4723),
.Y(n_4748)
);

NAND3xp33_ASAP7_75t_L g4749 ( 
.A(n_4728),
.B(n_3948),
.C(n_3901),
.Y(n_4749)
);

OR2x2_ASAP7_75t_L g4750 ( 
.A(n_4721),
.B(n_4734),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4707),
.Y(n_4751)
);

NAND4xp25_ASAP7_75t_L g4752 ( 
.A(n_4705),
.B(n_3425),
.C(n_3435),
.D(n_3417),
.Y(n_4752)
);

OAI21xp5_ASAP7_75t_SL g4753 ( 
.A1(n_4712),
.A2(n_3471),
.B(n_3439),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4732),
.B(n_722),
.Y(n_4754)
);

AOI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_4701),
.A2(n_3367),
.B1(n_3373),
.B2(n_3300),
.Y(n_4755)
);

INVx2_ASAP7_75t_L g4756 ( 
.A(n_4718),
.Y(n_4756)
);

NOR2x1_ASAP7_75t_L g4757 ( 
.A(n_4725),
.B(n_4722),
.Y(n_4757)
);

AOI22xp5_ASAP7_75t_L g4758 ( 
.A1(n_4708),
.A2(n_3726),
.B1(n_3713),
.B2(n_3347),
.Y(n_4758)
);

AOI21xp33_ASAP7_75t_L g4759 ( 
.A1(n_4729),
.A2(n_723),
.B(n_724),
.Y(n_4759)
);

NOR2xp33_ASAP7_75t_L g4760 ( 
.A(n_4726),
.B(n_724),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4733),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4719),
.B(n_725),
.Y(n_4762)
);

OR2x2_ASAP7_75t_L g4763 ( 
.A(n_4731),
.B(n_725),
.Y(n_4763)
);

HB1xp67_ASAP7_75t_L g4764 ( 
.A(n_4730),
.Y(n_4764)
);

INVx2_ASAP7_75t_L g4765 ( 
.A(n_4737),
.Y(n_4765)
);

XOR2xp5_ASAP7_75t_L g4766 ( 
.A(n_4751),
.B(n_4727),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4738),
.Y(n_4767)
);

NOR2xp33_ASAP7_75t_L g4768 ( 
.A(n_4744),
.B(n_4759),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4741),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4764),
.B(n_4727),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4739),
.Y(n_4771)
);

NOR2xp33_ASAP7_75t_L g4772 ( 
.A(n_4736),
.B(n_726),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4746),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4750),
.Y(n_4774)
);

AOI21xp33_ASAP7_75t_L g4775 ( 
.A1(n_4760),
.A2(n_726),
.B(n_727),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_4762),
.B(n_727),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4743),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4763),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4754),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4756),
.Y(n_4780)
);

AOI22xp5_ASAP7_75t_L g4781 ( 
.A1(n_4740),
.A2(n_3599),
.B1(n_3666),
.B2(n_3331),
.Y(n_4781)
);

XOR2xp5_ASAP7_75t_L g4782 ( 
.A(n_4748),
.B(n_728),
.Y(n_4782)
);

NOR2xp67_ASAP7_75t_SL g4783 ( 
.A(n_4735),
.B(n_3575),
.Y(n_4783)
);

AOI221xp5_ASAP7_75t_L g4784 ( 
.A1(n_4761),
.A2(n_3472),
.B1(n_3512),
.B2(n_3516),
.C(n_3495),
.Y(n_4784)
);

INVx1_ASAP7_75t_SL g4785 ( 
.A(n_4742),
.Y(n_4785)
);

AOI21xp5_ASAP7_75t_L g4786 ( 
.A1(n_4757),
.A2(n_4747),
.B(n_4745),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4753),
.B(n_728),
.Y(n_4787)
);

OR2x2_ASAP7_75t_L g4788 ( 
.A(n_4749),
.B(n_729),
.Y(n_4788)
);

AOI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4755),
.A2(n_3687),
.B(n_3789),
.Y(n_4789)
);

INVx2_ASAP7_75t_SL g4790 ( 
.A(n_4758),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4758),
.B(n_730),
.Y(n_4791)
);

NOR2x1_ASAP7_75t_L g4792 ( 
.A(n_4752),
.B(n_3653),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4751),
.B(n_730),
.Y(n_4793)
);

INVxp67_ASAP7_75t_L g4794 ( 
.A(n_4760),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4738),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4738),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4751),
.B(n_731),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4738),
.Y(n_4798)
);

NAND3xp33_ASAP7_75t_L g4799 ( 
.A(n_4768),
.B(n_3674),
.C(n_4049),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4772),
.B(n_732),
.Y(n_4800)
);

NAND4xp25_ASAP7_75t_L g4801 ( 
.A(n_4786),
.B(n_4013),
.C(n_3586),
.D(n_3605),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_SL g4802 ( 
.A(n_4765),
.B(n_3583),
.Y(n_4802)
);

NOR3xp33_ASAP7_75t_L g4803 ( 
.A(n_4787),
.B(n_3680),
.C(n_3678),
.Y(n_4803)
);

NOR2xp33_ASAP7_75t_L g4804 ( 
.A(n_4782),
.B(n_732),
.Y(n_4804)
);

NAND3xp33_ASAP7_75t_L g4805 ( 
.A(n_4767),
.B(n_3518),
.C(n_3607),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_SL g4806 ( 
.A(n_4795),
.B(n_3608),
.Y(n_4806)
);

BUFx3_ASAP7_75t_L g4807 ( 
.A(n_4769),
.Y(n_4807)
);

NOR4xp25_ASAP7_75t_L g4808 ( 
.A(n_4785),
.B(n_3720),
.C(n_3606),
.D(n_3644),
.Y(n_4808)
);

AND2x2_ASAP7_75t_L g4809 ( 
.A(n_4774),
.B(n_733),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_SL g4810 ( 
.A(n_4796),
.B(n_3609),
.Y(n_4810)
);

NOR2xp33_ASAP7_75t_L g4811 ( 
.A(n_4798),
.B(n_734),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4793),
.Y(n_4812)
);

AOI22xp5_ASAP7_75t_L g4813 ( 
.A1(n_4766),
.A2(n_3619),
.B1(n_3811),
.B2(n_3623),
.Y(n_4813)
);

OAI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4770),
.A2(n_3813),
.B1(n_3724),
.B2(n_3696),
.Y(n_4814)
);

OAI22xp5_ASAP7_75t_SL g4815 ( 
.A1(n_4790),
.A2(n_3227),
.B1(n_3363),
.B2(n_3213),
.Y(n_4815)
);

AOI22xp5_ASAP7_75t_L g4816 ( 
.A1(n_4794),
.A2(n_3491),
.B1(n_4054),
.B2(n_3812),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_SL g4817 ( 
.A(n_4780),
.B(n_3668),
.Y(n_4817)
);

NOR2xp33_ASAP7_75t_L g4818 ( 
.A(n_4797),
.B(n_734),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4783),
.B(n_4776),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4788),
.Y(n_4820)
);

OR2x2_ASAP7_75t_L g4821 ( 
.A(n_4791),
.B(n_735),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4771),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4778),
.B(n_735),
.Y(n_4823)
);

NOR2xp33_ASAP7_75t_L g4824 ( 
.A(n_4773),
.B(n_736),
.Y(n_4824)
);

NAND4xp25_ASAP7_75t_SL g4825 ( 
.A(n_4779),
.B(n_3708),
.C(n_3225),
.D(n_3890),
.Y(n_4825)
);

INVxp33_ASAP7_75t_L g4826 ( 
.A(n_4792),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4777),
.B(n_736),
.Y(n_4827)
);

AOI222xp33_ASAP7_75t_L g4828 ( 
.A1(n_4784),
.A2(n_3864),
.B1(n_3625),
.B2(n_3647),
.C1(n_3543),
.C2(n_3795),
.Y(n_4828)
);

NOR2xp33_ASAP7_75t_L g4829 ( 
.A(n_4775),
.B(n_737),
.Y(n_4829)
);

OAI21xp5_ASAP7_75t_SL g4830 ( 
.A1(n_4826),
.A2(n_4781),
.B(n_4789),
.Y(n_4830)
);

OAI21xp5_ASAP7_75t_L g4831 ( 
.A1(n_4824),
.A2(n_4811),
.B(n_4819),
.Y(n_4831)
);

AOI211xp5_ASAP7_75t_L g4832 ( 
.A1(n_4820),
.A2(n_4781),
.B(n_3700),
.C(n_3523),
.Y(n_4832)
);

AOI21xp33_ASAP7_75t_L g4833 ( 
.A1(n_4822),
.A2(n_737),
.B(n_738),
.Y(n_4833)
);

AOI222xp33_ASAP7_75t_L g4834 ( 
.A1(n_4807),
.A2(n_3792),
.B1(n_3799),
.B2(n_3797),
.C1(n_741),
.C2(n_745),
.Y(n_4834)
);

AND2x2_ASAP7_75t_L g4835 ( 
.A(n_4809),
.B(n_739),
.Y(n_4835)
);

AOI222xp33_ASAP7_75t_L g4836 ( 
.A1(n_4812),
.A2(n_741),
.B1(n_746),
.B2(n_739),
.C1(n_740),
.C2(n_743),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_4821),
.Y(n_4837)
);

O2A1O1Ixp33_ASAP7_75t_L g4838 ( 
.A1(n_4827),
.A2(n_747),
.B(n_743),
.C(n_746),
.Y(n_4838)
);

OAI221xp5_ASAP7_75t_SL g4839 ( 
.A1(n_4823),
.A2(n_4808),
.B1(n_4801),
.B2(n_4799),
.C(n_4813),
.Y(n_4839)
);

AOI221xp5_ASAP7_75t_L g4840 ( 
.A1(n_4804),
.A2(n_751),
.B1(n_748),
.B2(n_749),
.C(n_752),
.Y(n_4840)
);

OAI211xp5_ASAP7_75t_SL g4841 ( 
.A1(n_4817),
.A2(n_751),
.B(n_748),
.C(n_749),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4800),
.Y(n_4842)
);

O2A1O1Ixp33_ASAP7_75t_L g4843 ( 
.A1(n_4829),
.A2(n_754),
.B(n_752),
.C(n_753),
.Y(n_4843)
);

O2A1O1Ixp33_ASAP7_75t_L g4844 ( 
.A1(n_4818),
.A2(n_755),
.B(n_753),
.C(n_754),
.Y(n_4844)
);

AOI221xp5_ASAP7_75t_L g4845 ( 
.A1(n_4815),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.C(n_759),
.Y(n_4845)
);

OAI221xp5_ASAP7_75t_L g4846 ( 
.A1(n_4806),
.A2(n_3746),
.B1(n_761),
.B2(n_757),
.C(n_760),
.Y(n_4846)
);

OAI321xp33_ASAP7_75t_L g4847 ( 
.A1(n_4802),
.A2(n_3474),
.A3(n_3227),
.B1(n_3499),
.B2(n_3363),
.C(n_3213),
.Y(n_4847)
);

OAI221xp5_ASAP7_75t_SL g4848 ( 
.A1(n_4828),
.A2(n_763),
.B1(n_761),
.B2(n_762),
.C(n_765),
.Y(n_4848)
);

BUFx2_ASAP7_75t_L g4849 ( 
.A(n_4805),
.Y(n_4849)
);

OAI22xp5_ASAP7_75t_L g4850 ( 
.A1(n_4810),
.A2(n_3227),
.B1(n_3363),
.B2(n_3213),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4803),
.B(n_763),
.Y(n_4851)
);

AOI211xp5_ASAP7_75t_L g4852 ( 
.A1(n_4814),
.A2(n_768),
.B(n_766),
.C(n_767),
.Y(n_4852)
);

INVxp67_ASAP7_75t_L g4853 ( 
.A(n_4835),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4851),
.Y(n_4854)
);

AOI221xp5_ASAP7_75t_L g4855 ( 
.A1(n_4848),
.A2(n_4825),
.B1(n_4816),
.B2(n_3539),
.C(n_3551),
.Y(n_4855)
);

AOI221x1_ASAP7_75t_L g4856 ( 
.A1(n_4833),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.C(n_769),
.Y(n_4856)
);

AOI21xp5_ASAP7_75t_L g4857 ( 
.A1(n_4838),
.A2(n_770),
.B(n_771),
.Y(n_4857)
);

AOI221xp5_ASAP7_75t_L g4858 ( 
.A1(n_4839),
.A2(n_3539),
.B1(n_3551),
.B2(n_3499),
.C(n_3474),
.Y(n_4858)
);

NOR3xp33_ASAP7_75t_L g4859 ( 
.A(n_4840),
.B(n_771),
.C(n_772),
.Y(n_4859)
);

AOI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_4842),
.A2(n_3762),
.B1(n_3499),
.B2(n_3551),
.Y(n_4860)
);

HB1xp67_ASAP7_75t_L g4861 ( 
.A(n_4837),
.Y(n_4861)
);

OAI211xp5_ASAP7_75t_L g4862 ( 
.A1(n_4852),
.A2(n_775),
.B(n_773),
.C(n_774),
.Y(n_4862)
);

O2A1O1Ixp33_ASAP7_75t_L g4863 ( 
.A1(n_4843),
.A2(n_777),
.B(n_773),
.C(n_776),
.Y(n_4863)
);

O2A1O1Ixp33_ASAP7_75t_L g4864 ( 
.A1(n_4844),
.A2(n_779),
.B(n_776),
.C(n_778),
.Y(n_4864)
);

NOR3x1_ASAP7_75t_L g4865 ( 
.A(n_4830),
.B(n_778),
.C(n_780),
.Y(n_4865)
);

AOI211xp5_ASAP7_75t_L g4866 ( 
.A1(n_4846),
.A2(n_782),
.B(n_780),
.C(n_781),
.Y(n_4866)
);

AOI211xp5_ASAP7_75t_SL g4867 ( 
.A1(n_4845),
.A2(n_785),
.B(n_783),
.C(n_784),
.Y(n_4867)
);

OAI21xp5_ASAP7_75t_L g4868 ( 
.A1(n_4831),
.A2(n_4849),
.B(n_4836),
.Y(n_4868)
);

NAND3xp33_ASAP7_75t_L g4869 ( 
.A(n_4832),
.B(n_784),
.C(n_787),
.Y(n_4869)
);

OAI211xp5_ASAP7_75t_SL g4870 ( 
.A1(n_4834),
.A2(n_790),
.B(n_788),
.C(n_789),
.Y(n_4870)
);

AOI22xp5_ASAP7_75t_L g4871 ( 
.A1(n_4841),
.A2(n_3578),
.B1(n_3624),
.B2(n_3474),
.Y(n_4871)
);

AOI22xp5_ASAP7_75t_L g4872 ( 
.A1(n_4850),
.A2(n_3624),
.B1(n_3578),
.B2(n_3752),
.Y(n_4872)
);

NOR2xp33_ASAP7_75t_R g4873 ( 
.A(n_4847),
.B(n_788),
.Y(n_4873)
);

OAI21x1_ASAP7_75t_L g4874 ( 
.A1(n_4831),
.A2(n_790),
.B(n_791),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4867),
.B(n_791),
.Y(n_4875)
);

OAI211xp5_ASAP7_75t_L g4876 ( 
.A1(n_4873),
.A2(n_794),
.B(n_792),
.C(n_793),
.Y(n_4876)
);

NOR2xp33_ASAP7_75t_L g4877 ( 
.A(n_4853),
.B(n_792),
.Y(n_4877)
);

AND2x4_ASAP7_75t_L g4878 ( 
.A(n_4861),
.B(n_793),
.Y(n_4878)
);

BUFx6f_ASAP7_75t_L g4879 ( 
.A(n_4874),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4865),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4855),
.B(n_795),
.Y(n_4881)
);

INVxp67_ASAP7_75t_L g4882 ( 
.A(n_4869),
.Y(n_4882)
);

AOI22xp5_ASAP7_75t_L g4883 ( 
.A1(n_4859),
.A2(n_3624),
.B1(n_798),
.B2(n_796),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4856),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4863),
.Y(n_4885)
);

OAI22xp5_ASAP7_75t_SL g4886 ( 
.A1(n_4866),
.A2(n_799),
.B1(n_796),
.B2(n_797),
.Y(n_4886)
);

NOR2xp67_ASAP7_75t_L g4887 ( 
.A(n_4857),
.B(n_799),
.Y(n_4887)
);

INVx1_ASAP7_75t_SL g4888 ( 
.A(n_4854),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4860),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4864),
.Y(n_4890)
);

O2A1O1Ixp33_ASAP7_75t_L g4891 ( 
.A1(n_4881),
.A2(n_4868),
.B(n_4870),
.C(n_4862),
.Y(n_4891)
);

AND4x1_ASAP7_75t_L g4892 ( 
.A(n_4877),
.B(n_4858),
.C(n_4871),
.D(n_4872),
.Y(n_4892)
);

NOR3xp33_ASAP7_75t_L g4893 ( 
.A(n_4876),
.B(n_800),
.C(n_801),
.Y(n_4893)
);

OAI221xp5_ASAP7_75t_L g4894 ( 
.A1(n_4880),
.A2(n_803),
.B1(n_800),
.B2(n_802),
.C(n_804),
.Y(n_4894)
);

AND2x4_ASAP7_75t_L g4895 ( 
.A(n_4878),
.B(n_4889),
.Y(n_4895)
);

OAI321xp33_ASAP7_75t_L g4896 ( 
.A1(n_4885),
.A2(n_805),
.A3(n_806),
.B1(n_807),
.B2(n_808),
.C(n_809),
.Y(n_4896)
);

NOR2x1p5_ASAP7_75t_L g4897 ( 
.A(n_4875),
.B(n_807),
.Y(n_4897)
);

NOR3xp33_ASAP7_75t_L g4898 ( 
.A(n_4886),
.B(n_808),
.C(n_809),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4884),
.Y(n_4899)
);

NOR3xp33_ASAP7_75t_L g4900 ( 
.A(n_4888),
.B(n_810),
.C(n_811),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4887),
.B(n_810),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4899),
.Y(n_4902)
);

OA22x2_ASAP7_75t_L g4903 ( 
.A1(n_4895),
.A2(n_4883),
.B1(n_4890),
.B2(n_4882),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4901),
.Y(n_4904)
);

XNOR2xp5_ASAP7_75t_L g4905 ( 
.A(n_4892),
.B(n_4879),
.Y(n_4905)
);

INVx2_ASAP7_75t_L g4906 ( 
.A(n_4897),
.Y(n_4906)
);

BUFx3_ASAP7_75t_L g4907 ( 
.A(n_4894),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4905),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4902),
.Y(n_4909)
);

AOI22xp5_ASAP7_75t_L g4910 ( 
.A1(n_4903),
.A2(n_4893),
.B1(n_4898),
.B2(n_4900),
.Y(n_4910)
);

INVx2_ASAP7_75t_L g4911 ( 
.A(n_4906),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4908),
.B(n_4879),
.Y(n_4912)
);

OAI21x1_ASAP7_75t_SL g4913 ( 
.A1(n_4910),
.A2(n_4891),
.B(n_4904),
.Y(n_4913)
);

OAI22xp5_ASAP7_75t_L g4914 ( 
.A1(n_4909),
.A2(n_4907),
.B1(n_4896),
.B2(n_813),
.Y(n_4914)
);

OAI21xp5_ASAP7_75t_L g4915 ( 
.A1(n_4912),
.A2(n_4914),
.B(n_4911),
.Y(n_4915)
);

OAI22xp5_ASAP7_75t_L g4916 ( 
.A1(n_4913),
.A2(n_813),
.B1(n_811),
.B2(n_812),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4916),
.Y(n_4917)
);

AO22x2_ASAP7_75t_L g4918 ( 
.A1(n_4915),
.A2(n_816),
.B1(n_814),
.B2(n_815),
.Y(n_4918)
);

OA22x2_ASAP7_75t_SL g4919 ( 
.A1(n_4916),
.A2(n_818),
.B1(n_814),
.B2(n_817),
.Y(n_4919)
);

AOI22xp5_ASAP7_75t_L g4920 ( 
.A1(n_4917),
.A2(n_819),
.B1(n_817),
.B2(n_818),
.Y(n_4920)
);

AOI22xp33_ASAP7_75t_L g4921 ( 
.A1(n_4918),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.Y(n_4921)
);

XNOR2xp5_ASAP7_75t_L g4922 ( 
.A(n_4920),
.B(n_4919),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4921),
.B(n_820),
.Y(n_4923)
);

AOI22x1_ASAP7_75t_L g4924 ( 
.A1(n_4922),
.A2(n_4923),
.B1(n_823),
.B2(n_821),
.Y(n_4924)
);

XNOR2xp5_ASAP7_75t_L g4925 ( 
.A(n_4922),
.B(n_822),
.Y(n_4925)
);

AOI221xp5_ASAP7_75t_L g4926 ( 
.A1(n_4925),
.A2(n_825),
.B1(n_822),
.B2(n_824),
.C(n_826),
.Y(n_4926)
);

AOI211xp5_ASAP7_75t_L g4927 ( 
.A1(n_4926),
.A2(n_4924),
.B(n_827),
.C(n_824),
.Y(n_4927)
);


endmodule