module fake_jpeg_14345_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_21),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_35),
.B(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_14),
.B1(n_19),
.B2(n_16),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_43),
.B1(n_37),
.B2(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_14),
.B1(n_19),
.B2(n_16),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_27),
.B1(n_18),
.B2(n_14),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_19),
.B1(n_16),
.B2(n_14),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_65),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_43),
.B1(n_49),
.B2(n_46),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_22),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_26),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_76),
.B1(n_59),
.B2(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_18),
.B1(n_23),
.B2(n_50),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_51),
.A3(n_23),
.B1(n_17),
.B2(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_29),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_9),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_65),
.B1(n_57),
.B2(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_91),
.B1(n_95),
.B2(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_17),
.B1(n_44),
.B2(n_30),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_90),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_52),
.B1(n_60),
.B2(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_17),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_60),
.B(n_63),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_94),
.B(n_69),
.C(n_74),
.D(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_55),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_66),
.B1(n_63),
.B2(n_33),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_78),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_106),
.C(n_91),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.C(n_101),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_80),
.B(n_71),
.C(n_83),
.D(n_79),
.Y(n_100)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_80),
.B(n_71),
.C(n_79),
.D(n_30),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_105),
.B1(n_84),
.B2(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_86),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_44),
.C(n_1),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_87),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_114),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_89),
.B1(n_96),
.B2(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_111),
.B1(n_113),
.B2(n_106),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_99),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_84),
.B(n_96),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_101),
.B(n_100),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_112),
.A3(n_107),
.B1(n_44),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_110),
.C(n_114),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_123),
.C(n_11),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_5),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_12),
.Y(n_123)
);

OAI221xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_119),
.B1(n_116),
.B2(n_117),
.C(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

OAI221xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_2),
.B1(n_3),
.B2(n_9),
.C(n_10),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_127),
.B1(n_11),
.B2(n_0),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_0),
.C(n_130),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_0),
.Y(n_132)
);


endmodule