module real_aes_7326_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g189 ( .A1(n_0), .A2(n_190), .B(n_193), .C(n_197), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_1), .B(n_181), .Y(n_200) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_3), .B(n_191), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_4), .A2(n_154), .B(n_157), .C(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_5), .A2(n_149), .B(n_567), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_6), .A2(n_149), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_7), .B(n_181), .Y(n_573) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_8), .A2(n_183), .B(n_255), .Y(n_254) );
AND2x6_ASAP7_75t_L g154 ( .A(n_9), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_10), .A2(n_154), .B(n_157), .C(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g534 ( .A(n_11), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_12), .B(n_40), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_13), .B(n_196), .Y(n_545) );
INVx1_ASAP7_75t_L g175 ( .A(n_14), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_15), .B(n_191), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_16), .A2(n_192), .B(n_553), .C(n_555), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_17), .A2(n_105), .B1(n_118), .B2(n_767), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_18), .B(n_181), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_19), .B(n_169), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_20), .A2(n_157), .B(n_160), .C(n_168), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_21), .A2(n_195), .B(n_263), .C(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_22), .B(n_196), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_23), .B(n_196), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_24), .Y(n_515) );
INVx1_ASAP7_75t_L g495 ( .A(n_25), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_26), .A2(n_157), .B(n_168), .C(n_258), .Y(n_257) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_27), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_28), .Y(n_541) );
INVx1_ASAP7_75t_L g509 ( .A(n_29), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_30), .A2(n_149), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g152 ( .A(n_31), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_32), .A2(n_207), .B(n_208), .C(n_212), .Y(n_206) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_33), .A2(n_34), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_33), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_34), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_35), .A2(n_195), .B(n_570), .C(n_572), .Y(n_569) );
INVxp67_ASAP7_75t_L g510 ( .A(n_36), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_37), .B(n_260), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_38), .A2(n_157), .B(n_168), .C(n_494), .Y(n_493) );
CKINVDCx14_ASAP7_75t_R g568 ( .A(n_39), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_41), .A2(n_197), .B(n_532), .C(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_42), .B(n_148), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_43), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_44), .B(n_191), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_45), .B(n_149), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_46), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_47), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_48), .A2(n_207), .B(n_212), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g194 ( .A(n_49), .Y(n_194) );
INVx1_ASAP7_75t_L g238 ( .A(n_50), .Y(n_238) );
INVx1_ASAP7_75t_L g581 ( .A(n_51), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_52), .B(n_149), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_53), .Y(n_177) );
CKINVDCx14_ASAP7_75t_R g530 ( .A(n_54), .Y(n_530) );
AOI22xp5_ASAP7_75t_SL g467 ( .A1(n_55), .A2(n_114), .B1(n_468), .B2(n_764), .Y(n_467) );
INVx1_ASAP7_75t_L g155 ( .A(n_56), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_57), .B(n_149), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_58), .B(n_181), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_59), .A2(n_167), .B(n_223), .C(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g174 ( .A(n_60), .Y(n_174) );
INVx1_ASAP7_75t_SL g571 ( .A(n_61), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_62), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_63), .B(n_191), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_64), .B(n_181), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_65), .B(n_192), .Y(n_273) );
INVx1_ASAP7_75t_L g518 ( .A(n_66), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_67), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_68), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_69), .A2(n_157), .B(n_212), .C(n_221), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_70), .Y(n_247) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_72), .A2(n_149), .B(n_529), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_73), .A2(n_95), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_73), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_74), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_75), .A2(n_103), .B1(n_477), .B2(n_478), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_75), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_76), .A2(n_149), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_77), .A2(n_148), .B(n_505), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_78), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_79), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_79), .Y(n_474) );
INVx1_ASAP7_75t_L g551 ( .A(n_80), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_81), .B(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_82), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_83), .A2(n_149), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g554 ( .A(n_84), .Y(n_554) );
INVx2_ASAP7_75t_L g172 ( .A(n_85), .Y(n_172) );
INVx1_ASAP7_75t_L g544 ( .A(n_86), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_87), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_88), .B(n_196), .Y(n_274) );
INVx2_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
OR2x2_ASAP7_75t_L g461 ( .A(n_89), .B(n_114), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_90), .A2(n_157), .B(n_212), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_91), .B(n_149), .Y(n_205) );
INVx1_ASAP7_75t_L g209 ( .A(n_92), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_93), .B(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_L g250 ( .A(n_94), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_95), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_96), .A2(n_473), .B1(n_479), .B2(n_480), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_96), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_97), .B(n_183), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g222 ( .A(n_99), .Y(n_222) );
INVx1_ASAP7_75t_L g269 ( .A(n_100), .Y(n_269) );
INVx2_ASAP7_75t_L g584 ( .A(n_101), .Y(n_584) );
AND2x2_ASAP7_75t_L g240 ( .A(n_102), .B(n_171), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_103), .Y(n_477) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g768 ( .A(n_108), .Y(n_768) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_SL g764 ( .A(n_111), .Y(n_764) );
INVx3_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
NOR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx2_ASAP7_75t_L g469 ( .A(n_113), .Y(n_469) );
INVx1_ASAP7_75t_L g482 ( .A(n_113), .Y(n_482) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_466), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g766 ( .A(n_123), .Y(n_766) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_459), .B(n_462), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_128), .B(n_182), .Y(n_546) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B1(n_136), .B2(n_137), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_136), .A2(n_137), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_414), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_349), .Y(n_138) );
NAND4xp25_ASAP7_75t_SL g139 ( .A(n_140), .B(n_294), .C(n_318), .D(n_341), .Y(n_139) );
AOI221xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_231), .B1(n_265), .B2(n_278), .C(n_281), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_201), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_143), .A2(n_179), .B1(n_232), .B2(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_143), .B(n_202), .Y(n_352) );
AND2x2_ASAP7_75t_L g371 ( .A(n_143), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_143), .B(n_355), .Y(n_441) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_179), .Y(n_143) );
AND2x2_ASAP7_75t_L g309 ( .A(n_144), .B(n_202), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_144), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g332 ( .A(n_144), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g337 ( .A(n_144), .B(n_180), .Y(n_337) );
INVx2_ASAP7_75t_L g369 ( .A(n_144), .Y(n_369) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_144), .Y(n_413) );
AND2x2_ASAP7_75t_L g430 ( .A(n_144), .B(n_307), .Y(n_430) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g348 ( .A(n_145), .B(n_307), .Y(n_348) );
AND2x4_ASAP7_75t_L g362 ( .A(n_145), .B(n_179), .Y(n_362) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_145), .Y(n_366) );
AND2x2_ASAP7_75t_L g386 ( .A(n_145), .B(n_301), .Y(n_386) );
AND2x2_ASAP7_75t_L g436 ( .A(n_145), .B(n_203), .Y(n_436) );
AND2x2_ASAP7_75t_L g446 ( .A(n_145), .B(n_180), .Y(n_446) );
OR2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_176), .Y(n_145) );
AOI21xp5_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_156), .B(n_169), .Y(n_146) );
BUFx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g270 ( .A(n_150), .B(n_154), .Y(n_270) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx1_ASAP7_75t_L g264 ( .A(n_152), .Y(n_264) );
INVx1_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_153), .Y(n_163) );
INVx3_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
INVx1_ASAP7_75t_L g260 ( .A(n_153), .Y(n_260) );
BUFx3_ASAP7_75t_L g168 ( .A(n_154), .Y(n_168) );
INVx4_ASAP7_75t_SL g199 ( .A(n_154), .Y(n_199) );
INVx5_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx3_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_158), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_164), .B(n_166), .Y(n_160) );
INVx2_ASAP7_75t_L g165 ( .A(n_162), .Y(n_165) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx4_ASAP7_75t_L g224 ( .A(n_163), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_165), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_165), .A2(n_211), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_165), .A2(n_518), .B(n_519), .C(n_520), .Y(n_517) );
O2A1O1Ixp5_ASAP7_75t_L g543 ( .A1(n_165), .A2(n_520), .B(n_544), .C(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_166), .A2(n_191), .B(n_495), .C(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_167), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_170), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g178 ( .A(n_171), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_171), .A2(n_235), .B(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_171), .A2(n_270), .B(n_492), .C(n_493), .Y(n_491) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_171), .A2(n_528), .B(n_535), .Y(n_527) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_172), .B(n_173), .Y(n_171) );
AND2x2_ASAP7_75t_L g184 ( .A(n_172), .B(n_173), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_178), .A2(n_540), .B(n_546), .Y(n_539) );
AND2x2_ASAP7_75t_L g302 ( .A(n_179), .B(n_202), .Y(n_302) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_179), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_179), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g392 ( .A(n_179), .Y(n_392) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g280 ( .A(n_180), .B(n_217), .Y(n_280) );
AND2x2_ASAP7_75t_L g307 ( .A(n_180), .B(n_218), .Y(n_307) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_185), .B(n_200), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_182), .B(n_214), .Y(n_213) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_182), .A2(n_219), .B(n_229), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_182), .B(n_230), .Y(n_229) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_182), .A2(n_268), .B(n_275), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_182), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_182), .A2(n_514), .B(n_521), .Y(n_513) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_183), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_183), .A2(n_256), .B(n_257), .Y(n_255) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g277 ( .A(n_184), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_SL g186 ( .A1(n_187), .A2(n_188), .B(n_189), .C(n_199), .Y(n_186) );
INVx2_ASAP7_75t_L g207 ( .A(n_188), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_188), .A2(n_199), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_188), .A2(n_199), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_188), .A2(n_199), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_SL g550 ( .A1(n_188), .A2(n_199), .B(n_551), .C(n_552), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g567 ( .A1(n_188), .A2(n_199), .B(n_568), .C(n_569), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_SL g580 ( .A1(n_188), .A2(n_199), .B(n_581), .C(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_191), .B(n_250), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_191), .A2(n_224), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_192), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_195), .B(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g532 ( .A(n_196), .Y(n_532) );
INVx2_ASAP7_75t_L g520 ( .A(n_197), .Y(n_520) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_198), .Y(n_211) );
INVx1_ASAP7_75t_L g555 ( .A(n_198), .Y(n_555) );
INVx1_ASAP7_75t_L g212 ( .A(n_199), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_201), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_215), .Y(n_201) );
OR2x2_ASAP7_75t_L g333 ( .A(n_202), .B(n_216), .Y(n_333) );
AND2x2_ASAP7_75t_L g370 ( .A(n_202), .B(n_280), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_202), .B(n_301), .Y(n_381) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_202), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_202), .B(n_337), .Y(n_454) );
INVx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx2_ASAP7_75t_L g279 ( .A(n_203), .Y(n_279) );
AND2x2_ASAP7_75t_L g288 ( .A(n_203), .B(n_216), .Y(n_288) );
AND2x2_ASAP7_75t_L g404 ( .A(n_203), .B(n_299), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_203), .B(n_337), .Y(n_426) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_216), .Y(n_372) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_217), .Y(n_324) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g301 ( .A(n_218), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_228), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_225), .C(n_226), .Y(n_221) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_224), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_224), .B(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g572 ( .A(n_227), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_241), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_232), .B(n_314), .Y(n_433) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_233), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g285 ( .A(n_233), .B(n_286), .Y(n_285) );
INVx5_ASAP7_75t_SL g293 ( .A(n_233), .Y(n_293) );
OR2x2_ASAP7_75t_L g316 ( .A(n_233), .B(n_286), .Y(n_316) );
OR2x2_ASAP7_75t_L g326 ( .A(n_233), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g389 ( .A(n_233), .B(n_243), .Y(n_389) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_233), .B(n_242), .Y(n_427) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_233), .B(n_369), .C(n_449), .D(n_450), .Y(n_448) );
AND2x2_ASAP7_75t_L g458 ( .A(n_233), .B(n_290), .Y(n_458) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g283 ( .A(n_242), .B(n_279), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_242), .B(n_285), .Y(n_452) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
OR2x2_ASAP7_75t_L g292 ( .A(n_243), .B(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g299 ( .A(n_243), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_243), .B(n_267), .Y(n_311) );
INVxp67_ASAP7_75t_L g314 ( .A(n_243), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_243), .B(n_286), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_243), .B(n_253), .Y(n_380) );
AND2x2_ASAP7_75t_L g395 ( .A(n_243), .B(n_290), .Y(n_395) );
OR2x2_ASAP7_75t_L g424 ( .A(n_243), .B(n_253), .Y(n_424) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_251), .Y(n_243) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_244), .A2(n_549), .B(n_556), .Y(n_548) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_244), .A2(n_566), .B(n_573), .Y(n_565) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_244), .A2(n_579), .B(n_585), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_252), .B(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_252), .B(n_293), .Y(n_432) );
OR2x2_ASAP7_75t_L g453 ( .A(n_252), .B(n_330), .Y(n_453) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g266 ( .A(n_253), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g290 ( .A(n_253), .B(n_286), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_253), .B(n_267), .Y(n_305) );
AND2x2_ASAP7_75t_L g375 ( .A(n_253), .B(n_299), .Y(n_375) );
AND2x2_ASAP7_75t_L g409 ( .A(n_253), .B(n_293), .Y(n_409) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_254), .B(n_293), .Y(n_312) );
AND2x2_ASAP7_75t_L g340 ( .A(n_254), .B(n_267), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_261), .B(n_262), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_262), .A2(n_273), .B(n_274), .Y(n_272) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_265), .B(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_266), .A2(n_355), .B1(n_391), .B2(n_408), .C(n_410), .Y(n_407) );
INVx5_ASAP7_75t_SL g286 ( .A(n_267), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_271), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_270), .A2(n_515), .B(n_516), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_270), .A2(n_541), .B(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g503 ( .A(n_277), .Y(n_503) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OAI33xp33_ASAP7_75t_L g306 ( .A1(n_279), .A2(n_307), .A3(n_308), .B1(n_310), .B2(n_313), .B3(n_317), .Y(n_306) );
OR2x2_ASAP7_75t_L g322 ( .A(n_279), .B(n_323), .Y(n_322) );
AOI322xp5_ASAP7_75t_L g431 ( .A1(n_279), .A2(n_348), .A3(n_355), .B1(n_432), .B2(n_433), .C1(n_434), .C2(n_437), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_279), .B(n_307), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_SL g455 ( .A1(n_279), .A2(n_307), .B(n_456), .C(n_458), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_280), .A2(n_295), .B1(n_300), .B2(n_303), .C(n_306), .Y(n_294) );
INVx1_ASAP7_75t_L g387 ( .A(n_280), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_280), .B(n_436), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B1(n_287), .B2(n_289), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g364 ( .A(n_285), .B(n_299), .Y(n_364) );
AND2x2_ASAP7_75t_L g422 ( .A(n_285), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g330 ( .A(n_286), .B(n_293), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_286), .B(n_299), .Y(n_358) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_288), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_288), .B(n_366), .Y(n_420) );
OAI321xp33_ASAP7_75t_L g439 ( .A1(n_288), .A2(n_361), .A3(n_440), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g406 ( .A(n_289), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_290), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g345 ( .A(n_290), .B(n_293), .Y(n_345) );
AOI321xp33_ASAP7_75t_L g403 ( .A1(n_290), .A2(n_307), .A3(n_404), .B1(n_405), .B2(n_406), .C(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g320 ( .A(n_292), .B(n_305), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_293), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_293), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_293), .B(n_379), .Y(n_416) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g339 ( .A(n_297), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g304 ( .A(n_298), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g412 ( .A(n_299), .Y(n_412) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_302), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g335 ( .A(n_307), .Y(n_335) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_309), .B(n_344), .Y(n_393) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
OR2x2_ASAP7_75t_L g357 ( .A(n_312), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g402 ( .A(n_312), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_313), .A2(n_360), .B1(n_363), .B2(n_365), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g457 ( .A(n_316), .B(n_380), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B1(n_325), .B2(n_331), .C(n_334), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_SL g401 ( .A(n_327), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_329), .B(n_379), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_329), .A2(n_397), .B(n_399), .Y(n_396) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g442 ( .A(n_330), .B(n_424), .Y(n_442) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_SL g344 ( .A(n_333), .Y(n_344) );
AOI21xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B(n_338), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g450 ( .A(n_340), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_344), .B(n_362), .Y(n_398) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g419 ( .A(n_348), .Y(n_419) );
NAND5xp2_ASAP7_75t_L g349 ( .A(n_350), .B(n_367), .C(n_376), .D(n_396), .E(n_403), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B(n_356), .C(n_359), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_363), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g405 ( .A(n_365), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_371), .B(n_373), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_368), .A2(n_422), .B1(n_425), .B2(n_427), .C(n_428), .Y(n_421) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
AOI321xp33_ASAP7_75t_L g376 ( .A1(n_369), .A2(n_377), .A3(n_381), .B1(n_382), .B2(n_388), .C(n_390), .Y(n_376) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g447 ( .A(n_381), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_383), .B(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g399 ( .A(n_384), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
NOR2xp67_ASAP7_75t_SL g411 ( .A(n_385), .B(n_392), .Y(n_411) );
AOI321xp33_ASAP7_75t_SL g443 ( .A1(n_388), .A2(n_444), .A3(n_445), .B1(n_446), .B2(n_447), .C(n_448), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_393), .C(n_394), .Y(n_390) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_401), .B(n_409), .Y(n_438) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .C(n_413), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_439), .C(n_451), .Y(n_414) );
OAI211xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_417), .B(n_421), .C(n_431), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_420), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_420), .A2(n_452), .B1(n_453), .B2(n_454), .C(n_455), .Y(n_451) );
INVx1_ASAP7_75t_L g440 ( .A(n_422), .Y(n_440) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g444 ( .A(n_442), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx14_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g465 ( .A(n_461), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_462), .A2(n_467), .B(n_765), .Y(n_466) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B1(n_481), .B2(n_483), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_471), .A2(n_472), .B1(n_484), .B2(n_485), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_473), .Y(n_480) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR4x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_654), .C(n_701), .D(n_741), .Y(n_485) );
NAND3xp33_ASAP7_75t_SL g486 ( .A(n_487), .B(n_600), .C(n_629), .Y(n_486) );
AOI211xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_523), .B(n_557), .C(n_593), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_488), .A2(n_613), .B(n_630), .C(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_490), .B(n_592), .Y(n_591) );
INVx3_ASAP7_75t_SL g596 ( .A(n_490), .Y(n_596) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_490), .Y(n_608) );
AND2x4_ASAP7_75t_L g612 ( .A(n_490), .B(n_564), .Y(n_612) );
AND2x2_ASAP7_75t_L g623 ( .A(n_490), .B(n_513), .Y(n_623) );
OR2x2_ASAP7_75t_L g647 ( .A(n_490), .B(n_560), .Y(n_647) );
AND2x2_ASAP7_75t_L g660 ( .A(n_490), .B(n_565), .Y(n_660) );
AND2x2_ASAP7_75t_L g700 ( .A(n_490), .B(n_686), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_490), .B(n_670), .Y(n_707) );
AND2x2_ASAP7_75t_L g737 ( .A(n_490), .B(n_500), .Y(n_737) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_497), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_499), .B(n_664), .Y(n_676) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_512), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_500), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g614 ( .A(n_500), .B(n_512), .Y(n_614) );
BUFx3_ASAP7_75t_L g622 ( .A(n_500), .Y(n_622) );
OR2x2_ASAP7_75t_L g643 ( .A(n_500), .B(n_526), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_500), .B(n_664), .Y(n_754) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .B(n_511), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g561 ( .A(n_504), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_512), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g607 ( .A(n_512), .Y(n_607) );
AND2x2_ASAP7_75t_L g670 ( .A(n_512), .B(n_565), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_512), .A2(n_673), .B1(n_675), .B2(n_677), .C(n_678), .Y(n_672) );
AND2x2_ASAP7_75t_L g686 ( .A(n_512), .B(n_560), .Y(n_686) );
AND2x2_ASAP7_75t_L g712 ( .A(n_512), .B(n_596), .Y(n_712) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g592 ( .A(n_513), .B(n_565), .Y(n_592) );
BUFx2_ASAP7_75t_L g726 ( .A(n_513), .Y(n_726) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI32xp33_ASAP7_75t_L g692 ( .A1(n_524), .A2(n_653), .A3(n_667), .B1(n_693), .B2(n_694), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .Y(n_524) );
AND2x2_ASAP7_75t_L g633 ( .A(n_525), .B(n_577), .Y(n_633) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g615 ( .A(n_526), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_526), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g687 ( .A(n_526), .B(n_577), .Y(n_687) );
AND2x2_ASAP7_75t_L g698 ( .A(n_526), .B(n_590), .Y(n_698) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g599 ( .A(n_527), .B(n_578), .Y(n_599) );
AND2x2_ASAP7_75t_L g603 ( .A(n_527), .B(n_578), .Y(n_603) );
AND2x2_ASAP7_75t_L g638 ( .A(n_527), .B(n_589), .Y(n_638) );
AND2x2_ASAP7_75t_L g645 ( .A(n_527), .B(n_547), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_527), .A2(n_596), .B(n_607), .C(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g704 ( .A(n_527), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_527), .B(n_538), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_536), .B(n_587), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_536), .B(n_603), .Y(n_693) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g598 ( .A(n_537), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
AND2x2_ASAP7_75t_L g590 ( .A(n_538), .B(n_548), .Y(n_590) );
OR2x2_ASAP7_75t_L g605 ( .A(n_538), .B(n_548), .Y(n_605) );
AND2x2_ASAP7_75t_L g628 ( .A(n_538), .B(n_589), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_538), .Y(n_632) );
AND2x2_ASAP7_75t_L g651 ( .A(n_538), .B(n_588), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_538), .A2(n_616), .B1(n_662), .B2(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_538), .B(n_704), .Y(n_728) );
AND2x2_ASAP7_75t_L g743 ( .A(n_538), .B(n_603), .Y(n_743) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g575 ( .A(n_539), .Y(n_575) );
AND2x2_ASAP7_75t_L g617 ( .A(n_539), .B(n_548), .Y(n_617) );
AND2x2_ASAP7_75t_L g619 ( .A(n_539), .B(n_577), .Y(n_619) );
AND3x2_ASAP7_75t_L g681 ( .A(n_539), .B(n_645), .C(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g716 ( .A(n_547), .B(n_588), .Y(n_716) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g577 ( .A(n_548), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_548), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_548), .B(n_587), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_548), .B(n_628), .C(n_704), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_574), .B1(n_586), .B2(n_591), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_560), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g668 ( .A(n_560), .Y(n_668) );
OAI31xp33_ASAP7_75t_L g684 ( .A1(n_563), .A2(n_685), .A3(n_686), .B(n_687), .Y(n_684) );
AND2x2_ASAP7_75t_L g709 ( .A(n_563), .B(n_596), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_563), .B(n_622), .Y(n_755) );
AND2x2_ASAP7_75t_L g664 ( .A(n_564), .B(n_596), .Y(n_664) );
AND2x2_ASAP7_75t_L g725 ( .A(n_564), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g595 ( .A(n_565), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
CKINVDCx16_ASAP7_75t_R g674 ( .A(n_575), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_576), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AOI221x1_ASAP7_75t_SL g641 ( .A1(n_577), .A2(n_642), .B1(n_644), .B2(n_646), .C(n_648), .Y(n_641) );
INVx2_ASAP7_75t_L g589 ( .A(n_578), .Y(n_589) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_578), .Y(n_683) );
INVx1_ASAP7_75t_L g671 ( .A(n_586), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_587), .B(n_604), .Y(n_696) );
INVx1_ASAP7_75t_SL g759 ( .A(n_587), .Y(n_759) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g677 ( .A(n_590), .B(n_603), .Y(n_677) );
INVx1_ASAP7_75t_L g745 ( .A(n_591), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_591), .B(n_674), .Y(n_758) );
INVx2_ASAP7_75t_SL g597 ( .A(n_592), .Y(n_597) );
AND2x2_ASAP7_75t_L g640 ( .A(n_592), .B(n_596), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_592), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_592), .B(n_667), .Y(n_694) );
AOI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_597), .B(n_598), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_595), .B(n_667), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_595), .B(n_622), .Y(n_763) );
OR2x2_ASAP7_75t_L g635 ( .A(n_596), .B(n_614), .Y(n_635) );
AND2x2_ASAP7_75t_L g734 ( .A(n_596), .B(n_725), .Y(n_734) );
OAI22xp5_ASAP7_75t_SL g609 ( .A1(n_597), .A2(n_610), .B1(n_615), .B2(n_618), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_597), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g657 ( .A(n_599), .B(n_605), .Y(n_657) );
INVx1_ASAP7_75t_L g721 ( .A(n_599), .Y(n_721) );
AOI311xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_606), .A3(n_608), .B(n_609), .C(n_620), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_604), .A2(n_736), .B1(n_748), .B2(n_751), .C(n_753), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_604), .B(n_759), .Y(n_761) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g658 ( .A(n_606), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_607), .A2(n_649), .B(n_650), .C(n_652), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_SL g717 ( .A1(n_611), .A2(n_613), .B(n_718), .C(n_719), .Y(n_717) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_612), .B(n_686), .Y(n_752) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_615), .A2(n_635), .B1(n_636), .B2(n_639), .C(n_641), .Y(n_634) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g637 ( .A(n_617), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g720 ( .A(n_617), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_621), .A2(n_679), .B(n_680), .C(n_684), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_622), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_622), .B(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g644 ( .A(n_628), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_632), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g746 ( .A(n_635), .Y(n_746) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_638), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g673 ( .A(n_638), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g750 ( .A(n_638), .Y(n_750) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g691 ( .A(n_640), .B(n_667), .Y(n_691) );
INVx1_ASAP7_75t_SL g685 ( .A(n_647), .Y(n_685) );
INVx1_ASAP7_75t_L g662 ( .A(n_653), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_672), .C(n_688), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .A3(n_659), .B1(n_661), .B2(n_665), .C1(n_669), .C2(n_671), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g708 ( .A1(n_656), .A2(n_709), .B(n_710), .C(n_717), .Y(n_708) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_659), .A2(n_680), .B1(n_711), .B2(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g669 ( .A(n_667), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g706 ( .A(n_667), .B(n_707), .Y(n_706) );
AOI32xp33_ASAP7_75t_L g757 ( .A1(n_667), .A2(n_758), .A3(n_759), .B1(n_760), .B2(n_762), .Y(n_757) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g679 ( .A(n_670), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_670), .A2(n_723), .B1(n_727), .B2(n_729), .C(n_732), .Y(n_722) );
AND2x2_ASAP7_75t_L g736 ( .A(n_670), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g739 ( .A(n_674), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g749 ( .A(n_674), .B(n_750), .Y(n_749) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g740 ( .A(n_683), .B(n_704), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_692), .C(n_695), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI211xp5_ASAP7_75t_SL g701 ( .A1(n_702), .A2(n_705), .B(n_708), .C(n_722), .Y(n_701) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_716), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g731 ( .A(n_728), .Y(n_731) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B(n_738), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_744), .B(n_747), .C(n_757), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
endmodule