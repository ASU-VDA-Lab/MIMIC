module fake_jpeg_501_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_16),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_58),
.Y(n_66)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_45),
.B(n_47),
.Y(n_62)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_53),
.B(n_48),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_67),
.B(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_78),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_38),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_85),
.Y(n_88)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_38),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_4),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_50),
.B1(n_44),
.B2(n_52),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_61),
.B1(n_52),
.B2(n_50),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_85),
.B1(n_79),
.B2(n_75),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_61),
.B1(n_1),
.B2(n_2),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_0),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_98),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_21),
.Y(n_106)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_20),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_111),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_5),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_110),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_117),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_6),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_116),
.B1(n_11),
.B2(n_12),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_96),
.B(n_27),
.C(n_28),
.D(n_36),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_125),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_130),
.B1(n_103),
.B2(n_102),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_11),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_23),
.C(n_34),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_103),
.C(n_31),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_13),
.B(n_14),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_22),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_127),
.B1(n_121),
.B2(n_125),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_35),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_140),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_135),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_138),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_141),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_133),
.C(n_139),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_119),
.B(n_118),
.C(n_124),
.D(n_134),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_126),
.B(n_122),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_29),
.Y(n_149)
);


endmodule