module fake_jpeg_7112_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_42),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_51),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_19),
.B1(n_33),
.B2(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_58),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_19),
.B1(n_21),
.B2(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_19),
.B1(n_20),
.B2(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_19),
.B1(n_33),
.B2(n_28),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_25),
.C(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_34),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_30),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_78),
.C(n_84),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_72),
.Y(n_104)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_80),
.Y(n_107)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_76),
.B1(n_28),
.B2(n_65),
.Y(n_116)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_83),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_92),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_16),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_65),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_45),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_110),
.B(n_99),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_48),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_108),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_34),
.CON(n_110),
.SN(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_117),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_68),
.B1(n_55),
.B2(n_33),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_86),
.B1(n_85),
.B2(n_81),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_60),
.C(n_45),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_119),
.C(n_17),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_122),
.B1(n_73),
.B2(n_72),
.Y(n_147)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_89),
.C(n_69),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_23),
.C(n_30),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_128),
.B1(n_17),
.B2(n_27),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_31),
.B1(n_23),
.B2(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_129),
.B(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_142),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_143),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_20),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_135),
.A2(n_115),
.B(n_125),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_145),
.B(n_120),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_82),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_144),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_124),
.B1(n_106),
.B2(n_126),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_34),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_16),
.B(n_27),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_86),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_34),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_34),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_27),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_0),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_159),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_76),
.B1(n_75),
.B2(n_23),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_154),
.A2(n_24),
.B1(n_120),
.B2(n_32),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_107),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_102),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_71),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_0),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_169),
.B(n_175),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_106),
.B1(n_126),
.B2(n_123),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_170),
.B1(n_173),
.B2(n_191),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_120),
.C(n_21),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_183),
.C(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_20),
.B(n_24),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_22),
.B1(n_18),
.B2(n_32),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_18),
.B(n_22),
.C(n_2),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_177),
.B(n_157),
.Y(n_194)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_142),
.C(n_148),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_102),
.C(n_22),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_131),
.B1(n_154),
.B2(n_143),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_18),
.B(n_22),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_188),
.B(n_138),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_18),
.B(n_22),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_18),
.B1(n_32),
.B2(n_102),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_135),
.B(n_7),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_140),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_129),
.Y(n_197)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_139),
.A3(n_145),
.B1(n_152),
.B2(n_136),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_210),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_179),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_209),
.B1(n_214),
.B2(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_136),
.B1(n_130),
.B2(n_156),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_175),
.B1(n_186),
.B2(n_190),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_207),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_130),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_192),
.C(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_211),
.A2(n_212),
.B(n_213),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_155),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_9),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_220),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_2),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_2),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_222),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_3),
.B(n_4),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_167),
.B(n_183),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_231),
.C(n_235),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_166),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_244),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_201),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_172),
.C(n_169),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_188),
.B1(n_173),
.B2(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_212),
.B(n_197),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_211),
.B(n_219),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_162),
.C(n_176),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_180),
.C(n_175),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_175),
.C(n_4),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_3),
.C(n_5),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_205),
.C(n_203),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_246),
.C(n_247),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_199),
.A2(n_3),
.B1(n_15),
.B2(n_8),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_213),
.B1(n_207),
.B2(n_216),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_6),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_6),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_198),
.B(n_6),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_223),
.B(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_248),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_214),
.B(n_199),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_264),
.B(n_209),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_201),
.Y(n_282)
);

AOI221xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_220),
.B1(n_244),
.B2(n_242),
.C(n_246),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_240),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_231),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_273),
.Y(n_291)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_242),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_286),
.B(n_262),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_226),
.C(n_206),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_254),
.C(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_250),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_253),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_280),
.A2(n_259),
.B1(n_263),
.B2(n_257),
.Y(n_289)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_271),
.B(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_297),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_269),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_301),
.C(n_302),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_270),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_261),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_287),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_261),
.B(n_258),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_258),
.C(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_284),
.B1(n_251),
.B2(n_286),
.Y(n_303)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_298),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_306),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_295),
.B(n_291),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_292),
.A2(n_278),
.B(n_281),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_SL g315 ( 
.A(n_312),
.B(n_302),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_287),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_291),
.C(n_9),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_316),
.Y(n_330)
);

AOI21x1_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_307),
.B(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_310),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_319),
.C(n_322),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_311),
.B(n_309),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_8),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_10),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_9),
.C(n_10),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_329),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_314),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_328),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_310),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_15),
.Y(n_329)
);

AOI321xp33_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_330),
.A3(n_327),
.B1(n_324),
.B2(n_14),
.C(n_13),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_331),
.B(n_333),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_10),
.C(n_12),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_12),
.Y(n_338)
);


endmodule