module fake_netlist_5_1177_n_1778 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1778);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1778;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_85),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_16),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_119),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_56),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_32),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_81),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_18),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_125),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_98),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_99),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_65),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_41),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_61),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_40),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_49),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_41),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_115),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_25),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_14),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_63),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_66),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_74),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_54),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_149),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_145),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_25),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_0),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_48),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_14),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_42),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_150),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_169),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_111),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_127),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_164),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_129),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_50),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_64),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_140),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_87),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_11),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_116),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_75),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_23),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_96),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_10),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_77),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_4),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_58),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_95),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_126),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_102),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_80),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_104),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_34),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_83),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_38),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_27),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_28),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_20),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_142),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_34),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_152),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_97),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_123),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_73),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_92),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_110),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_89),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_68),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_23),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_171),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_54),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_118),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_71),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_107),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_165),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_22),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_162),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_100),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_161),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_144),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_141),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_93),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_132),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_160),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_91),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_21),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_120),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_46),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_135),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_19),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_117),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_42),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_16),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_33),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_40),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_57),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_19),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_69),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_109),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_31),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_67),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_1),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_167),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_90),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_174),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_148),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_170),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_3),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_2),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_94),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_39),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_17),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_131),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_153),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_29),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_35),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_15),
.Y(n_330)
);

BUFx8_ASAP7_75t_SL g331 ( 
.A(n_8),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_30),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_22),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_62),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_52),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_7),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_137),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_21),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_10),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_36),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_155),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_105),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_173),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_35),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_124),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_53),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_52),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_31),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_39),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_59),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_3),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_45),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_82),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_38),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_220),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_185),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_220),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_220),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_205),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_185),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_220),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_195),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_331),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_197),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_256),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_178),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_210),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_246),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_269),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_311),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_181),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_184),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_182),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_182),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_219),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_192),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_244),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_193),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_195),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_288),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_188),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_276),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_219),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_189),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_288),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_242),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_242),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_293),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_249),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_249),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_260),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_179),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_260),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_345),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_261),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_261),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_194),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_268),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_276),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_239),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_196),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_239),
.Y(n_412)
);

INVxp33_ASAP7_75t_SL g413 ( 
.A(n_191),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_268),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_202),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_199),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_315),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_280),
.Y(n_418)
);

BUFx2_ASAP7_75t_SL g419 ( 
.A(n_183),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_267),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_280),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_179),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_276),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_297),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_206),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_297),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_200),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_201),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_214),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_215),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_345),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_299),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_239),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_299),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_300),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_300),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_316),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_325),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_221),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_229),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_325),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_328),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_328),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_183),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_355),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_367),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_222),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_374),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_430),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_398),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_263),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_372),
.B(n_222),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_356),
.B(n_267),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_L g459 ( 
.A(n_402),
.B(n_263),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_361),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_361),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_389),
.B(n_275),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_380),
.B(n_275),
.Y(n_463)
);

CKINVDCx8_ASAP7_75t_R g464 ( 
.A(n_410),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_386),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_363),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_363),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_422),
.Y(n_469)
);

BUFx8_ASAP7_75t_L g470 ( 
.A(n_366),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_360),
.A2(n_247),
.B1(n_354),
.B2(n_294),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_362),
.B(n_296),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_422),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_383),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_368),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_364),
.B(n_319),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_390),
.B(n_319),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_368),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_388),
.B(n_207),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_383),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_384),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_395),
.B(n_296),
.Y(n_482)
);

BUFx8_ASAP7_75t_L g483 ( 
.A(n_366),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_404),
.B(n_207),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_369),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_431),
.B(n_243),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_407),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_411),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_410),
.B(n_316),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_385),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_416),
.B(n_243),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_385),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_412),
.A2(n_245),
.B1(n_227),
.B2(n_226),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_415),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_420),
.B(n_251),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_396),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_R g501 ( 
.A(n_427),
.B(n_230),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_375),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_425),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_394),
.B(n_413),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_428),
.B(n_251),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_397),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_399),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_412),
.B(n_316),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_429),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_433),
.A2(n_305),
.B1(n_320),
.B2(n_332),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_433),
.A2(n_324),
.B1(n_258),
.B2(n_349),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_439),
.B(n_321),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_420),
.B(n_321),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_440),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_419),
.B(n_252),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_370),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_400),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_455),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_449),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

AND3x2_ASAP7_75t_L g524 ( 
.A(n_465),
.B(n_248),
.C(n_357),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_449),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_476),
.B(n_477),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_446),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_512),
.A2(n_377),
.B1(n_417),
.B2(n_379),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_469),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_451),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_476),
.B(n_419),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_494),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_458),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_461),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_476),
.B(n_477),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_494),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_491),
.A2(n_387),
.B1(n_426),
.B2(n_208),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_472),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_477),
.A2(n_329),
.B1(n_333),
.B2(n_335),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_472),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_469),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_454),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_479),
.B(n_437),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_487),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_506),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_482),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_506),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_506),
.Y(n_550)
);

OAI21xp33_ASAP7_75t_SL g551 ( 
.A1(n_491),
.A2(n_333),
.B(n_329),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_505),
.B(n_387),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_461),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_493),
.B(n_437),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_469),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_482),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_446),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_473),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_453),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_473),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_444),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_501),
.B(n_365),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_454),
.Y(n_565)
);

INVx8_ASAP7_75t_L g566 ( 
.A(n_484),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_510),
.B(n_392),
.Y(n_567)
);

INVxp33_ASAP7_75t_L g568 ( 
.A(n_497),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_464),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_451),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_473),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_445),
.A2(n_187),
.B(n_186),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_451),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_453),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_464),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_506),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_507),
.B(n_180),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_508),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_L g582 ( 
.A(n_457),
.B(n_217),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_450),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_463),
.B(n_217),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_514),
.B(n_186),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_510),
.A2(n_277),
.B1(n_312),
.B2(n_307),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_509),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_484),
.B(n_231),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_452),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_509),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_484),
.B(n_486),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_466),
.B(n_409),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_486),
.B(n_232),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_460),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_466),
.B(n_423),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_467),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_509),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_517),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_517),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_517),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_486),
.B(n_234),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_520),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_471),
.A2(n_283),
.B1(n_274),
.B2(n_309),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_488),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_470),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_520),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_518),
.A2(n_190),
.B(n_187),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_504),
.A2(n_259),
.B1(n_237),
.B2(n_314),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_488),
.A2(n_330),
.B1(n_348),
.B2(n_347),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_520),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_520),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_444),
.A2(n_335),
.B1(n_339),
.B2(n_351),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_474),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_475),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_475),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_478),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_481),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_489),
.Y(n_624)
);

AND3x2_ASAP7_75t_L g625 ( 
.A(n_444),
.B(n_198),
.C(n_190),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_470),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_503),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_478),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_492),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_496),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_448),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_448),
.B(n_235),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_485),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_500),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_490),
.B(n_236),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_502),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_448),
.B(n_198),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_490),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_462),
.B(n_203),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_462),
.A2(n_339),
.B1(n_351),
.B2(n_352),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_511),
.B(n_240),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_499),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_519),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_519),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_498),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_456),
.B(n_204),
.C(n_203),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_462),
.A2(n_352),
.B1(n_337),
.B2(n_216),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_498),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_498),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_515),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_515),
.B(n_241),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_SL g654 ( 
.A1(n_470),
.A2(n_322),
.B1(n_211),
.B2(n_212),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_515),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_459),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_459),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_511),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_495),
.Y(n_659)
);

BUFx4f_ASAP7_75t_L g660 ( 
.A(n_516),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_483),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_483),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_513),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_503),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_483),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_505),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_449),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_469),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_458),
.B(n_370),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_449),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_655),
.B(n_204),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_655),
.B(n_209),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_655),
.B(n_209),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_629),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_618),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_534),
.B(n_217),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_629),
.Y(n_678)
);

AO22x2_ASAP7_75t_L g679 ( 
.A1(n_659),
.A2(n_213),
.B1(n_216),
.B2(n_233),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_527),
.A2(n_342),
.B1(n_213),
.B2(n_233),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_521),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_618),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_562),
.B(n_238),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_629),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_562),
.B(n_632),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_534),
.B(n_322),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_632),
.B(n_238),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_522),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_537),
.B(n_253),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_623),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_656),
.B(n_253),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_656),
.B(n_271),
.Y(n_692)
);

O2A1O1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_612),
.A2(n_271),
.B(n_342),
.C(n_337),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_620),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_657),
.B(n_278),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_540),
.A2(n_270),
.B1(n_353),
.B2(n_350),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_623),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_624),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_540),
.A2(n_291),
.B1(n_327),
.B2(n_278),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_657),
.B(n_593),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_566),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_548),
.B(n_217),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_548),
.B(n_322),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_647),
.B(n_282),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_546),
.B(n_250),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_535),
.B(n_400),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_647),
.B(n_282),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_535),
.B(n_218),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_661),
.B(n_284),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_624),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_521),
.B(n_528),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_542),
.B(n_217),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_659),
.A2(n_664),
.B1(n_542),
.B2(n_557),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_650),
.B(n_284),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_630),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_651),
.B(n_308),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_575),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_525),
.Y(n_718)
);

BUFx5_ASAP7_75t_L g719 ( 
.A(n_523),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_536),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_651),
.B(n_308),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_652),
.B(n_326),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_557),
.B(n_272),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_532),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_670),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_566),
.B(n_327),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_566),
.B(n_334),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_553),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_658),
.B(n_254),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_631),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_566),
.B(n_334),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_R g732 ( 
.A(n_569),
.B(n_255),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_670),
.B(n_401),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_664),
.A2(n_257),
.B1(n_262),
.B2(n_264),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_578),
.B(n_265),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_558),
.B(n_401),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_619),
.B(n_266),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_658),
.B(n_403),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_619),
.B(n_273),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_638),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_560),
.B(n_403),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_619),
.B(n_279),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_590),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_619),
.B(n_281),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_619),
.B(n_285),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_635),
.B(n_286),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_545),
.B(n_287),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_620),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_L g749 ( 
.A1(n_573),
.A2(n_443),
.B(n_442),
.C(n_441),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_554),
.B(n_223),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_635),
.B(n_289),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_635),
.B(n_290),
.Y(n_752)
);

AO22x2_ASAP7_75t_L g753 ( 
.A1(n_648),
.A2(n_443),
.B1(n_442),
.B2(n_441),
.Y(n_753)
);

INVxp33_ASAP7_75t_L g754 ( 
.A(n_568),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_579),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_621),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_625),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_638),
.B(n_405),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_584),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_553),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_635),
.B(n_292),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_539),
.B(n_224),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_627),
.B(n_405),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_668),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_595),
.B(n_225),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_581),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_635),
.B(n_295),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_637),
.B(n_298),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_555),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_658),
.B(n_302),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_606),
.B(n_228),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_586),
.B(n_301),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_551),
.A2(n_438),
.B(n_436),
.C(n_435),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_555),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_591),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_637),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_551),
.B(n_438),
.C(n_436),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_556),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_663),
.B(n_406),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_637),
.B(n_310),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_591),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_638),
.B(n_406),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_586),
.A2(n_435),
.B1(n_434),
.B2(n_432),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_663),
.B(n_408),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_637),
.B(n_313),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_596),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_637),
.B(n_317),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_586),
.B(n_304),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_600),
.B(n_318),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_653),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_596),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_523),
.B(n_323),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_614),
.B(n_434),
.C(n_432),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_526),
.B(n_341),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_541),
.A2(n_424),
.B(n_421),
.C(n_418),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_621),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_586),
.A2(n_633),
.B1(n_552),
.B2(n_640),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_533),
.B(n_343),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_538),
.B(n_421),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_602),
.B(n_340),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_538),
.B(n_418),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_547),
.B(n_414),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_547),
.B(n_414),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_586),
.A2(n_408),
.B1(n_344),
.B2(n_346),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_598),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_622),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_598),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_549),
.B(n_550),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_588),
.B(n_0),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_599),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_599),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_550),
.B(n_381),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_622),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_588),
.B(n_636),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_628),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_665),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_661),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_602),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_613),
.B(n_378),
.C(n_376),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_580),
.B(n_378),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_649),
.A2(n_373),
.B1(n_371),
.B2(n_376),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_643),
.B(n_5),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_628),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_668),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_638),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_556),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_634),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_700),
.B(n_641),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_740),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_694),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_740),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_755),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_815),
.B(n_660),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_759),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_724),
.B(n_641),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_780),
.B(n_609),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_815),
.B(n_660),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_819),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_761),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_738),
.B(n_660),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_776),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_725),
.B(n_609),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_810),
.A2(n_638),
.B1(n_640),
.B2(n_583),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_685),
.A2(n_589),
.B(n_577),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_694),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_743),
.B(n_609),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_743),
.B(n_667),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_748),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_724),
.A2(n_587),
.B(n_605),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_748),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_782),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_732),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_681),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_787),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_798),
.B(n_667),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_711),
.Y(n_857)
);

NAND2x1p5_ASAP7_75t_L g858 ( 
.A(n_777),
.B(n_577),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_756),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_758),
.B(n_640),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_691),
.B(n_634),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_754),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_740),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_692),
.A2(n_601),
.B(n_580),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_819),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_785),
.B(n_639),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_750),
.B(n_639),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_695),
.B(n_644),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_792),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_806),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_733),
.B(n_791),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_810),
.A2(n_640),
.B1(n_587),
.B2(n_583),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_736),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_819),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_713),
.B(n_569),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_717),
.B(n_544),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_756),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_758),
.B(n_640),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_783),
.B(n_576),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_819),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_783),
.B(n_576),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_R g882 ( 
.A(n_817),
.B(n_544),
.Y(n_882)
);

O2A1O1Ixp5_ASAP7_75t_L g883 ( 
.A1(n_677),
.A2(n_573),
.B(n_616),
.C(n_615),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_741),
.Y(n_884)
);

NAND2x1p5_ASAP7_75t_L g885 ( 
.A(n_777),
.B(n_577),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_808),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_770),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_763),
.A2(n_617),
.B1(n_642),
.B2(n_648),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_SL g889 ( 
.A1(n_805),
.A2(n_529),
.B1(n_654),
.B2(n_665),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_811),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_764),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_812),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_706),
.B(n_644),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_SL g894 ( 
.A(n_818),
.B(n_662),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_686),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_770),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_766),
.A2(n_567),
.B1(n_604),
.B2(n_605),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_797),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_826),
.B(n_662),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_757),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_797),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_689),
.B(n_645),
.Y(n_902)
);

AND2x6_ASAP7_75t_L g903 ( 
.A(n_823),
.B(n_666),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_805),
.B(n_567),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_814),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_676),
.B(n_645),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_682),
.B(n_646),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_750),
.B(n_594),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_703),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_726),
.A2(n_577),
.B(n_589),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_816),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_807),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_690),
.B(n_646),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_697),
.B(n_592),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_828),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_698),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_807),
.Y(n_917)
);

INVx3_ASAP7_75t_SL g918 ( 
.A(n_709),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_710),
.Y(n_919)
);

AND2x6_ASAP7_75t_L g920 ( 
.A(n_823),
.B(n_666),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_824),
.Y(n_921)
);

NAND2x1_ASAP7_75t_L g922 ( 
.A(n_777),
.B(n_589),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_775),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_715),
.B(n_592),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_730),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_824),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_773),
.A2(n_601),
.B1(n_611),
.B2(n_604),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_SL g928 ( 
.A(n_773),
.B(n_565),
.C(n_529),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_766),
.B(n_597),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_772),
.B(n_564),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_777),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_701),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_772),
.B(n_613),
.Y(n_933)
);

BUFx4f_ASAP7_75t_L g934 ( 
.A(n_709),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_708),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_729),
.B(n_610),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_789),
.A2(n_611),
.B1(n_615),
.B2(n_616),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_679),
.A2(n_671),
.B1(n_582),
.B2(n_585),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_789),
.A2(n_571),
.B1(n_559),
.B2(n_561),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_813),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_821),
.Y(n_941)
);

AND2x2_ASAP7_75t_SL g942 ( 
.A(n_699),
.B(n_589),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_771),
.B(n_626),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_701),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_784),
.B(n_671),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_784),
.B(n_607),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_767),
.B(n_607),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_767),
.B(n_607),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_818),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_779),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_688),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_753),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_718),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_732),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_693),
.A2(n_608),
.B(n_559),
.C(n_571),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_699),
.B(n_581),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_701),
.Y(n_957)
);

NOR2x2_ASAP7_75t_L g958 ( 
.A(n_709),
.B(n_608),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_679),
.A2(n_371),
.B1(n_373),
.B2(n_581),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_679),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_719),
.B(n_574),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_723),
.A2(n_572),
.B1(n_574),
.B2(n_563),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_735),
.B(n_572),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_708),
.B(n_524),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_820),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_720),
.Y(n_966)
);

INVx8_ASAP7_75t_L g967 ( 
.A(n_779),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_734),
.B(n_669),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_719),
.B(n_669),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_705),
.B(n_669),
.Y(n_970)
);

AND2x4_ASAP7_75t_SL g971 ( 
.A(n_794),
.B(n_778),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_827),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_774),
.A2(n_563),
.B1(n_543),
.B2(n_530),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_728),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_696),
.B(n_563),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_760),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_723),
.Y(n_977)
);

NAND2x1p5_ASAP7_75t_L g978 ( 
.A(n_827),
.B(n_543),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_801),
.B(n_530),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_765),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_683),
.B(n_543),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_825),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_800),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_719),
.B(n_530),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_802),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_803),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_804),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_801),
.B(n_570),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_778),
.B(n_570),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_719),
.B(n_570),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_794),
.B(n_531),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_719),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_SL g993 ( 
.A(n_680),
.B(n_6),
.C(n_7),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_727),
.A2(n_531),
.B1(n_603),
.B2(n_175),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_675),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_678),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_687),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_684),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_731),
.A2(n_531),
.B1(n_603),
.B2(n_163),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_672),
.A2(n_673),
.B1(n_674),
.B2(n_712),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_753),
.B(n_8),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_809),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_744),
.A2(n_603),
.B1(n_156),
.B2(n_146),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_704),
.B(n_9),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_747),
.B(n_9),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_712),
.A2(n_603),
.B(n_143),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_719),
.B(n_707),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_714),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_862),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_935),
.B(n_793),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_854),
.Y(n_1011)
);

INVx3_ASAP7_75t_SL g1012 ( 
.A(n_853),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_831),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_935),
.B(n_795),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_916),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_932),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_866),
.B(n_753),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_837),
.B(n_774),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_933),
.A2(n_680),
.B1(n_722),
.B2(n_721),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1002),
.B(n_716),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_846),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_849),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_882),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_SL g1024 ( 
.A1(n_908),
.A2(n_751),
.B(n_746),
.C(n_737),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_932),
.B(n_944),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_L g1026 ( 
.A(n_909),
.B(n_744),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_932),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1007),
.A2(n_992),
.B(n_990),
.Y(n_1028)
);

AO32x1_ASAP7_75t_L g1029 ( 
.A1(n_959),
.A2(n_749),
.A3(n_702),
.B1(n_677),
.B2(n_745),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_1007),
.A2(n_768),
.B(n_742),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_867),
.B(n_799),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_857),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_851),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_992),
.A2(n_762),
.B(n_752),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_859),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_865),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_884),
.Y(n_1037)
);

OAI22x1_ASAP7_75t_L g1038 ( 
.A1(n_904),
.A2(n_929),
.B1(n_918),
.B2(n_848),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_871),
.B(n_702),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_871),
.B(n_790),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_888),
.A2(n_796),
.B1(n_822),
.B2(n_745),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_977),
.A2(n_786),
.B(n_749),
.C(n_796),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_876),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_954),
.B(n_739),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_SL g1045 ( 
.A1(n_1005),
.A2(n_788),
.B(n_781),
.C(n_769),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_990),
.A2(n_603),
.B(n_822),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_960),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_888),
.A2(n_603),
.B1(n_13),
.B2(n_15),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_949),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_856),
.A2(n_12),
.B(n_17),
.C(n_24),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_877),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_898),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_901),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_969),
.A2(n_139),
.B(n_138),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_900),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_834),
.A2(n_133),
.B(n_121),
.C(n_113),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_L g1057 ( 
.A(n_830),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_969),
.A2(n_112),
.B(n_106),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_912),
.Y(n_1059)
);

NAND2x2_ASAP7_75t_L g1060 ( 
.A(n_873),
.B(n_12),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_838),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_891),
.B(n_26),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_925),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_917),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1008),
.B(n_101),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_984),
.A2(n_84),
.B(n_79),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_984),
.A2(n_78),
.B(n_76),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_829),
.A2(n_72),
.B(n_70),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_829),
.A2(n_60),
.B(n_30),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_944),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_919),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_921),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_875),
.A2(n_29),
.B(n_33),
.C(n_36),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_977),
.A2(n_37),
.B(n_43),
.C(n_44),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_961),
.A2(n_37),
.B(n_43),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_895),
.B(n_46),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_944),
.B(n_47),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_957),
.Y(n_1078)
);

O2A1O1Ixp5_ASAP7_75t_SL g1079 ( 
.A1(n_959),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_949),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_926),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_906),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_879),
.B(n_51),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_881),
.B(n_51),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_865),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_961),
.A2(n_893),
.B(n_910),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_942),
.A2(n_53),
.B1(n_55),
.B2(n_952),
.Y(n_1087)
);

AOI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_1004),
.A2(n_55),
.B(n_893),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_965),
.B(n_964),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_897),
.B(n_836),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_906),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_942),
.A2(n_952),
.B1(n_844),
.B2(n_945),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_907),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_997),
.B(n_889),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_983),
.B(n_985),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_SL g1096 ( 
.A(n_928),
.B(n_847),
.C(n_841),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_860),
.B(n_878),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_860),
.B(n_878),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_907),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_945),
.A2(n_1001),
.B1(n_971),
.B2(n_836),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_986),
.B(n_987),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_957),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_940),
.B(n_941),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1001),
.A2(n_958),
.B1(n_993),
.B2(n_872),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_955),
.A2(n_973),
.A3(n_979),
.B(n_988),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_913),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_850),
.A2(n_991),
.B(n_864),
.C(n_934),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_957),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_910),
.A2(n_948),
.B(n_947),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_SL g1110 ( 
.A(n_843),
.B(n_894),
.C(n_936),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_913),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_947),
.A2(n_948),
.B(n_902),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_914),
.Y(n_1113)
);

INVx6_ASAP7_75t_L g1114 ( 
.A(n_830),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_934),
.B(n_943),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_902),
.A2(n_868),
.B(n_861),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_861),
.A2(n_868),
.B(n_963),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_899),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_943),
.B(n_928),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_914),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_830),
.B(n_832),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_924),
.B(n_903),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_956),
.A2(n_946),
.B1(n_938),
.B2(n_1000),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_883),
.A2(n_956),
.B(n_946),
.Y(n_1124)
);

AOI221xp5_ASAP7_75t_L g1125 ( 
.A1(n_993),
.A2(n_899),
.B1(n_833),
.B2(n_835),
.C(n_892),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_832),
.B(n_863),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_845),
.A2(n_885),
.B(n_858),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_924),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_903),
.B(n_920),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_953),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_938),
.A2(n_927),
.B1(n_1003),
.B2(n_840),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_845),
.A2(n_885),
.B(n_858),
.Y(n_1132)
);

XOR2x2_ASAP7_75t_L g1133 ( 
.A(n_968),
.B(n_975),
.Y(n_1133)
);

INVx5_ASAP7_75t_L g1134 ( 
.A(n_931),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_905),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_931),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_865),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_911),
.Y(n_1138)
);

INVx8_ASAP7_75t_L g1139 ( 
.A(n_967),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_915),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_L g1141 ( 
.A(n_903),
.B(n_920),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_842),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_966),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_976),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_852),
.B(n_890),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_920),
.B(n_855),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_869),
.B(n_886),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_870),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_L g1149 ( 
.A(n_832),
.B(n_863),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_SL g1150 ( 
.A(n_970),
.B(n_999),
.C(n_994),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_972),
.A2(n_922),
.B(n_981),
.Y(n_1151)
);

INVx3_ASAP7_75t_SL g1152 ( 
.A(n_863),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_972),
.A2(n_989),
.B(n_839),
.Y(n_1153)
);

NAND2x1p5_ASAP7_75t_L g1154 ( 
.A(n_931),
.B(n_880),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_980),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_972),
.A2(n_874),
.B(n_967),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_880),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1127),
.A2(n_883),
.B(n_973),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1055),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1139),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_L g1161 ( 
.A(n_1095),
.B(n_967),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1145),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_SL g1163 ( 
.A(n_1023),
.B(n_880),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1123),
.A2(n_1006),
.B(n_939),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_1011),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1034),
.A2(n_978),
.B(n_937),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1015),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1088),
.A2(n_982),
.B1(n_951),
.B2(n_974),
.C(n_962),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1028),
.A2(n_978),
.B(n_998),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1089),
.B(n_998),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1123),
.A2(n_995),
.B(n_996),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1030),
.A2(n_972),
.B(n_896),
.Y(n_1172)
);

OR2x6_ASAP7_75t_L g1173 ( 
.A(n_1139),
.B(n_1115),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1128),
.B(n_887),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1116),
.A2(n_995),
.B(n_996),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1031),
.A2(n_887),
.B(n_896),
.C(n_923),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1112),
.A2(n_923),
.B(n_950),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1071),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1107),
.A2(n_950),
.B(n_1131),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1124),
.A2(n_1117),
.B(n_1042),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1151),
.A2(n_1153),
.B(n_1124),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1082),
.B(n_1091),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1045),
.A2(n_1024),
.B(n_1141),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1017),
.B(n_1098),
.Y(n_1184)
);

AOI211x1_ASAP7_75t_L g1185 ( 
.A1(n_1087),
.A2(n_1048),
.B(n_1095),
.C(n_1101),
.Y(n_1185)
);

NOR2xp67_ASAP7_75t_L g1186 ( 
.A(n_1043),
.B(n_1009),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1150),
.A2(n_1122),
.B(n_1100),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1037),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1129),
.A2(n_1146),
.B(n_1046),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_1012),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1094),
.B(n_1101),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1103),
.A2(n_1090),
.B1(n_1092),
.B2(n_1087),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1040),
.A2(n_1088),
.B(n_1103),
.C(n_1019),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1100),
.A2(n_1092),
.A3(n_1131),
.B(n_1041),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1093),
.B(n_1099),
.Y(n_1195)
);

AOI221x1_ASAP7_75t_L g1196 ( 
.A1(n_1038),
.A2(n_1048),
.B1(n_1104),
.B2(n_1096),
.C(n_1019),
.Y(n_1196)
);

NAND3x1_ASAP7_75t_L g1197 ( 
.A(n_1119),
.B(n_1084),
.C(n_1083),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1156),
.A2(n_1065),
.B(n_1041),
.Y(n_1198)
);

AOI221xp5_ASAP7_75t_L g1199 ( 
.A1(n_1104),
.A2(n_1073),
.B1(n_1050),
.B2(n_1061),
.C(n_1074),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1065),
.A2(n_1058),
.B(n_1054),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1020),
.A2(n_1010),
.B(n_1014),
.C(n_1026),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1133),
.A2(n_1106),
.B(n_1111),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1062),
.A2(n_1037),
.B(n_1069),
.C(n_1075),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1018),
.B(n_1039),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1079),
.A2(n_1068),
.B(n_1067),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1066),
.A2(n_1154),
.B(n_1081),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1154),
.A2(n_1013),
.B(n_1053),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1021),
.A2(n_1035),
.B(n_1022),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1139),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1063),
.A2(n_1097),
.B1(n_1147),
.B2(n_1125),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1029),
.A2(n_1149),
.B(n_1134),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1033),
.A2(n_1064),
.B(n_1052),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1029),
.A2(n_1105),
.A3(n_1135),
.B(n_1148),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1138),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1051),
.A2(n_1072),
.B(n_1059),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1121),
.A2(n_1126),
.B(n_1025),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1016),
.B(n_1108),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1140),
.B(n_1142),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1057),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1076),
.A2(n_1056),
.B(n_1110),
.Y(n_1220)
);

AOI221xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1130),
.A2(n_1155),
.B1(n_1143),
.B2(n_1144),
.C(n_1157),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1118),
.B(n_1032),
.C(n_1047),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1036),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1152),
.B(n_1085),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1137),
.A2(n_1077),
.B(n_1105),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1044),
.B(n_1105),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1057),
.A2(n_1136),
.B(n_1134),
.C(n_1027),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1157),
.B(n_1027),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_SL g1229 ( 
.A(n_1080),
.B(n_1027),
.Y(n_1229)
);

CKINVDCx14_ASAP7_75t_R g1230 ( 
.A(n_1049),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1114),
.B(n_1070),
.Y(n_1231)
);

INVxp67_ASAP7_75t_SL g1232 ( 
.A(n_1078),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1102),
.B(n_1060),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1102),
.A2(n_1132),
.B(n_1127),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1037),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1031),
.A2(n_933),
.B(n_908),
.C(n_815),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1145),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1043),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1116),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1127),
.A2(n_1132),
.B(n_1086),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1145),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1017),
.B(n_866),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1031),
.A2(n_933),
.B(n_908),
.C(n_815),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1017),
.B(n_866),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1145),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1127),
.A2(n_1132),
.B(n_1086),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1009),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1043),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1127),
.A2(n_1132),
.B(n_1086),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1145),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1123),
.A2(n_1100),
.A3(n_1109),
.B(n_1092),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1089),
.A2(n_933),
.B1(n_908),
.B2(n_867),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1116),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1031),
.A2(n_933),
.B(n_908),
.C(n_815),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1089),
.B(n_658),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1145),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1123),
.A2(n_933),
.B(n_1086),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1127),
.A2(n_1132),
.B(n_1086),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1123),
.A2(n_1100),
.A3(n_1109),
.B(n_1092),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1123),
.A2(n_1100),
.A3(n_1109),
.B(n_1092),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1127),
.A2(n_1132),
.B(n_1086),
.Y(n_1269)
);

AOI21xp33_ASAP7_75t_L g1270 ( 
.A1(n_1019),
.A2(n_933),
.B(n_908),
.Y(n_1270)
);

AOI21xp33_ASAP7_75t_L g1271 ( 
.A1(n_1019),
.A2(n_933),
.B(n_908),
.Y(n_1271)
);

OAI21xp33_ASAP7_75t_L g1272 ( 
.A1(n_1095),
.A2(n_933),
.B(n_908),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1157),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1116),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1116),
.Y(n_1276)
);

AOI221x1_ASAP7_75t_L g1277 ( 
.A1(n_1087),
.A2(n_1100),
.B1(n_1038),
.B2(n_1048),
.C(n_1104),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1089),
.B(n_933),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_SL g1279 ( 
.A1(n_1107),
.A2(n_933),
.B(n_1065),
.C(n_834),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1145),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1017),
.B(n_866),
.Y(n_1281)
);

O2A1O1Ixp5_ASAP7_75t_SL g1282 ( 
.A1(n_1100),
.A2(n_838),
.B(n_834),
.C(n_1088),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1017),
.B(n_866),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_SL g1284 ( 
.A1(n_1119),
.A2(n_1122),
.B(n_1129),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1145),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1017),
.B(n_866),
.Y(n_1286)
);

INVx6_ASAP7_75t_SL g1287 ( 
.A(n_1097),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1123),
.A2(n_933),
.B(n_1086),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1097),
.B(n_1098),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_SL g1290 ( 
.A(n_1087),
.B(n_933),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1090),
.B(n_528),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1095),
.A2(n_933),
.B1(n_1103),
.B2(n_1101),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1145),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1278),
.B(n_1191),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1237),
.A2(n_1261),
.B(n_1246),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1208),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1239),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1236),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1218),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1259),
.B(n_1290),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1212),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1183),
.A2(n_1196),
.A3(n_1277),
.B(n_1211),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1255),
.A2(n_1269),
.B(n_1266),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1291),
.B(n_1162),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1159),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1270),
.B(n_1271),
.C(n_1272),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1188),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1184),
.B(n_1245),
.Y(n_1308)
);

OAI21xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1235),
.A2(n_1242),
.B(n_1241),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1205),
.A2(n_1288),
.B(n_1265),
.Y(n_1310)
);

INVx6_ASAP7_75t_SL g1311 ( 
.A(n_1173),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1292),
.A2(n_1210),
.B1(n_1202),
.B2(n_1242),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1247),
.B(n_1281),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1292),
.B(n_1235),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1244),
.B(n_1256),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1241),
.B(n_1250),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1218),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1167),
.Y(n_1318)
);

BUFx2_ASAP7_75t_SL g1319 ( 
.A(n_1219),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1163),
.B(n_1273),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1192),
.A2(n_1199),
.B1(n_1286),
.B2(n_1283),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1165),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1230),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1181),
.A2(n_1177),
.B(n_1172),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1205),
.A2(n_1180),
.B(n_1164),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1178),
.Y(n_1326)
);

NAND2x1p5_ASAP7_75t_L g1327 ( 
.A(n_1273),
.B(n_1160),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1158),
.A2(n_1189),
.B(n_1169),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1193),
.A2(n_1201),
.B(n_1282),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1192),
.A2(n_1164),
.B1(n_1204),
.B2(n_1262),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1219),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1180),
.A2(n_1198),
.B(n_1200),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1166),
.A2(n_1206),
.B(n_1175),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1203),
.A2(n_1279),
.B(n_1170),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1219),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1221),
.A2(n_1171),
.B(n_1175),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1238),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1284),
.A2(n_1225),
.B(n_1171),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1250),
.B(n_1252),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_1229),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1179),
.A2(n_1207),
.B(n_1220),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_SL g1342 ( 
.A1(n_1220),
.A2(n_1176),
.B(n_1204),
.C(n_1254),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1214),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1289),
.B(n_1293),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1252),
.B(n_1263),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1254),
.B(n_1258),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1221),
.A2(n_1168),
.B(n_1182),
.Y(n_1347)
);

INVx3_ASAP7_75t_R g1348 ( 
.A(n_1224),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1215),
.A2(n_1174),
.B(n_1216),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1187),
.A2(n_1161),
.B(n_1258),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1274),
.A2(n_1197),
.B1(n_1182),
.B2(n_1195),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1274),
.B(n_1251),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1185),
.B(n_1173),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1248),
.B(n_1280),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1213),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1160),
.B(n_1209),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1264),
.B(n_1285),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_SL g1358 ( 
.A1(n_1227),
.A2(n_1233),
.B(n_1223),
.C(n_1228),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1194),
.A2(n_1222),
.B(n_1229),
.C(n_1268),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1232),
.B(n_1194),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1186),
.B(n_1194),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1231),
.B(n_1217),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1257),
.B(n_1267),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1257),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1267),
.B(n_1268),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1267),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1287),
.A2(n_1217),
.B1(n_1190),
.B2(n_1273),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1287),
.A2(n_1259),
.B1(n_1237),
.B2(n_1246),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1268),
.B(n_1253),
.Y(n_1369)
);

AOI31xp67_ASAP7_75t_L g1370 ( 
.A1(n_1226),
.A2(n_834),
.A3(n_838),
.B(n_856),
.Y(n_1370)
);

AO21x2_ASAP7_75t_L g1371 ( 
.A1(n_1183),
.A2(n_1260),
.B(n_1240),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1218),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1179),
.B(n_1185),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1218),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1219),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1270),
.A2(n_1271),
.B1(n_1290),
.B2(n_1278),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1290),
.A2(n_1259),
.B1(n_1278),
.B2(n_810),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1237),
.A2(n_1246),
.B(n_1261),
.C(n_933),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1179),
.B(n_1185),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1218),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1184),
.B(n_1245),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1219),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1240),
.A2(n_1260),
.A3(n_1276),
.B(n_1275),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1278),
.A2(n_933),
.B1(n_1259),
.B2(n_1290),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1218),
.Y(n_1385)
);

INVx3_ASAP7_75t_SL g1386 ( 
.A(n_1239),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1208),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1219),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1291),
.B(n_1162),
.Y(n_1389)
);

NAND3xp33_ASAP7_75t_L g1390 ( 
.A(n_1237),
.B(n_1261),
.C(n_1246),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1208),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1239),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1184),
.B(n_1245),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1184),
.B(n_1245),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1184),
.B(n_1245),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1159),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1163),
.B(n_1273),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1219),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1278),
.B(n_1191),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1184),
.B(n_1245),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1218),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1219),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1234),
.A2(n_1249),
.B(n_1243),
.Y(n_1403)
);

NAND4xp25_ASAP7_75t_L g1404 ( 
.A(n_1191),
.B(n_1278),
.C(n_763),
.D(n_810),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1183),
.A2(n_1260),
.B(n_1240),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1240),
.A2(n_1260),
.A3(n_1276),
.B(n_1275),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1218),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1208),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1230),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1404),
.A2(n_1377),
.B(n_1378),
.C(n_1399),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1384),
.A2(n_1378),
.B(n_1377),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1294),
.A2(n_1300),
.B(n_1312),
.C(n_1295),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1313),
.B(n_1308),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1300),
.A2(n_1368),
.B(n_1376),
.C(n_1334),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1304),
.B(n_1389),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1346),
.B(n_1314),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1376),
.A2(n_1351),
.B(n_1359),
.C(n_1390),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1359),
.A2(n_1329),
.B(n_1306),
.C(n_1358),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1346),
.A2(n_1340),
.B1(n_1339),
.B2(n_1316),
.Y(n_1419)
);

CKINVDCx6p67_ASAP7_75t_R g1420 ( 
.A(n_1386),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1381),
.B(n_1393),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1345),
.B(n_1309),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1423)
);

BUFx8_ASAP7_75t_SL g1424 ( 
.A(n_1323),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1315),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1311),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1321),
.A2(n_1352),
.B1(n_1330),
.B2(n_1337),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1321),
.A2(n_1352),
.B1(n_1330),
.B2(n_1379),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1361),
.B(n_1400),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1373),
.A2(n_1379),
.B1(n_1407),
.B2(n_1317),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1299),
.B(n_1372),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1374),
.B(n_1380),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1373),
.A2(n_1379),
.B1(n_1401),
.B2(n_1385),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1358),
.A2(n_1342),
.B(n_1298),
.C(n_1373),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1297),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_SL g1436 ( 
.A1(n_1369),
.A2(n_1363),
.B(n_1356),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1302),
.B(n_1360),
.Y(n_1437)
);

AOI21x1_ASAP7_75t_SL g1438 ( 
.A1(n_1369),
.A2(n_1356),
.B(n_1354),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1344),
.B(n_1362),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1353),
.A2(n_1326),
.B1(n_1318),
.B2(n_1343),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1357),
.B(n_1307),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1342),
.A2(n_1353),
.B(n_1367),
.C(n_1325),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1311),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1302),
.B(n_1347),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1392),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1353),
.A2(n_1322),
.B(n_1388),
.C(n_1398),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1375),
.A2(n_1388),
.B(n_1398),
.C(n_1305),
.Y(n_1447)
);

AOI211xp5_ASAP7_75t_L g1448 ( 
.A1(n_1386),
.A2(n_1341),
.B(n_1396),
.C(n_1331),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1302),
.B(n_1347),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1302),
.B(n_1347),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1392),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1310),
.B(n_1350),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1311),
.A2(n_1365),
.B1(n_1397),
.B2(n_1320),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1320),
.A2(n_1397),
.B(n_1327),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1335),
.A2(n_1364),
.B(n_1366),
.C(n_1350),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1396),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1327),
.A2(n_1336),
.B(n_1382),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1338),
.A2(n_1333),
.B(n_1328),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1349),
.Y(n_1459)
);

O2A1O1Ixp5_ASAP7_75t_L g1460 ( 
.A1(n_1296),
.A2(n_1301),
.B(n_1408),
.C(n_1387),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1336),
.A2(n_1402),
.B(n_1405),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1348),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1319),
.Y(n_1463)
);

AND2x4_ASAP7_75t_SL g1464 ( 
.A(n_1409),
.B(n_1323),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1371),
.B(n_1355),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1338),
.A2(n_1333),
.B(n_1328),
.Y(n_1466)
);

AND2x4_ASAP7_75t_SL g1467 ( 
.A(n_1409),
.B(n_1296),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1341),
.B(n_1332),
.Y(n_1468)
);

AOI21x1_ASAP7_75t_SL g1469 ( 
.A1(n_1370),
.A2(n_1332),
.B(n_1383),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1391),
.Y(n_1470)
);

AOI21x1_ASAP7_75t_SL g1471 ( 
.A1(n_1383),
.A2(n_1406),
.B(n_1324),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1383),
.B(n_1406),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1406),
.B(n_1303),
.Y(n_1473)
);

O2A1O1Ixp5_ASAP7_75t_L g1474 ( 
.A1(n_1403),
.A2(n_1271),
.B(n_1270),
.C(n_1237),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1384),
.A2(n_1246),
.B(n_1237),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1346),
.B(n_1314),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1313),
.B(n_1308),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1404),
.A2(n_1246),
.B(n_1261),
.C(n_1237),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_SL g1479 ( 
.A1(n_1300),
.A2(n_933),
.B(n_867),
.C(n_930),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1384),
.A2(n_1246),
.B(n_1237),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1329),
.A2(n_1205),
.B(n_1183),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1313),
.B(n_1308),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1313),
.B(n_1308),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1384),
.A2(n_1246),
.B(n_1237),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1396),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1428),
.A2(n_1427),
.B1(n_1419),
.B2(n_1462),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1416),
.B(n_1476),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1429),
.B(n_1437),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1458),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1470),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1479),
.A2(n_1411),
.B(n_1475),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1415),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1416),
.B(n_1476),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1427),
.A2(n_1428),
.B1(n_1410),
.B2(n_1412),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1468),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1437),
.B(n_1481),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1460),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1422),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1422),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1465),
.B(n_1452),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1419),
.A2(n_1425),
.B1(n_1441),
.B2(n_1413),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1459),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1444),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1444),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1449),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1506)
);

BUFx4f_ASAP7_75t_SL g1507 ( 
.A(n_1420),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1457),
.B(n_1461),
.Y(n_1508)
);

BUFx4f_ASAP7_75t_SL g1509 ( 
.A(n_1485),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1450),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1464),
.Y(n_1511)
);

OR2x6_ASAP7_75t_L g1512 ( 
.A(n_1442),
.B(n_1446),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1440),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1467),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1431),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1466),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1474),
.A2(n_1472),
.B(n_1473),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1440),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1431),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1481),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1466),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1430),
.B(n_1433),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1432),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1432),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1430),
.A2(n_1433),
.A3(n_1453),
.B(n_1469),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1453),
.B(n_1484),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1455),
.Y(n_1527)
);

AO21x1_ASAP7_75t_SL g1528 ( 
.A1(n_1448),
.A2(n_1438),
.B(n_1417),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1418),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1423),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1421),
.B(n_1483),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1508),
.B(n_1434),
.Y(n_1532)
);

INVx4_ASAP7_75t_SL g1533 ( 
.A(n_1525),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1500),
.B(n_1482),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1502),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1496),
.B(n_1477),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1494),
.A2(n_1414),
.B1(n_1439),
.B2(n_1478),
.Y(n_1537)
);

AND2x2_ASAP7_75t_SL g1538 ( 
.A(n_1518),
.B(n_1436),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1498),
.B(n_1456),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1497),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1516),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1499),
.B(n_1456),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1495),
.B(n_1471),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1489),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1506),
.B(n_1426),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1495),
.B(n_1520),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1489),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1488),
.B(n_1447),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1515),
.B(n_1519),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1527),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1520),
.B(n_1443),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1529),
.B(n_1454),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1503),
.Y(n_1555)
);

BUFx2_ASAP7_75t_SL g1556 ( 
.A(n_1514),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1545),
.A2(n_1521),
.B(n_1497),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1537),
.A2(n_1491),
.B1(n_1486),
.B2(n_1529),
.C(n_1526),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1535),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1548),
.B(n_1517),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1539),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1539),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1535),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1548),
.B(n_1517),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1536),
.B(n_1517),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1556),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1537),
.A2(n_1501),
.B1(n_1518),
.B2(n_1526),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1541),
.Y(n_1569)
);

AOI33xp33_ASAP7_75t_L g1570 ( 
.A1(n_1553),
.A2(n_1501),
.A3(n_1492),
.B1(n_1527),
.B2(n_1524),
.B3(n_1523),
.Y(n_1570)
);

OAI211xp5_ASAP7_75t_L g1571 ( 
.A1(n_1532),
.A2(n_1513),
.B(n_1487),
.C(n_1493),
.Y(n_1571)
);

OAI33xp33_ASAP7_75t_L g1572 ( 
.A1(n_1552),
.A2(n_1510),
.A3(n_1505),
.B1(n_1504),
.B2(n_1523),
.B3(n_1524),
.Y(n_1572)
);

OAI221xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1552),
.A2(n_1512),
.B1(n_1530),
.B2(n_1522),
.C(n_1511),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1538),
.A2(n_1512),
.B(n_1530),
.Y(n_1574)
);

AO21x1_ASAP7_75t_SL g1575 ( 
.A1(n_1550),
.A2(n_1522),
.B(n_1510),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1538),
.B(n_1554),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_SL g1577 ( 
.A(n_1550),
.B(n_1528),
.C(n_1463),
.D(n_1531),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_SL g1578 ( 
.A(n_1534),
.B(n_1490),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1536),
.B(n_1517),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1546),
.B(n_1506),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1555),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1505),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1542),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1581),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1583),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1558),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1558),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1581),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1583),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1583),
.B(n_1533),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1574),
.A2(n_1549),
.B(n_1544),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1562),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1578),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1562),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1583),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1563),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1560),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1560),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_SL g1599 ( 
.A(n_1577),
.B(n_1435),
.C(n_1445),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1583),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1564),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1569),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1578),
.Y(n_1603)
);

INVx4_ASAP7_75t_SL g1604 ( 
.A(n_1583),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1582),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1586),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1593),
.B(n_1566),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1592),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1593),
.B(n_1603),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1593),
.A2(n_1576),
.B(n_1574),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1603),
.B(n_1591),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1591),
.B(n_1566),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1591),
.B(n_1579),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1592),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1591),
.A2(n_1576),
.B1(n_1577),
.B2(n_1559),
.Y(n_1616)
);

NAND3xp33_ASAP7_75t_L g1617 ( 
.A(n_1599),
.B(n_1571),
.C(n_1559),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1605),
.B(n_1570),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1602),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1591),
.B(n_1579),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1604),
.B(n_1579),
.Y(n_1622)
);

OAI33xp33_ASAP7_75t_L g1623 ( 
.A1(n_1584),
.A2(n_1568),
.A3(n_1580),
.B1(n_1551),
.B2(n_1547),
.B3(n_1543),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1604),
.B(n_1561),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1586),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

OAI321xp33_ASAP7_75t_L g1628 ( 
.A1(n_1589),
.A2(n_1571),
.A3(n_1568),
.B1(n_1573),
.B2(n_1512),
.C(n_1540),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1596),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1604),
.B(n_1561),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1604),
.B(n_1561),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1605),
.B(n_1570),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1604),
.B(n_1565),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1604),
.B(n_1565),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1588),
.B(n_1569),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1595),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1587),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1597),
.B(n_1580),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1617),
.A2(n_1599),
.B(n_1573),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1624),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1618),
.B(n_1534),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1610),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1630),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1618),
.B(n_1534),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1630),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1633),
.B(n_1610),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1624),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1609),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1633),
.B(n_1531),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1609),
.B(n_1590),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1609),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1625),
.B(n_1575),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1640),
.B(n_1598),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1617),
.A2(n_1528),
.B1(n_1538),
.B2(n_1512),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1619),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1619),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1616),
.A2(n_1538),
.B1(n_1512),
.B2(n_1567),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1628),
.A2(n_1572),
.B(n_1451),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1608),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1625),
.B(n_1575),
.Y(n_1663)
);

NOR2xp67_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1595),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1638),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1606),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1606),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1640),
.B(n_1557),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1625),
.B(n_1590),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1606),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1631),
.B(n_1590),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1623),
.B(n_1424),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1638),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1608),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1642),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1649),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1652),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1672),
.B(n_1507),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1649),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_L g1681 ( 
.A1(n_1648),
.A2(n_1612),
.B(n_1611),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1644),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1657),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1666),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1641),
.B(n_1612),
.C(n_1638),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1652),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1664),
.A2(n_1612),
.B(n_1637),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1650),
.B(n_1607),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1653),
.B(n_1607),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1669),
.B(n_1631),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1657),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1669),
.B(n_1631),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1652),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1665),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1658),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1661),
.B(n_1607),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1666),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1667),
.Y(n_1698)
);

INVxp33_ASAP7_75t_L g1699 ( 
.A(n_1651),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1671),
.B(n_1632),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1679),
.B(n_1682),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1690),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1675),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1696),
.B(n_1643),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1688),
.B(n_1646),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1675),
.B(n_1656),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1690),
.B(n_1671),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1699),
.B(n_1685),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1692),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1685),
.A2(n_1623),
.B1(n_1660),
.B2(n_1647),
.C(n_1645),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1678),
.Y(n_1713)
);

OAI322xp33_ASAP7_75t_L g1714 ( 
.A1(n_1676),
.A2(n_1647),
.A3(n_1655),
.B1(n_1659),
.B2(n_1662),
.C1(n_1674),
.C2(n_1665),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1687),
.B(n_1673),
.C(n_1662),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

AOI311xp33_ASAP7_75t_L g1717 ( 
.A1(n_1677),
.A2(n_1674),
.A3(n_1668),
.B(n_1629),
.C(n_1615),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1681),
.A2(n_1654),
.B1(n_1663),
.B2(n_1673),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1692),
.B(n_1654),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1704),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1704),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1713),
.B(n_1686),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1712),
.B(n_1681),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1709),
.B(n_1715),
.Y(n_1725)
);

CKINVDCx16_ASAP7_75t_R g1726 ( 
.A(n_1701),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1713),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1711),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1708),
.B(n_1719),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1711),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1720),
.B(n_1686),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1714),
.B(n_1694),
.Y(n_1732)
);

AND5x1_ASAP7_75t_L g1733 ( 
.A(n_1724),
.B(n_1718),
.C(n_1705),
.D(n_1717),
.E(n_1720),
.Y(n_1733)
);

AOI22x1_ASAP7_75t_L g1734 ( 
.A1(n_1726),
.A2(n_1694),
.B1(n_1710),
.B2(n_1702),
.Y(n_1734)
);

NOR3xp33_ASAP7_75t_L g1735 ( 
.A(n_1725),
.B(n_1707),
.C(n_1703),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1725),
.B(n_1721),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1729),
.B(n_1677),
.Y(n_1737)
);

OAI21xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1724),
.A2(n_1700),
.B(n_1689),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1732),
.A2(n_1706),
.B(n_1716),
.C(n_1680),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1727),
.B(n_1680),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1723),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1722),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1728),
.A2(n_1700),
.B1(n_1691),
.B2(n_1695),
.Y(n_1743)
);

AOI221x1_ASAP7_75t_L g1744 ( 
.A1(n_1739),
.A2(n_1730),
.B1(n_1731),
.B2(n_1683),
.C(n_1691),
.Y(n_1744)
);

NOR4xp25_ASAP7_75t_L g1745 ( 
.A(n_1742),
.B(n_1695),
.C(n_1697),
.D(n_1698),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1736),
.A2(n_1655),
.B1(n_1611),
.B2(n_1585),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1736),
.A2(n_1698),
.B(n_1697),
.C(n_1684),
.Y(n_1747)
);

AOI322xp5_ASAP7_75t_L g1748 ( 
.A1(n_1735),
.A2(n_1614),
.A3(n_1620),
.B1(n_1613),
.B2(n_1611),
.C1(n_1622),
.C2(n_1632),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1737),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1738),
.A2(n_1733),
.B(n_1741),
.C(n_1740),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1747),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1749),
.B(n_1743),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1750),
.B(n_1734),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1744),
.B(n_1698),
.Y(n_1754)
);

NOR3xp33_ASAP7_75t_L g1755 ( 
.A(n_1746),
.B(n_1697),
.C(n_1684),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1745),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1748),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1753),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1752),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1754),
.B(n_1638),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_R g1761 ( 
.A(n_1751),
.B(n_1509),
.Y(n_1761)
);

AOI322xp5_ASAP7_75t_L g1762 ( 
.A1(n_1757),
.A2(n_1614),
.A3(n_1620),
.B1(n_1613),
.B2(n_1684),
.C1(n_1622),
.C2(n_1632),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1760),
.Y(n_1763)
);

AND4x1_ASAP7_75t_L g1764 ( 
.A(n_1761),
.B(n_1756),
.C(n_1755),
.D(n_1759),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1758),
.A2(n_1638),
.B1(n_1636),
.B2(n_1659),
.Y(n_1765)
);

NAND3x1_ASAP7_75t_L g1766 ( 
.A(n_1764),
.B(n_1762),
.C(n_1635),
.Y(n_1766)
);

AOI22x1_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1763),
.B1(n_1765),
.B2(n_1667),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1767),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1767),
.A2(n_1670),
.B1(n_1595),
.B2(n_1600),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1768),
.Y(n_1770)
);

AO22x1_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_1670),
.B1(n_1634),
.B2(n_1635),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1770),
.A2(n_1585),
.B1(n_1490),
.B2(n_1636),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1772),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1773),
.B(n_1771),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1774),
.B(n_1636),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1627),
.B1(n_1621),
.B2(n_1626),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1634),
.B1(n_1635),
.B2(n_1626),
.Y(n_1777)
);

AOI211xp5_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1627),
.B(n_1626),
.C(n_1639),
.Y(n_1778)
);


endmodule