module fake_jpeg_18836_n_123 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_66),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_0),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_49),
.C(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_77),
.Y(n_82)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_0),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_51),
.B1(n_46),
.B2(n_52),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_6),
.B(n_8),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_48),
.B1(n_58),
.B2(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_60),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_19),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_54),
.B1(n_47),
.B2(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_12),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_16),
.B1(n_41),
.B2(n_33),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_1),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_2),
.B(n_3),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_9),
.B(n_11),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_21),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_99),
.B1(n_98),
.B2(n_27),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_111),
.Y(n_114)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_98),
.C(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_115),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_118),
.B(n_110),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_114),
.B(n_109),
.C(n_112),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_23),
.C(n_24),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_121),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_28),
.C(n_32),
.Y(n_123)
);


endmodule