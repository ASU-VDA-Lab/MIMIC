module fake_jpeg_837_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_74),
.B1(n_52),
.B2(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_60),
.Y(n_73)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_56),
.B1(n_48),
.B2(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_60),
.B1(n_59),
.B2(n_41),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_87),
.B1(n_65),
.B2(n_52),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_64),
.B1(n_51),
.B2(n_6),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_73),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_59),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_89),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_44),
.B1(n_41),
.B2(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_50),
.Y(n_89)
);

BUFx2_ASAP7_75t_SL g91 ( 
.A(n_88),
.Y(n_91)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_99),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_104),
.B1(n_9),
.B2(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_24),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_101),
.Y(n_113)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_8),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_51),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_22),
.C(n_39),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_119),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_76),
.B1(n_75),
.B2(n_51),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_27),
.B1(n_14),
.B2(n_15),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_121),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_7),
.B(n_8),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_110),
.B(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_7),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_11),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_25),
.C(n_38),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_28),
.C(n_18),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_138),
.B1(n_111),
.B2(n_116),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_135),
.B(n_137),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_31),
.B(n_19),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_13),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_136),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_124),
.B1(n_21),
.B2(n_23),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_148),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_129),
.C(n_133),
.Y(n_148)
);

OAI22x1_ASAP7_75t_SL g151 ( 
.A1(n_149),
.A2(n_140),
.B1(n_141),
.B2(n_128),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_147),
.C(n_148),
.Y(n_152)
);

NAND4xp25_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_150),
.C(n_139),
.D(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_145),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_125),
.C(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_134),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_20),
.B(n_32),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_40),
.Y(n_159)
);


endmodule