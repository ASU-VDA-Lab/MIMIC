module fake_jpeg_20865_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_53),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_0),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_37),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_48),
.B1(n_41),
.B2(n_46),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_60),
.B1(n_38),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_3),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_45),
.B1(n_19),
.B2(n_22),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_63),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_5),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_40),
.B(n_2),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_77),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_4),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_88),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_74),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_87),
.B1(n_75),
.B2(n_85),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_70),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_86),
.A3(n_87),
.B1(n_14),
.B2(n_16),
.C1(n_17),
.C2(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_10),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_99),
.B1(n_92),
.B2(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_96),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_26),
.CI(n_27),
.CON(n_105),
.SN(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_28),
.B(n_30),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_105),
.Y(n_107)
);


endmodule