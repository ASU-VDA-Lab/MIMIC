module real_aes_10730_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_1801, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_1801;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_1382;
wire n_1199;
wire n_951;
wire n_875;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_1767;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_1779;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_1772;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_1369;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_0), .A2(n_152), .B1(n_459), .B2(n_700), .C(n_701), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_0), .A2(n_308), .B1(n_757), .B2(n_758), .C(n_760), .Y(n_756) );
INVx1_ASAP7_75t_L g787 ( .A(n_1), .Y(n_787) );
INVx1_ASAP7_75t_L g921 ( .A(n_2), .Y(n_921) );
INVx1_ASAP7_75t_L g1505 ( .A(n_3), .Y(n_1505) );
INVxp33_ASAP7_75t_L g1245 ( .A(n_4), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1325 ( .A1(n_4), .A2(n_86), .B1(n_1143), .B2(n_1317), .Y(n_1325) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_5), .A2(n_136), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_5), .A2(n_47), .B1(n_998), .B2(n_1170), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1767 ( .A1(n_6), .A2(n_233), .B1(n_1199), .B2(n_1352), .C(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1796 ( .A(n_6), .Y(n_1796) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_7), .A2(n_54), .B1(n_601), .B2(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g676 ( .A(n_7), .Y(n_676) );
XNOR2x2_ASAP7_75t_L g1134 ( .A(n_8), .B(n_1135), .Y(n_1134) );
AOI22xp33_ASAP7_75t_SL g1145 ( .A1(n_9), .A2(n_47), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
AOI21xp33_ASAP7_75t_L g1171 ( .A1(n_9), .A2(n_580), .B(n_822), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g1382 ( .A(n_10), .Y(n_1382) );
AOI22xp5_ASAP7_75t_L g1475 ( .A1(n_11), .A2(n_105), .B1(n_1476), .B2(n_1484), .Y(n_1475) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_12), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_12), .A2(n_50), .B1(n_391), .B2(n_418), .C(n_916), .Y(n_1063) );
INVxp33_ASAP7_75t_L g1251 ( .A(n_13), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_13), .A2(n_179), .B1(n_675), .B2(n_1319), .Y(n_1324) );
INVxp33_ASAP7_75t_L g797 ( .A(n_14), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_14), .A2(n_64), .B1(n_860), .B2(n_862), .C(n_863), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_15), .A2(n_60), .B1(n_1339), .B2(n_1340), .C(n_1341), .Y(n_1338) );
INVx1_ASAP7_75t_L g1366 ( .A(n_15), .Y(n_1366) );
INVx1_ASAP7_75t_L g1161 ( .A(n_16), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_16), .A2(n_264), .B1(n_822), .B2(n_998), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_17), .A2(n_303), .B1(n_570), .B2(n_618), .C(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g659 ( .A(n_17), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_18), .A2(n_301), .B1(n_376), .B2(n_381), .Y(n_375) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_18), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g1764 ( .A1(n_19), .A2(n_310), .B1(n_912), .B2(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1783 ( .A(n_19), .Y(n_1783) );
INVx1_ASAP7_75t_L g973 ( .A(n_20), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_20), .A2(n_44), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1032 ( .A1(n_21), .A2(n_109), .B1(n_936), .B2(n_937), .C(n_1033), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_21), .A2(n_109), .B1(n_912), .B2(n_1061), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1432 ( .A(n_22), .Y(n_1432) );
AOI221xp5_ASAP7_75t_L g1454 ( .A1(n_22), .A2(n_293), .B1(n_647), .B2(n_757), .C(n_916), .Y(n_1454) );
INVxp33_ASAP7_75t_L g965 ( .A(n_23), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_23), .A2(n_66), .B1(n_997), .B2(n_998), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_24), .A2(n_298), .B1(n_773), .B2(n_826), .Y(n_825) );
INVxp67_ASAP7_75t_SL g877 ( .A(n_24), .Y(n_877) );
INVx1_ASAP7_75t_L g1354 ( .A(n_25), .Y(n_1354) );
INVx1_ASAP7_75t_L g318 ( .A(n_26), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g1494 ( .A1(n_27), .A2(n_100), .B1(n_1476), .B2(n_1484), .Y(n_1494) );
INVx1_ASAP7_75t_L g1526 ( .A(n_28), .Y(n_1526) );
INVx1_ASAP7_75t_L g1772 ( .A(n_29), .Y(n_1772) );
AOI22xp33_ASAP7_75t_L g1791 ( .A1(n_29), .A2(n_278), .B1(n_488), .B2(n_860), .Y(n_1791) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_30), .A2(n_170), .B1(n_707), .B2(n_713), .C(n_717), .Y(n_970) );
OAI33xp33_ASAP7_75t_L g1003 ( .A1(n_30), .A2(n_170), .A3(n_432), .B1(n_752), .B2(n_1004), .B3(n_1801), .Y(n_1003) );
INVx1_ASAP7_75t_L g1188 ( .A(n_31), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_32), .A2(n_52), .B1(n_381), .B2(n_912), .Y(n_911) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_32), .A2(n_52), .B1(n_936), .B2(n_937), .C(n_938), .Y(n_935) );
AOI21xp33_ASAP7_75t_L g1388 ( .A1(n_33), .A2(n_626), .B(n_1011), .Y(n_1388) );
AOI221xp5_ASAP7_75t_L g1406 ( .A1(n_33), .A2(n_75), .B1(n_461), .B2(n_492), .C(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g399 ( .A(n_34), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_34), .A2(n_260), .B1(n_449), .B2(n_459), .C(n_466), .Y(n_448) );
INVx1_ASAP7_75t_L g807 ( .A(n_35), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_36), .A2(n_296), .B1(n_452), .B2(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_36), .A2(n_213), .B1(n_601), .B2(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g1778 ( .A(n_37), .Y(n_1778) );
AOI22xp33_ASAP7_75t_L g1788 ( .A1(n_37), .A2(n_285), .B1(n_495), .B2(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_L g1714 ( .A(n_38), .Y(n_1714) );
AOI22xp33_ASAP7_75t_L g1731 ( .A1(n_38), .A2(n_254), .B1(n_565), .B2(n_1732), .Y(n_1731) );
OAI222xp33_ASAP7_75t_L g1094 ( .A1(n_39), .A2(n_155), .B1(n_237), .B2(n_1095), .C1(n_1097), .C2(n_1098), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g1128 ( .A1(n_39), .A2(n_155), .B1(n_1129), .B2(n_1131), .C(n_1132), .Y(n_1128) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_40), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g1139 ( .A(n_41), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_42), .A2(n_62), .B1(n_1488), .B2(n_1492), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g639 ( .A(n_43), .Y(n_639) );
INVx1_ASAP7_75t_L g978 ( .A(n_44), .Y(n_978) );
INVxp67_ASAP7_75t_SL g1431 ( .A(n_45), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_45), .A2(n_187), .B1(n_909), .B2(n_1456), .Y(n_1455) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_46), .A2(n_98), .B1(n_707), .B2(n_712), .C(n_717), .Y(n_706) );
OAI221xp5_ASAP7_75t_SL g749 ( .A1(n_46), .A2(n_98), .B1(n_750), .B2(n_751), .C(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g983 ( .A(n_48), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_49), .A2(n_175), .B1(n_832), .B2(n_833), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_49), .A2(n_175), .B1(n_892), .B2(n_894), .Y(n_891) );
INVxp33_ASAP7_75t_L g1042 ( .A(n_50), .Y(n_1042) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_51), .A2(n_83), .B1(n_757), .B2(n_916), .C(n_1199), .Y(n_1198) );
INVxp67_ASAP7_75t_L g1231 ( .A(n_51), .Y(n_1231) );
INVx1_ASAP7_75t_L g545 ( .A(n_53), .Y(n_545) );
INVx1_ASAP7_75t_L g678 ( .A(n_54), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_55), .A2(n_135), .B1(n_551), .B2(n_554), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_55), .A2(n_189), .B1(n_569), .B2(n_570), .C(n_573), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_56), .A2(n_180), .B1(n_386), .B2(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_56), .A2(n_180), .B1(n_488), .B2(n_490), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_57), .A2(n_182), .B1(n_1476), .B2(n_1484), .Y(n_1512) );
OAI221xp5_ASAP7_75t_L g1383 ( .A1(n_58), .A2(n_123), .B1(n_606), .B2(n_1004), .C(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1411 ( .A(n_58), .Y(n_1411) );
AO22x1_ASAP7_75t_SL g1551 ( .A1(n_59), .A2(n_106), .B1(n_1476), .B2(n_1484), .Y(n_1551) );
AOI221xp5_ASAP7_75t_L g1362 ( .A1(n_60), .A2(n_181), .B1(n_1119), .B2(n_1363), .C(n_1365), .Y(n_1362) );
INVx1_ASAP7_75t_L g960 ( .A(n_61), .Y(n_960) );
XOR2x2_ASAP7_75t_L g782 ( .A(n_62), .B(n_783), .Y(n_782) );
INVxp33_ASAP7_75t_L g968 ( .A(n_63), .Y(n_968) );
AOI21xp33_ASAP7_75t_L g1000 ( .A1(n_63), .A2(n_593), .B(n_1001), .Y(n_1000) );
INVxp33_ASAP7_75t_L g801 ( .A(n_64), .Y(n_801) );
INVx1_ASAP7_75t_L g1205 ( .A(n_65), .Y(n_1205) );
INVxp33_ASAP7_75t_L g969 ( .A(n_66), .Y(n_969) );
XNOR2x2_ASAP7_75t_L g614 ( .A(n_67), .B(n_615), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g1513 ( .A1(n_67), .A2(n_202), .B1(n_1492), .B2(n_1514), .Y(n_1513) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_68), .A2(n_232), .B1(n_826), .B2(n_1305), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_68), .A2(n_232), .B1(n_1143), .B2(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g532 ( .A(n_69), .Y(n_532) );
OAI211xp5_ASAP7_75t_SL g1719 ( .A1(n_70), .A2(n_1449), .B(n_1720), .C(n_1723), .Y(n_1719) );
AOI22xp33_ASAP7_75t_L g1735 ( .A1(n_70), .A2(n_167), .B1(n_885), .B2(n_1129), .Y(n_1735) );
CKINVDCx5p33_ASAP7_75t_R g1158 ( .A(n_71), .Y(n_1158) );
AOI221xp5_ASAP7_75t_L g903 ( .A1(n_72), .A2(n_302), .B1(n_904), .B2(n_905), .C(n_906), .Y(n_903) );
INVxp33_ASAP7_75t_L g931 ( .A(n_72), .Y(n_931) );
INVxp33_ASAP7_75t_L g1031 ( .A(n_73), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_73), .A2(n_311), .B1(n_909), .B2(n_1059), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_74), .A2(n_157), .B1(n_492), .B2(n_1149), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_74), .A2(n_157), .B1(n_583), .B2(n_1181), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_75), .A2(n_205), .B1(n_572), .B2(n_998), .Y(n_1387) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_76), .A2(n_158), .B1(n_827), .B2(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1372 ( .A(n_76), .Y(n_1372) );
INVxp33_ASAP7_75t_SL g437 ( .A(n_77), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_77), .A2(n_299), .B1(n_490), .B2(n_494), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g1517 ( .A1(n_78), .A2(n_94), .B1(n_1492), .B2(n_1514), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_79), .A2(n_261), .B1(n_918), .B2(n_919), .Y(n_917) );
INVxp67_ASAP7_75t_SL g951 ( .A(n_79), .Y(n_951) );
INVx1_ASAP7_75t_L g1463 ( .A(n_80), .Y(n_1463) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_81), .A2(n_200), .B1(n_908), .B2(n_909), .Y(n_907) );
INVxp33_ASAP7_75t_SL g934 ( .A(n_81), .Y(n_934) );
OR2x2_ASAP7_75t_L g347 ( .A(n_82), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g351 ( .A(n_82), .Y(n_351) );
BUFx2_ASAP7_75t_L g446 ( .A(n_82), .Y(n_446) );
INVx1_ASAP7_75t_L g456 ( .A(n_82), .Y(n_456) );
INVxp33_ASAP7_75t_SL g1229 ( .A(n_83), .Y(n_1229) );
AOI22xp33_ASAP7_75t_SL g1150 ( .A1(n_84), .A2(n_97), .B1(n_1142), .B2(n_1143), .Y(n_1150) );
INVx1_ASAP7_75t_L g1179 ( .A(n_84), .Y(n_1179) );
INVx1_ASAP7_75t_L g1528 ( .A(n_85), .Y(n_1528) );
INVxp67_ASAP7_75t_L g1263 ( .A(n_86), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_87), .A2(n_258), .B1(n_1476), .B2(n_1484), .Y(n_1538) );
AOI221xp5_ASAP7_75t_SL g1347 ( .A1(n_88), .A2(n_93), .B1(n_426), .B2(n_906), .C(n_1082), .Y(n_1347) );
INVx1_ASAP7_75t_L g1361 ( .A(n_88), .Y(n_1361) );
INVxp33_ASAP7_75t_L g1297 ( .A(n_89), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_89), .A2(n_268), .B1(n_826), .B2(n_904), .Y(n_1311) );
INVx1_ASAP7_75t_L g1343 ( .A(n_90), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_91), .A2(n_222), .B1(n_1488), .B2(n_1492), .Y(n_1495) );
INVx1_ASAP7_75t_L g733 ( .A(n_92), .Y(n_733) );
INVx1_ASAP7_75t_L g1359 ( .A(n_93), .Y(n_1359) );
XOR2x2_ASAP7_75t_L g1375 ( .A(n_94), .B(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1213 ( .A(n_95), .Y(n_1213) );
INVxp67_ASAP7_75t_SL g979 ( .A(n_96), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_96), .A2(n_266), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_97), .B(n_436), .Y(n_1164) );
INVxp33_ASAP7_75t_L g1290 ( .A(n_99), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_99), .A2(n_244), .B1(n_1015), .B2(n_1087), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_101), .Y(n_745) );
INVx1_ASAP7_75t_L g1554 ( .A(n_102), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_103), .A2(n_225), .B1(n_629), .B2(n_822), .Y(n_1393) );
OAI211xp5_ASAP7_75t_L g1395 ( .A1(n_103), .A2(n_1396), .B(n_1397), .C(n_1399), .Y(n_1395) );
OAI22xp33_ASAP7_75t_SL g645 ( .A1(n_104), .A2(n_134), .B1(n_574), .B2(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g683 ( .A(n_104), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g1350 ( .A1(n_107), .A2(n_164), .B1(n_391), .B2(n_757), .C(n_916), .Y(n_1350) );
AOI221xp5_ASAP7_75t_L g1368 ( .A1(n_107), .A2(n_158), .B1(n_1369), .B2(n_1370), .C(n_1371), .Y(n_1368) );
XNOR2x1_ASAP7_75t_L g1022 ( .A(n_108), .B(n_1023), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_110), .Y(n_632) );
INVx1_ASAP7_75t_L g598 ( .A(n_111), .Y(n_598) );
OAI222xp33_ASAP7_75t_L g1099 ( .A1(n_112), .A2(n_172), .B1(n_294), .B2(n_1100), .C1(n_1101), .C2(n_1102), .Y(n_1099) );
INVx1_ASAP7_75t_L g1114 ( .A(n_112), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g1722 ( .A(n_113), .Y(n_1722) );
OAI22xp33_ASAP7_75t_L g1380 ( .A1(n_114), .A2(n_274), .B1(n_387), .B2(n_606), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_114), .A2(n_162), .B1(n_861), .B2(n_1360), .Y(n_1405) );
AOI221xp5_ASAP7_75t_L g1773 ( .A1(n_115), .A2(n_271), .B1(n_580), .B2(n_640), .C(n_1774), .Y(n_1773) );
AOI22xp33_ASAP7_75t_L g1787 ( .A1(n_115), .A2(n_196), .B1(n_495), .B2(n_954), .Y(n_1787) );
AOI21xp5_ASAP7_75t_L g1394 ( .A1(n_116), .A2(n_593), .B(n_1001), .Y(n_1394) );
INVx1_ASAP7_75t_L g1400 ( .A(n_116), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_117), .A2(n_162), .B1(n_601), .B2(n_646), .Y(n_1379) );
AOI22xp5_ASAP7_75t_L g1404 ( .A1(n_117), .A2(n_274), .B1(n_470), .B2(n_1146), .Y(n_1404) );
OAI221xp5_ASAP7_75t_L g1425 ( .A1(n_118), .A2(n_154), .B1(n_714), .B2(n_936), .C(n_1033), .Y(n_1425) );
OAI22xp33_ASAP7_75t_L g1461 ( .A1(n_118), .A2(n_154), .B1(n_1102), .B2(n_1462), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_119), .A2(n_267), .B1(n_391), .B2(n_417), .C(n_421), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_119), .A2(n_267), .B1(n_494), .B2(n_496), .Y(n_493) );
INVx1_ASAP7_75t_L g535 ( .A(n_120), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g1718 ( .A1(n_121), .A2(n_580), .B(n_584), .Y(n_1718) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_121), .A2(n_149), .B1(n_1129), .B2(n_1734), .Y(n_1733) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_122), .Y(n_1386) );
INVx1_ASAP7_75t_L g1398 ( .A(n_123), .Y(n_1398) );
INVx1_ASAP7_75t_L g1345 ( .A(n_124), .Y(n_1345) );
OAI22xp33_ASAP7_75t_L g1728 ( .A1(n_125), .A2(n_167), .B1(n_436), .B2(n_439), .Y(n_1728) );
AOI22xp33_ASAP7_75t_L g1736 ( .A1(n_125), .A2(n_228), .B1(n_565), .B2(n_1142), .Y(n_1736) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_126), .A2(n_265), .B1(n_418), .B2(n_580), .C(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1126 ( .A(n_126), .Y(n_1126) );
INVx1_ASAP7_75t_L g696 ( .A(n_127), .Y(n_696) );
INVx1_ASAP7_75t_L g1265 ( .A(n_128), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_128), .A2(n_252), .B1(n_1284), .B2(n_1286), .Y(n_1283) );
INVxp33_ASAP7_75t_SL g434 ( .A(n_129), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_129), .A2(n_247), .B1(n_488), .B2(n_496), .Y(n_499) );
INVx1_ASAP7_75t_L g1047 ( .A(n_130), .Y(n_1047) );
INVx1_ASAP7_75t_L g1480 ( .A(n_131), .Y(n_1480) );
CKINVDCx5p33_ASAP7_75t_R g1721 ( .A(n_132), .Y(n_1721) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_133), .Y(n_991) );
INVx1_ASAP7_75t_L g673 ( .A(n_134), .Y(n_673) );
INVx1_ASAP7_75t_L g576 ( .A(n_135), .Y(n_576) );
INVx1_ASAP7_75t_L g1167 ( .A(n_136), .Y(n_1167) );
AOI221xp5_ASAP7_75t_L g1522 ( .A1(n_137), .A2(n_210), .B1(n_1523), .B2(n_1524), .C(n_1525), .Y(n_1522) );
INVx1_ASAP7_75t_L g966 ( .A(n_138), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_138), .B(n_401), .Y(n_1002) );
INVx1_ASAP7_75t_L g736 ( .A(n_139), .Y(n_736) );
INVx1_ASAP7_75t_L g813 ( .A(n_140), .Y(n_813) );
INVx1_ASAP7_75t_L g1049 ( .A(n_141), .Y(n_1049) );
INVx1_ASAP7_75t_L g1481 ( .A(n_142), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_142), .B(n_1479), .Y(n_1486) );
XNOR2xp5_ASAP7_75t_L g1758 ( .A(n_143), .B(n_1759), .Y(n_1758) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_144), .A2(n_211), .B1(n_908), .B2(n_919), .Y(n_1348) );
OAI221xp5_ASAP7_75t_L g1357 ( .A1(n_144), .A2(n_211), .B1(n_724), .B2(n_857), .C(n_1358), .Y(n_1357) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_145), .A2(n_168), .B1(n_821), .B2(n_823), .Y(n_820) );
INVxp67_ASAP7_75t_SL g874 ( .A(n_145), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g1775 ( .A1(n_146), .A2(n_196), .B1(n_758), .B2(n_1085), .Y(n_1775) );
AOI22xp33_ASAP7_75t_SL g1785 ( .A1(n_146), .A2(n_271), .B1(n_1360), .B2(n_1786), .Y(n_1785) );
AOI21xp5_ASAP7_75t_L g1770 ( .A1(n_147), .A2(n_406), .B(n_1202), .Y(n_1770) );
INVx1_ASAP7_75t_L g1795 ( .A(n_147), .Y(n_1795) );
INVx2_ASAP7_75t_L g330 ( .A(n_148), .Y(n_330) );
INVx1_ASAP7_75t_L g1715 ( .A(n_149), .Y(n_1715) );
OAI22x1_ASAP7_75t_SL g1239 ( .A1(n_150), .A2(n_1240), .B1(n_1326), .B2(n_1327), .Y(n_1239) );
INVx1_ASAP7_75t_L g1326 ( .A(n_150), .Y(n_1326) );
AO221x2_ASAP7_75t_L g1498 ( .A1(n_150), .A2(n_191), .B1(n_1488), .B2(n_1499), .C(n_1501), .Y(n_1498) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_151), .A2(n_286), .B1(n_370), .B2(n_915), .C(n_916), .Y(n_914) );
INVxp33_ASAP7_75t_SL g944 ( .A(n_151), .Y(n_944) );
INVx1_ASAP7_75t_L g755 ( .A(n_152), .Y(n_755) );
BUFx3_ASAP7_75t_L g360 ( .A(n_153), .Y(n_360) );
INVx1_ASAP7_75t_L g390 ( .A(n_153), .Y(n_390) );
INVx1_ASAP7_75t_L g792 ( .A(n_156), .Y(n_792) );
INVx1_ASAP7_75t_L g985 ( .A(n_159), .Y(n_985) );
INVxp33_ASAP7_75t_L g1423 ( .A(n_160), .Y(n_1423) );
AOI221xp5_ASAP7_75t_L g1459 ( .A1(n_160), .A2(n_201), .B1(n_418), .B2(n_593), .C(n_1001), .Y(n_1459) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_161), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_163), .Y(n_1217) );
INVx1_ASAP7_75t_L g1373 ( .A(n_164), .Y(n_1373) );
INVxp67_ASAP7_75t_L g721 ( .A(n_165), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_165), .A2(n_284), .B1(n_425), .B2(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g703 ( .A(n_166), .Y(n_703) );
INVxp67_ASAP7_75t_SL g883 ( .A(n_168), .Y(n_883) );
INVx1_ASAP7_75t_L g1344 ( .A(n_169), .Y(n_1344) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_171), .Y(n_841) );
INVx1_ASAP7_75t_L g1107 ( .A(n_172), .Y(n_1107) );
INVxp33_ASAP7_75t_SL g526 ( .A(n_173), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_173), .A2(n_217), .B1(n_569), .B2(n_582), .C(n_585), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_174), .A2(n_256), .B1(n_832), .B2(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1113 ( .A(n_174), .Y(n_1113) );
INVxp67_ASAP7_75t_L g1040 ( .A(n_176), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_176), .A2(n_224), .B1(n_905), .B2(n_909), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1214 ( .A1(n_177), .A2(n_272), .B1(n_406), .B2(n_757), .C(n_758), .Y(n_1214) );
INVxp33_ASAP7_75t_SL g1223 ( .A(n_177), .Y(n_1223) );
INVx1_ASAP7_75t_L g355 ( .A(n_178), .Y(n_355) );
INVx1_ASAP7_75t_L g408 ( .A(n_178), .Y(n_408) );
INVxp33_ASAP7_75t_L g1260 ( .A(n_179), .Y(n_1260) );
INVx1_ASAP7_75t_L g1342 ( .A(n_181), .Y(n_1342) );
INVxp33_ASAP7_75t_SL g1420 ( .A(n_183), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g1460 ( .A1(n_183), .A2(n_188), .B1(n_391), .B2(n_603), .Y(n_1460) );
INVx1_ASAP7_75t_L g982 ( .A(n_184), .Y(n_982) );
INVx1_ASAP7_75t_L g1207 ( .A(n_185), .Y(n_1207) );
OAI221xp5_ASAP7_75t_L g1224 ( .A1(n_185), .A2(n_212), .B1(n_936), .B2(n_937), .C(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g910 ( .A(n_186), .Y(n_910) );
INVx1_ASAP7_75t_L g1437 ( .A(n_187), .Y(n_1437) );
INVxp33_ASAP7_75t_SL g1424 ( .A(n_188), .Y(n_1424) );
INVx1_ASAP7_75t_L g549 ( .A(n_189), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g1390 ( .A(n_190), .Y(n_1390) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_192), .A2(n_275), .B1(n_626), .B2(n_628), .C(n_630), .Y(n_625) );
INVx1_ASAP7_75t_L g688 ( .A(n_192), .Y(n_688) );
INVx1_ASAP7_75t_L g1044 ( .A(n_193), .Y(n_1044) );
AOI22xp33_ASAP7_75t_SL g828 ( .A1(n_194), .A2(n_243), .B1(n_823), .B2(n_829), .Y(n_828) );
OAI211xp5_ASAP7_75t_SL g851 ( .A1(n_194), .A2(n_852), .B(n_856), .C(n_865), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g1516 ( .A1(n_195), .A2(n_231), .B1(n_1476), .B2(n_1484), .Y(n_1516) );
AOI22xp5_ASAP7_75t_L g1539 ( .A1(n_197), .A2(n_257), .B1(n_1492), .B2(n_1514), .Y(n_1539) );
AOI221xp5_ASAP7_75t_L g1081 ( .A1(n_198), .A2(n_270), .B1(n_426), .B2(n_906), .C(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1111 ( .A(n_198), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1726 ( .A1(n_199), .A2(n_235), .B1(n_370), .B2(n_629), .Y(n_1726) );
OAI22xp5_ASAP7_75t_L g1741 ( .A1(n_199), .A2(n_306), .B1(n_1742), .B2(n_1743), .Y(n_1741) );
INVxp33_ASAP7_75t_L g929 ( .A(n_200), .Y(n_929) );
INVxp33_ASAP7_75t_L g1421 ( .A(n_201), .Y(n_1421) );
INVx1_ASAP7_75t_L g1052 ( .A(n_203), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_204), .Y(n_1138) );
INVx1_ASAP7_75t_L g1408 ( .A(n_205), .Y(n_1408) );
INVx1_ASAP7_75t_L g1555 ( .A(n_206), .Y(n_1555) );
INVx1_ASAP7_75t_L g1162 ( .A(n_207), .Y(n_1162) );
OAI211xp5_ASAP7_75t_L g1177 ( .A1(n_207), .A2(n_1100), .B(n_1178), .C(n_1182), .Y(n_1177) );
CKINVDCx20_ASAP7_75t_R g1502 ( .A(n_208), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_209), .A2(n_253), .B1(n_833), .B2(n_1201), .Y(n_1200) );
INVxp67_ASAP7_75t_L g1228 ( .A(n_209), .Y(n_1228) );
INVx1_ASAP7_75t_L g1208 ( .A(n_212), .Y(n_1208) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_213), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_214), .Y(n_1054) );
XNOR2x1_ASAP7_75t_L g1077 ( .A(n_215), .B(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1204 ( .A(n_216), .Y(n_1204) );
INVxp33_ASAP7_75t_SL g530 ( .A(n_217), .Y(n_530) );
INVx1_ASAP7_75t_L g734 ( .A(n_218), .Y(n_734) );
BUFx3_ASAP7_75t_L g362 ( .A(n_219), .Y(n_362) );
INVx1_ASAP7_75t_L g372 ( .A(n_219), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_220), .Y(n_622) );
AOI21xp33_ASAP7_75t_L g1727 ( .A1(n_221), .A2(n_634), .B(n_799), .Y(n_1727) );
INVx1_ASAP7_75t_L g1739 ( .A(n_221), .Y(n_1739) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_223), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_223), .B(n_290), .Y(n_348) );
AND2x2_ASAP7_75t_L g457 ( .A(n_223), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g507 ( .A(n_223), .Y(n_507) );
INVxp67_ASAP7_75t_L g1038 ( .A(n_224), .Y(n_1038) );
INVx1_ASAP7_75t_L g1401 ( .A(n_225), .Y(n_1401) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_226), .A2(n_401), .B(n_405), .Y(n_400) );
INVx1_ASAP7_75t_L g474 ( .A(n_226), .Y(n_474) );
INVx1_ASAP7_75t_L g923 ( .A(n_227), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g1712 ( .A1(n_228), .A2(n_1176), .B1(n_1453), .B2(n_1713), .C(n_1716), .Y(n_1712) );
INVx1_ASAP7_75t_L g597 ( .A(n_229), .Y(n_597) );
INVx2_ASAP7_75t_L g357 ( .A(n_230), .Y(n_357) );
OR2x2_ASAP7_75t_L g374 ( .A(n_230), .B(n_355), .Y(n_374) );
INVx1_ASAP7_75t_L g1793 ( .A(n_233), .Y(n_1793) );
INVx1_ASAP7_75t_L g1216 ( .A(n_234), .Y(n_1216) );
INVx1_ASAP7_75t_L g1740 ( .A(n_235), .Y(n_1740) );
INVxp67_ASAP7_75t_L g726 ( .A(n_236), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_236), .A2(n_283), .B1(n_766), .B2(n_767), .C(n_771), .Y(n_765) );
INVx1_ASAP7_75t_L g1133 ( .A(n_237), .Y(n_1133) );
CKINVDCx16_ASAP7_75t_R g1334 ( .A(n_238), .Y(n_1334) );
INVx1_ASAP7_75t_L g1440 ( .A(n_239), .Y(n_1440) );
INVx1_ASAP7_75t_L g1779 ( .A(n_240), .Y(n_1779) );
INVx1_ASAP7_75t_L g924 ( .A(n_241), .Y(n_924) );
INVx1_ASAP7_75t_L g1197 ( .A(n_242), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g870 ( .A1(n_243), .A2(n_871), .B1(n_873), .B2(n_880), .C(n_890), .Y(n_870) );
INVxp67_ASAP7_75t_L g1294 ( .A(n_244), .Y(n_1294) );
INVx1_ASAP7_75t_L g1256 ( .A(n_245), .Y(n_1256) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_246), .A2(n_269), .B1(n_909), .B2(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1124 ( .A(n_246), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_247), .Y(n_415) );
INVx1_ASAP7_75t_L g739 ( .A(n_248), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_249), .A2(n_260), .B1(n_386), .B2(n_391), .C(n_392), .Y(n_385) );
INVxp33_ASAP7_75t_L g467 ( .A(n_249), .Y(n_467) );
INVx1_ASAP7_75t_L g1211 ( .A(n_250), .Y(n_1211) );
INVx1_ASAP7_75t_L g958 ( .A(n_251), .Y(n_958) );
INVx1_ASAP7_75t_L g1270 ( .A(n_252), .Y(n_1270) );
INVxp67_ASAP7_75t_L g1233 ( .A(n_253), .Y(n_1233) );
INVx1_ASAP7_75t_L g1717 ( .A(n_254), .Y(n_1717) );
INVx1_ASAP7_75t_L g1153 ( .A(n_255), .Y(n_1153) );
AOI21xp5_ASAP7_75t_L g1175 ( .A1(n_255), .A2(n_572), .B(n_634), .Y(n_1175) );
INVx1_ASAP7_75t_L g1109 ( .A(n_256), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1708 ( .A1(n_258), .A2(n_1709), .B1(n_1744), .B2(n_1745), .Y(n_1708) );
INVxp67_ASAP7_75t_SL g1744 ( .A(n_258), .Y(n_1744) );
AOI22xp33_ASAP7_75t_L g1752 ( .A1(n_258), .A2(n_1753), .B1(n_1757), .B2(n_1797), .Y(n_1752) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_259), .A2(n_277), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_259), .A2(n_277), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
INVxp33_ASAP7_75t_L g941 ( .A(n_261), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_262), .Y(n_621) );
INVx1_ASAP7_75t_L g987 ( .A(n_263), .Y(n_987) );
INVx1_ASAP7_75t_L g1157 ( .A(n_264), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1118 ( .A1(n_265), .A2(n_269), .B1(n_1119), .B2(n_1121), .C(n_1123), .Y(n_1118) );
INVxp33_ASAP7_75t_L g974 ( .A(n_266), .Y(n_974) );
INVxp67_ASAP7_75t_L g1277 ( .A(n_268), .Y(n_1277) );
INVx1_ASAP7_75t_L g1117 ( .A(n_270), .Y(n_1117) );
INVxp33_ASAP7_75t_SL g1221 ( .A(n_272), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_273), .Y(n_1093) );
INVx1_ASAP7_75t_L g690 ( .A(n_275), .Y(n_690) );
INVx1_ASAP7_75t_L g925 ( .A(n_276), .Y(n_925) );
INVx1_ASAP7_75t_L g1777 ( .A(n_278), .Y(n_1777) );
INVx1_ASAP7_75t_L g1415 ( .A(n_279), .Y(n_1415) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_280), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_280), .B(n_318), .Y(n_1483) );
AND3x2_ASAP7_75t_L g1491 ( .A(n_280), .B(n_318), .C(n_1480), .Y(n_1491) );
INVx2_ASAP7_75t_L g331 ( .A(n_281), .Y(n_331) );
XNOR2x2_ASAP7_75t_L g522 ( .A(n_282), .B(n_523), .Y(n_522) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_283), .Y(n_730) );
INVxp33_ASAP7_75t_SL g723 ( .A(n_284), .Y(n_723) );
INVx1_ASAP7_75t_L g1763 ( .A(n_285), .Y(n_1763) );
INVxp67_ASAP7_75t_SL g947 ( .A(n_286), .Y(n_947) );
INVx1_ASAP7_75t_L g528 ( .A(n_287), .Y(n_528) );
INVx1_ASAP7_75t_L g1443 ( .A(n_288), .Y(n_1443) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_289), .Y(n_654) );
INVx1_ASAP7_75t_L g333 ( .A(n_290), .Y(n_333) );
INVx2_ASAP7_75t_L g458 ( .A(n_290), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_291), .Y(n_652) );
OR2x2_ASAP7_75t_L g1710 ( .A(n_292), .B(n_345), .Y(n_1710) );
INVxp67_ASAP7_75t_SL g1436 ( .A(n_293), .Y(n_1436) );
INVx1_ASAP7_75t_L g1106 ( .A(n_294), .Y(n_1106) );
INVxp33_ASAP7_75t_L g1030 ( .A(n_295), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_295), .A2(n_297), .B1(n_426), .B2(n_904), .C(n_906), .Y(n_1057) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_296), .A2(n_305), .B1(n_605), .B2(n_606), .Y(n_604) );
INVxp33_ASAP7_75t_L g1028 ( .A(n_297), .Y(n_1028) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_298), .Y(n_889) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_299), .Y(n_366) );
INVx1_ASAP7_75t_L g1441 ( .A(n_300), .Y(n_1441) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_301), .Y(n_513) );
INVxp33_ASAP7_75t_L g933 ( .A(n_302), .Y(n_933) );
INVx1_ASAP7_75t_L g671 ( .A(n_303), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_304), .Y(n_363) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_305), .Y(n_561) );
INVx1_ASAP7_75t_L g1724 ( .A(n_306), .Y(n_1724) );
INVx1_ASAP7_75t_L g1444 ( .A(n_307), .Y(n_1444) );
INVxp33_ASAP7_75t_SL g702 ( .A(n_308), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g1769 ( .A(n_309), .Y(n_1769) );
INVx1_ASAP7_75t_L g1782 ( .A(n_310), .Y(n_1782) );
INVxp33_ASAP7_75t_L g1027 ( .A(n_311), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_334), .B(n_1465), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g1751 ( .A(n_316), .B(n_322), .Y(n_1751) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_SL g1756 ( .A(n_317), .Y(n_1756) );
NAND2xp5_ASAP7_75t_L g1799 ( .A(n_317), .B(n_319), .Y(n_1799) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g1755 ( .A(n_319), .B(n_1756), .Y(n_1755) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_324), .B(n_351), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g486 ( .A(n_325), .B(n_333), .Y(n_486) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g538 ( .A(n_326), .B(n_539), .Y(n_538) );
INVx8_ASAP7_75t_L g1296 ( .A(n_327), .Y(n_1296) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
OR2x2_ASAP7_75t_L g346 ( .A(n_328), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g661 ( .A(n_328), .Y(n_661) );
INVx2_ASAP7_75t_SL g876 ( .A(n_328), .Y(n_876) );
BUFx6f_ASAP7_75t_L g943 ( .A(n_328), .Y(n_943) );
INVx2_ASAP7_75t_SL g977 ( .A(n_328), .Y(n_977) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_328), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1132 ( .A1(n_328), .A2(n_681), .B1(n_1093), .B2(n_1133), .Y(n_1132) );
OR2x6_ASAP7_75t_L g1299 ( .A(n_328), .B(n_1289), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_328), .A2(n_681), .B1(n_1386), .B2(n_1408), .Y(n_1407) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g454 ( .A(n_330), .B(n_331), .Y(n_454) );
INVx2_ASAP7_75t_L g463 ( .A(n_330), .Y(n_463) );
AND2x4_ASAP7_75t_L g472 ( .A(n_330), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g479 ( .A(n_330), .Y(n_479) );
INVx1_ASAP7_75t_L g517 ( .A(n_330), .Y(n_517) );
INVx1_ASAP7_75t_L g465 ( .A(n_331), .Y(n_465) );
INVx2_ASAP7_75t_L g473 ( .A(n_331), .Y(n_473) );
INVx1_ASAP7_75t_L g511 ( .A(n_331), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_331), .B(n_463), .Y(n_544) );
INVx1_ASAP7_75t_L g666 ( .A(n_331), .Y(n_666) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_332), .B(n_511), .Y(n_1285) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_333), .B(n_516), .Y(n_1286) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_1329), .B1(n_1330), .B2(n_1464), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_1070), .B2(n_1071), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g1464 ( .A1(n_336), .A2(n_337), .B1(n_1070), .B2(n_1071), .Y(n_1464) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AO22x2_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_779), .B1(n_1068), .B2(n_1069), .Y(n_337) );
INVx1_ASAP7_75t_L g1069 ( .A(n_338), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_694), .B1(n_695), .B2(n_778), .Y(n_338) );
INVx2_ASAP7_75t_L g778 ( .A(n_339), .Y(n_778) );
AO22x2_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_520), .B1(n_521), .B2(n_693), .Y(n_339) );
INVx2_ASAP7_75t_SL g693 ( .A(n_340), .Y(n_693) );
XNOR2x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_447), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_363), .B(n_364), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g1445 ( .A1(n_344), .A2(n_442), .B1(n_1446), .B2(n_1463), .Y(n_1445) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx5_ASAP7_75t_L g744 ( .A(n_345), .Y(n_744) );
INVx1_ASAP7_75t_L g990 ( .A(n_345), .Y(n_990) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
INVx2_ASAP7_75t_L g533 ( .A(n_346), .Y(n_533) );
INVx3_ASAP7_75t_L g512 ( .A(n_347), .Y(n_512) );
INVx1_ASAP7_75t_L g848 ( .A(n_348), .Y(n_848) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x6_ASAP7_75t_L g842 ( .A(n_350), .B(n_843), .Y(n_842) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x4_ASAP7_75t_L g835 ( .A(n_351), .B(n_407), .Y(n_835) );
INVx2_ASAP7_75t_L g1100 ( .A(n_352), .Y(n_1100) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_358), .Y(n_352) );
AND2x4_ASAP7_75t_L g377 ( .A(n_353), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g382 ( .A(n_353), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g432 ( .A(n_353), .Y(n_432) );
BUFx2_ASAP7_75t_L g595 ( .A(n_353), .Y(n_595) );
AND2x4_ASAP7_75t_L g651 ( .A(n_353), .B(n_378), .Y(n_651) );
AND2x4_ASAP7_75t_L g653 ( .A(n_353), .B(n_383), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g812 ( .A(n_353), .B(n_504), .Y(n_812) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_353), .B(n_383), .Y(n_1766) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g407 ( .A(n_356), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g423 ( .A(n_357), .B(n_408), .Y(n_423) );
INVx1_ASAP7_75t_L g1249 ( .A(n_357), .Y(n_1249) );
INVx1_ASAP7_75t_L g1254 ( .A(n_357), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_357), .Y(n_1259) );
INVx6_ASAP7_75t_L g428 ( .A(n_358), .Y(n_428) );
BUFx2_ASAP7_75t_L g593 ( .A(n_358), .Y(n_593) );
INVx2_ASAP7_75t_L g800 ( .A(n_358), .Y(n_800) );
AND2x4_ASAP7_75t_L g1257 ( .A(n_358), .B(n_1258), .Y(n_1257) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g371 ( .A(n_360), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g414 ( .A(n_360), .B(n_362), .Y(n_414) );
INVx1_ASAP7_75t_L g380 ( .A(n_361), .Y(n_380) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g389 ( .A(n_362), .B(n_390), .Y(n_389) );
AOI31xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_409), .A3(n_433), .B(n_441), .Y(n_364) );
AOI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_375), .C(n_385), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g993 ( .A1(n_367), .A2(n_982), .B(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_369), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g902 ( .A1(n_369), .A2(n_903), .B1(n_907), .B2(n_910), .C(n_911), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g1056 ( .A1(n_369), .A2(n_1044), .B1(n_1057), .B2(n_1058), .C(n_1060), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_369), .B(n_1216), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g1776 ( .A1(n_369), .A2(n_435), .B1(n_1777), .B2(n_1778), .Y(n_1776) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_373), .Y(n_369) );
INVx2_ASAP7_75t_SL g754 ( .A(n_370), .Y(n_754) );
BUFx3_ASAP7_75t_L g908 ( .A(n_370), .Y(n_908) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g391 ( .A(n_371), .Y(n_391) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_371), .Y(n_578) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_371), .Y(n_584) );
INVx2_ASAP7_75t_SL g627 ( .A(n_371), .Y(n_627) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_371), .Y(n_647) );
BUFx3_ASAP7_75t_L g822 ( .A(n_371), .Y(n_822) );
BUFx2_ASAP7_75t_L g997 ( .A(n_371), .Y(n_997) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_371), .Y(n_1087) );
AND2x6_ASAP7_75t_L g1252 ( .A(n_371), .B(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g398 ( .A(n_372), .Y(n_398) );
AND2x4_ASAP7_75t_L g412 ( .A(n_373), .B(n_413), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_373), .A2(n_600), .B(n_604), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_373), .A2(n_643), .B(n_645), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_373), .A2(n_435), .B1(n_1093), .B2(n_1094), .C(n_1099), .Y(n_1092) );
A2O1A1Ixp33_ASAP7_75t_L g1178 ( .A1(n_373), .A2(n_904), .B(n_1179), .C(n_1180), .Y(n_1178) );
AOI222xp33_ASAP7_75t_L g1337 ( .A1(n_373), .A2(n_377), .B1(n_382), .B2(n_1338), .C1(n_1344), .C2(n_1345), .Y(n_1337) );
OAI21xp5_ASAP7_75t_L g1378 ( .A1(n_373), .A2(n_1379), .B(n_1380), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_373), .B(n_647), .Y(n_1450) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g436 ( .A(n_374), .B(n_396), .Y(n_436) );
OR2x2_ASAP7_75t_L g439 ( .A(n_374), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g791 ( .A(n_374), .B(n_456), .Y(n_791) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_377), .A2(n_382), .B1(n_597), .B2(n_598), .Y(n_596) );
INVx2_ASAP7_75t_SL g750 ( .A(n_377), .Y(n_750) );
INVx2_ASAP7_75t_SL g912 ( .A(n_377), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_377), .A2(n_382), .B1(n_1207), .B2(n_1208), .Y(n_1206) );
INVxp67_ASAP7_75t_L g1004 ( .A(n_378), .Y(n_1004) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g810 ( .A(n_379), .Y(n_810) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g1269 ( .A(n_380), .Y(n_1269) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g752 ( .A(n_383), .Y(n_752) );
INVx1_ASAP7_75t_L g1384 ( .A(n_383), .Y(n_1384) );
BUFx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x6_ASAP7_75t_L g1271 ( .A(n_384), .B(n_1254), .Y(n_1271) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_387), .A2(n_703), .B1(n_754), .B2(n_755), .C(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g1085 ( .A(n_387), .Y(n_1085) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_388), .Y(n_569) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_388), .Y(n_618) );
INVx1_ASAP7_75t_L g774 ( .A(n_388), .Y(n_774) );
INVx1_ASAP7_75t_L g1016 ( .A(n_388), .Y(n_1016) );
AND2x6_ASAP7_75t_L g1261 ( .A(n_388), .B(n_1248), .Y(n_1261) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_389), .Y(n_629) );
INVx1_ASAP7_75t_L g795 ( .A(n_389), .Y(n_795) );
INVx1_ASAP7_75t_L g920 ( .A(n_389), .Y(n_920) );
INVx1_ASAP7_75t_L g397 ( .A(n_390), .Y(n_397) );
OAI21xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_399), .B(n_400), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g601 ( .A(n_395), .Y(n_601) );
INVx2_ASAP7_75t_L g1339 ( .A(n_395), .Y(n_1339) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g589 ( .A(n_396), .Y(n_589) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g404 ( .A(n_397), .B(n_398), .Y(n_404) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g575 ( .A(n_404), .Y(n_575) );
BUFx4f_ASAP7_75t_L g587 ( .A(n_404), .Y(n_587) );
INVx2_ASAP7_75t_L g804 ( .A(n_404), .Y(n_804) );
INVx1_ASAP7_75t_L g1096 ( .A(n_404), .Y(n_1096) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_407), .Y(n_590) );
INVx2_ASAP7_75t_SL g634 ( .A(n_407), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_407), .Y(n_906) );
INVx1_ASAP7_75t_L g1001 ( .A(n_407), .Y(n_1001) );
INVx1_ASAP7_75t_L g1242 ( .A(n_408), .Y(n_1242) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_415), .B1(n_416), .B2(n_424), .C(n_429), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_412), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_412), .A2(n_430), .B1(n_914), .B2(n_917), .C(n_921), .Y(n_913) );
INVx1_ASAP7_75t_L g1007 ( .A(n_412), .Y(n_1007) );
INVx1_ASAP7_75t_L g1196 ( .A(n_412), .Y(n_1196) );
INVx2_ASAP7_75t_SL g1453 ( .A(n_412), .Y(n_1453) );
BUFx3_ASAP7_75t_L g757 ( .A(n_413), .Y(n_757) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_413), .Y(n_824) );
BUFx4f_ASAP7_75t_L g904 ( .A(n_413), .Y(n_904) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_413), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_413), .B(n_595), .Y(n_1091) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_414), .Y(n_420) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g592 ( .A1(n_418), .A2(n_532), .B(n_593), .C(n_594), .Y(n_592) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g430 ( .A(n_419), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g641 ( .A(n_419), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g1341 ( .A1(n_419), .A2(n_647), .B1(n_1342), .B2(n_1343), .Y(n_1341) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g770 ( .A(n_420), .Y(n_770) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_420), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g916 ( .A(n_422), .Y(n_916) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g580 ( .A(n_423), .Y(n_580) );
INVx1_ASAP7_75t_L g624 ( .A(n_423), .Y(n_624) );
INVx2_ASAP7_75t_L g819 ( .A(n_423), .Y(n_819) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g759 ( .A(n_427), .Y(n_759) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g572 ( .A(n_428), .Y(n_572) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_428), .Y(n_638) );
INVx1_ASAP7_75t_L g827 ( .A(n_428), .Y(n_827) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_428), .Y(n_1090) );
INVx2_ASAP7_75t_SL g1170 ( .A(n_428), .Y(n_1170) );
INVx2_ASAP7_75t_L g1202 ( .A(n_428), .Y(n_1202) );
INVx2_ASAP7_75t_L g1250 ( .A(n_428), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g776 ( .A(n_430), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g1005 ( .A1(n_430), .A2(n_987), .B1(n_1006), .B2(n_1008), .C(n_1013), .Y(n_1005) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_430), .A2(n_764), .B1(n_1052), .B2(n_1063), .C(n_1064), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1194 ( .A1(n_430), .A2(n_1195), .B1(n_1197), .B2(n_1198), .C(n_1200), .Y(n_1194) );
AOI21xp33_ASAP7_75t_L g1346 ( .A1(n_430), .A2(n_1347), .B(n_1348), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g1451 ( .A1(n_430), .A2(n_1444), .B1(n_1452), .B2(n_1454), .C(n_1455), .Y(n_1451) );
AOI221xp5_ASAP7_75t_L g1771 ( .A1(n_430), .A2(n_1452), .B1(n_1772), .B2(n_1773), .C(n_1775), .Y(n_1771) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g751 ( .A(n_432), .B(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_435), .A2(n_438), .B1(n_734), .B2(n_736), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_435), .A2(n_438), .B1(n_923), .B2(n_924), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_435), .A2(n_438), .B1(n_983), .B2(n_985), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_435), .A2(n_438), .B1(n_1047), .B2(n_1049), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_435), .A2(n_438), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
AOI22xp5_ASAP7_75t_L g1447 ( .A1(n_435), .A2(n_1440), .B1(n_1443), .B2(n_1448), .Y(n_1447) );
INVx6_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g1458 ( .A1(n_438), .A2(n_1441), .B1(n_1459), .B2(n_1460), .C(n_1461), .Y(n_1458) );
AOI211xp5_ASAP7_75t_L g1762 ( .A1(n_438), .A2(n_1763), .B(n_1764), .C(n_1767), .Y(n_1762) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g603 ( .A(n_440), .Y(n_603) );
INVx2_ASAP7_75t_L g999 ( .A(n_440), .Y(n_999) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx5_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI31xp33_ASAP7_75t_L g746 ( .A1(n_443), .A2(n_747), .A3(n_761), .B(n_777), .Y(n_746) );
OAI31xp33_ASAP7_75t_L g850 ( .A1(n_443), .A2(n_851), .A3(n_870), .B(n_891), .Y(n_850) );
AOI31xp33_ASAP7_75t_L g1055 ( .A1(n_443), .A2(n_1056), .A3(n_1062), .B(n_1065), .Y(n_1055) );
BUFx8_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g900 ( .A(n_444), .Y(n_900) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g655 ( .A(n_445), .Y(n_655) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_445), .B(n_1242), .Y(n_1241) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g485 ( .A(n_446), .Y(n_485) );
OR2x6_ASAP7_75t_L g537 ( .A(n_446), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_480), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_450), .A2(n_632), .B(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_450), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
BUFx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_451), .A2(n_535), .B(n_536), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_451), .A2(n_691), .B1(n_933), .B2(n_934), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_451), .A2(n_531), .B1(n_968), .B2(n_969), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_451), .A2(n_460), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_451), .B(n_1153), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_451), .A2(n_691), .B1(n_1211), .B2(n_1223), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_451), .A2(n_1110), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
AOI221xp5_ASAP7_75t_L g1738 ( .A1(n_451), .A2(n_1110), .B1(n_1739), .B2(n_1740), .C(n_1741), .Y(n_1738) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_451), .A2(n_1110), .B1(n_1795), .B2(n_1796), .Y(n_1794) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
BUFx2_ASAP7_75t_L g1732 ( .A(n_452), .Y(n_1732) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g489 ( .A(n_453), .Y(n_489) );
INVx2_ASAP7_75t_SL g849 ( .A(n_453), .Y(n_849) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_454), .Y(n_553) );
AND2x2_ASAP7_75t_L g460 ( .A(n_455), .B(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g469 ( .A(n_455), .B(n_470), .Y(n_469) );
AND2x6_ASAP7_75t_L g476 ( .A(n_455), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g531 ( .A(n_455), .B(n_461), .Y(n_531) );
AND2x2_ASAP7_75t_L g691 ( .A(n_455), .B(n_461), .Y(n_691) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_455), .B(n_461), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_455), .B(n_849), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_455), .B(n_461), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_455), .B(n_1046), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_455), .A2(n_685), .B1(n_1357), .B2(n_1362), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_455), .B(n_861), .Y(n_1409) );
AND2x4_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g504 ( .A(n_456), .Y(n_504) );
INVx2_ASAP7_75t_L g855 ( .A(n_457), .Y(n_855) );
AND2x4_ASAP7_75t_L g872 ( .A(n_457), .B(n_553), .Y(n_872) );
AND2x2_ASAP7_75t_L g893 ( .A(n_457), .B(n_462), .Y(n_893) );
INVx1_ASAP7_75t_L g506 ( .A(n_458), .Y(n_506) );
INVx1_ASAP7_75t_L g539 ( .A(n_458), .Y(n_539) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g495 ( .A(n_462), .Y(n_495) );
INVx1_ASAP7_75t_L g1120 ( .A(n_462), .Y(n_1120) );
INVx1_ASAP7_75t_L g1130 ( .A(n_462), .Y(n_1130) );
BUFx6f_ASAP7_75t_L g1146 ( .A(n_462), .Y(n_1146) );
BUFx6f_ASAP7_75t_L g1149 ( .A(n_462), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1288 ( .A(n_462), .B(n_1289), .Y(n_1288) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g716 ( .A(n_463), .Y(n_716) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_474), .B2(n_475), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_468), .A2(n_533), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g527 ( .A(n_469), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_469), .A2(n_476), .B1(n_631), .B2(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g705 ( .A(n_469), .Y(n_705) );
BUFx2_ASAP7_75t_L g930 ( .A(n_469), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_469), .A2(n_476), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
BUFx3_ASAP7_75t_L g954 ( .A(n_470), .Y(n_954) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_471), .Y(n_548) );
INVx3_ASAP7_75t_L g1046 ( .A(n_471), .Y(n_1046) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_472), .Y(n_492) );
INVx1_ASAP7_75t_L g888 ( .A(n_472), .Y(n_888) );
INVx1_ASAP7_75t_L g1293 ( .A(n_472), .Y(n_1293) );
AND2x4_ASAP7_75t_L g478 ( .A(n_473), .B(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_475), .Y(n_700) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_476), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_476), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_476), .A2(n_705), .B1(n_965), .B2(n_966), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_476), .A2(n_1109), .B1(n_1110), .B2(n_1111), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_476), .A2(n_1156), .B1(n_1157), .B2(n_1158), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_476), .A2(n_705), .B1(n_1213), .B2(n_1221), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_476), .A2(n_930), .B1(n_1420), .B2(n_1421), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1792 ( .A1(n_476), .A2(n_930), .B1(n_1769), .B2(n_1793), .Y(n_1792) );
NAND2x1p5_ASAP7_75t_L g717 ( .A(n_477), .B(n_512), .Y(n_717) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g497 ( .A(n_478), .Y(n_497) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_478), .Y(n_556) );
BUFx3_ASAP7_75t_L g566 ( .A(n_478), .Y(n_566) );
BUFx6f_ASAP7_75t_L g861 ( .A(n_478), .Y(n_861) );
INVx1_ASAP7_75t_L g1144 ( .A(n_478), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1280 ( .A(n_478), .B(n_1281), .Y(n_1280) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_481), .B(n_508), .Y(n_480) );
AOI33xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_487), .A3(n_493), .B1(n_498), .B2(n_499), .B3(n_500), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g1315 ( .A(n_484), .Y(n_1315) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
BUFx2_ASAP7_75t_L g608 ( .A(n_485), .Y(n_608) );
OR2x6_ASAP7_75t_L g818 ( .A(n_485), .B(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g844 ( .A(n_485), .Y(n_844) );
AOI31xp33_ASAP7_75t_L g992 ( .A1(n_485), .A2(n_993), .A3(n_1005), .B(n_1017), .Y(n_992) );
AND2x4_ASAP7_75t_L g1127 ( .A(n_485), .B(n_486), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_485), .B(n_864), .Y(n_1151) );
INVx1_ASAP7_75t_L g879 ( .A(n_486), .Y(n_879) );
BUFx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_491), .A2(n_1036), .B1(n_1037), .B2(n_1038), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1433 ( .A1(n_491), .A2(n_1434), .B1(n_1436), .B2(n_1437), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1438 ( .A1(n_491), .A2(n_1439), .B1(n_1440), .B2(n_1441), .Y(n_1438) );
INVx4_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_SL g562 ( .A(n_492), .Y(n_562) );
INVx2_ASAP7_75t_SL g724 ( .A(n_492), .Y(n_724) );
INVx2_ASAP7_75t_SL g858 ( .A(n_492), .Y(n_858) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g519 ( .A(n_497), .B(n_512), .Y(n_519) );
INVx1_ASAP7_75t_L g1279 ( .A(n_497), .Y(n_1279) );
INVx1_ASAP7_75t_L g740 ( .A(n_500), .Y(n_740) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_501), .A2(n_537), .B1(n_540), .B2(n_557), .Y(n_536) );
OAI33xp33_ASAP7_75t_L g939 ( .A1(n_501), .A2(n_537), .A3(n_940), .B1(n_946), .B2(n_952), .B3(n_955), .Y(n_939) );
OAI33xp33_ASAP7_75t_L g1034 ( .A1(n_501), .A2(n_537), .A3(n_1035), .B1(n_1039), .B2(n_1043), .B3(n_1048), .Y(n_1034) );
OAI33xp33_ASAP7_75t_L g1426 ( .A1(n_501), .A2(n_1427), .A3(n_1428), .B1(n_1433), .B2(n_1438), .B3(n_1442), .Y(n_1426) );
CKINVDCx8_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
INVx5_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx6_ASAP7_75t_L g685 ( .A(n_503), .Y(n_685) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g864 ( .A(n_505), .Y(n_864) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g1282 ( .A(n_506), .Y(n_1282) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_513), .B1(n_514), .B2(n_518), .C(n_519), .Y(n_508) );
INVx1_ASAP7_75t_L g613 ( .A(n_509), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_509), .A2(n_514), .B1(n_519), .B2(n_1106), .C(n_1107), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_509), .A2(n_514), .B1(n_519), .B2(n_1138), .C(n_1139), .Y(n_1137) );
AOI221xp5_ASAP7_75t_L g1374 ( .A1(n_509), .A2(n_514), .B1(n_519), .B2(n_1344), .C(n_1345), .Y(n_1374) );
AOI21xp5_ASAP7_75t_L g1410 ( .A1(n_509), .A2(n_519), .B(n_1411), .Y(n_1410) );
AOI221xp5_ASAP7_75t_L g1737 ( .A1(n_509), .A2(n_514), .B1(n_519), .B2(n_1721), .C(n_1722), .Y(n_1737) );
AOI221xp5_ASAP7_75t_L g1781 ( .A1(n_509), .A2(n_514), .B1(n_519), .B2(n_1782), .C(n_1783), .Y(n_1781) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
AND2x2_ASAP7_75t_L g867 ( .A(n_510), .B(n_846), .Y(n_867) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g711 ( .A(n_511), .Y(n_711) );
AND2x4_ASAP7_75t_L g514 ( .A(n_512), .B(n_515), .Y(n_514) );
NAND2x1_ASAP7_75t_SL g709 ( .A(n_512), .B(n_710), .Y(n_709) );
NAND2x1p5_ASAP7_75t_L g714 ( .A(n_512), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g611 ( .A(n_514), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g1397 ( .A1(n_514), .A2(n_533), .B1(n_1382), .B2(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g665 ( .A(n_517), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_517), .B(n_666), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_519), .A2(n_597), .B1(n_598), .B2(n_610), .C(n_612), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_519), .A2(n_610), .B1(n_612), .B2(n_652), .C(n_654), .Y(n_692) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
XOR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_614), .Y(n_521) );
NAND4xp25_ASAP7_75t_L g523 ( .A(n_524), .B(n_534), .C(n_567), .D(n_609), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g585 ( .A1(n_528), .A2(n_535), .B1(n_586), .B2(n_588), .C(n_590), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_531), .B1(n_532), .B2(n_533), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_533), .A2(n_639), .B1(n_690), .B2(n_691), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_533), .A2(n_1160), .B1(n_1161), .B2(n_1162), .Y(n_1159) );
AOI22xp5_ASAP7_75t_L g1367 ( .A1(n_533), .A2(n_1127), .B1(n_1354), .B2(n_1368), .Y(n_1367) );
OAI33xp33_ASAP7_75t_L g657 ( .A1(n_537), .A2(n_658), .A3(n_667), .B1(n_672), .B2(n_677), .B3(n_684), .Y(n_657) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_537), .Y(n_719) );
OAI33xp33_ASAP7_75t_L g1226 ( .A1(n_537), .A2(n_684), .A3(n_1227), .B1(n_1230), .B2(n_1234), .B3(n_1235), .Y(n_1226) );
HB1xp67_ASAP7_75t_L g1427 ( .A(n_537), .Y(n_1427) );
INVx1_ASAP7_75t_L g1289 ( .A(n_539), .Y(n_1289) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_545), .B1(n_546), .B2(n_549), .C(n_550), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g560 ( .A(n_544), .Y(n_560) );
INVx1_ASAP7_75t_L g670 ( .A(n_544), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_545), .A2(n_574), .B1(n_576), .B2(n_577), .C(n_579), .Y(n_573) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_548), .A2(n_622), .B1(n_668), .B2(n_671), .Y(n_667) );
INVx3_ASAP7_75t_L g675 ( .A(n_548), .Y(n_675) );
INVx2_ASAP7_75t_L g1147 ( .A(n_548), .Y(n_1147) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g862 ( .A(n_552), .Y(n_862) );
INVx2_ASAP7_75t_L g1142 ( .A(n_552), .Y(n_1142) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g1317 ( .A(n_553), .Y(n_1317) );
BUFx6f_ASAP7_75t_L g1360 ( .A(n_553), .Y(n_1360) );
AOI22xp5_ASAP7_75t_L g1358 ( .A1(n_554), .A2(n_1359), .B1(n_1360), .B2(n_1361), .Y(n_1358) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g1786 ( .A(n_555), .Y(n_1786) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B1(n_562), .B2(n_563), .C(n_564), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_558), .A2(n_673), .B1(n_674), .B2(n_676), .Y(n_672) );
BUFx2_ASAP7_75t_L g981 ( .A(n_558), .Y(n_981) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g729 ( .A(n_559), .Y(n_729) );
INVx2_ASAP7_75t_L g857 ( .A(n_559), .Y(n_857) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g950 ( .A(n_560), .Y(n_950) );
OAI22xp5_ASAP7_75t_SL g946 ( .A1(n_562), .A2(n_947), .B1(n_948), .B2(n_951), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_562), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_980) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g853 ( .A(n_566), .B(n_854), .Y(n_853) );
OAI31xp33_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_581), .A3(n_591), .B(n_607), .Y(n_567) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_572), .Y(n_1014) );
OAI21xp5_ASAP7_75t_SL g1768 ( .A1(n_574), .A2(n_1769), .B(n_1770), .Y(n_1768) );
INVx2_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g620 ( .A(n_575), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_577), .A2(n_620), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_619) );
INVx1_ASAP7_75t_L g1774 ( .A(n_577), .Y(n_1774) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g771 ( .A(n_580), .Y(n_771) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g605 ( .A(n_584), .Y(n_605) );
BUFx2_ASAP7_75t_L g766 ( .A(n_584), .Y(n_766) );
BUFx3_ASAP7_75t_L g832 ( .A(n_584), .Y(n_832) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_SL g606 ( .A(n_587), .Y(n_606) );
INVx1_ASAP7_75t_L g1168 ( .A(n_587), .Y(n_1168) );
INVx1_ASAP7_75t_L g1725 ( .A(n_587), .Y(n_1725) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_588), .A2(n_606), .B1(n_631), .B2(n_632), .C(n_633), .Y(n_630) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_596), .C(n_599), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_SL g636 ( .A1(n_594), .A2(n_637), .B(n_639), .C(n_640), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g1381 ( .A1(n_594), .A2(n_637), .B(n_1382), .C(n_1383), .Y(n_1381) );
BUFx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g1199 ( .A(n_605), .Y(n_1199) );
OAI21xp33_ASAP7_75t_L g1716 ( .A1(n_606), .A2(n_1717), .B(n_1718), .Y(n_1716) );
CKINVDCx8_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g615 ( .A(n_616), .B(n_656), .C(n_686), .D(n_692), .Y(n_615) );
OAI31xp33_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_625), .A3(n_635), .B(n_655), .Y(n_616) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_618), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_621), .A2(n_659), .B1(n_660), .B2(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g789 ( .A(n_627), .Y(n_789) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g644 ( .A(n_629), .Y(n_644) );
INVx1_ASAP7_75t_L g834 ( .A(n_629), .Y(n_834) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_629), .Y(n_909) );
INVx1_ASAP7_75t_L g760 ( .A(n_633), .Y(n_760) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_642), .C(n_648), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g830 ( .A(n_638), .Y(n_830) );
INVx4_ASAP7_75t_L g905 ( .A(n_638), .Y(n_905) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g915 ( .A(n_641), .Y(n_915) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g1309 ( .A(n_647), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .B1(n_653), .B2(n_654), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx4_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g1101 ( .A(n_651), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_651), .A2(n_653), .B1(n_1138), .B2(n_1139), .Y(n_1182) );
INVx2_ASAP7_75t_L g1462 ( .A(n_651), .Y(n_1462) );
AOI22xp5_ASAP7_75t_L g1720 ( .A1(n_651), .A2(n_653), .B1(n_1721), .B2(n_1722), .Y(n_1720) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_653), .Y(n_1061) );
INVx2_ASAP7_75t_L g1102 ( .A(n_653), .Y(n_1102) );
INVx2_ASAP7_75t_L g1103 ( .A(n_655), .Y(n_1103) );
OAI31xp33_ASAP7_75t_L g1163 ( .A1(n_655), .A2(n_1164), .A3(n_1165), .B(n_1177), .Y(n_1163) );
AOI22xp5_ASAP7_75t_L g1760 ( .A1(n_655), .A2(n_744), .B1(n_1761), .B2(n_1779), .Y(n_1760) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_660), .A2(n_678), .B1(n_679), .B2(n_683), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g1227 ( .A1(n_660), .A2(n_1041), .B1(n_1228), .B2(n_1229), .Y(n_1227) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g722 ( .A(n_661), .Y(n_722) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g890 ( .A(n_664), .B(n_847), .Y(n_890) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_664), .Y(n_986) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g945 ( .A(n_665), .Y(n_945) );
BUFx2_ASAP7_75t_L g957 ( .A(n_665), .Y(n_957) );
INVx3_ASAP7_75t_L g1051 ( .A(n_665), .Y(n_1051) );
BUFx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_670), .Y(n_882) );
INVx2_ASAP7_75t_L g1435 ( .A(n_670), .Y(n_1435) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g1232 ( .A(n_675), .Y(n_1232) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g731 ( .A(n_680), .Y(n_731) );
INVx1_ASAP7_75t_L g1041 ( .A(n_680), .Y(n_1041) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx3_ASAP7_75t_L g738 ( .A(n_681), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_681), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1123) );
BUFx3_ASAP7_75t_L g1237 ( .A(n_681), .Y(n_1237) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g988 ( .A(n_685), .Y(n_988) );
AOI222xp33_ASAP7_75t_L g1115 ( .A1(n_685), .A2(n_1116), .B1(n_1117), .B2(n_1118), .C1(n_1127), .C2(n_1128), .Y(n_1115) );
AOI33xp33_ASAP7_75t_L g1314 ( .A1(n_685), .A2(n_1315), .A3(n_1316), .B1(n_1318), .B2(n_1324), .B3(n_1325), .Y(n_1314) );
AOI322xp5_ASAP7_75t_L g1403 ( .A1(n_685), .A2(n_1127), .A3(n_1390), .B1(n_1404), .B2(n_1405), .C1(n_1406), .C2(n_1409), .Y(n_1403) );
AOI33xp33_ASAP7_75t_L g1784 ( .A1(n_685), .A2(n_1127), .A3(n_1785), .B1(n_1787), .B2(n_1788), .B3(n_1791), .Y(n_1784) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
XNOR2x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_741), .Y(n_697) );
NOR3xp33_ASAP7_75t_SL g698 ( .A(n_699), .B(n_706), .C(n_718), .Y(n_698) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g936 ( .A(n_708), .Y(n_936) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx4f_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx4f_ASAP7_75t_L g937 ( .A(n_714), .Y(n_937) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x6_ASAP7_75t_L g869 ( .A(n_716), .B(n_847), .Y(n_869) );
BUFx3_ASAP7_75t_L g938 ( .A(n_717), .Y(n_938) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_717), .Y(n_1033) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_717), .Y(n_1225) );
OAI33xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .A3(n_725), .B1(n_732), .B2(n_735), .B3(n_740), .Y(n_718) );
OAI33xp33_ASAP7_75t_L g971 ( .A1(n_719), .A2(n_972), .A3(n_975), .B1(n_980), .B2(n_984), .B3(n_988), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_722), .A2(n_736), .B1(n_737), .B2(n_739), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_724), .A2(n_727), .B1(n_733), .B2(n_734), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_730), .B2(n_731), .Y(n_725) );
OAI22xp33_ASAP7_75t_SL g975 ( .A1(n_727), .A2(n_976), .B1(n_978), .B2(n_979), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_727), .A2(n_1231), .B1(n_1232), .B2(n_1233), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_727), .A2(n_1205), .B1(n_1216), .B2(n_1232), .Y(n_1234) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_731), .A2(n_858), .B1(n_973), .B2(n_974), .Y(n_972) );
OAI22xp33_ASAP7_75t_L g1442 ( .A1(n_731), .A2(n_1429), .B1(n_1443), .B2(n_1444), .Y(n_1442) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_733), .A2(n_748), .B(n_749), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g873 ( .A1(n_737), .A2(n_874), .B1(n_875), .B2(n_877), .C(n_878), .Y(n_873) );
BUFx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_739), .A2(n_762), .B1(n_765), .B2(n_772), .C(n_775), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_744), .A2(n_900), .B1(n_901), .B2(n_925), .Y(n_899) );
AOI21xp33_ASAP7_75t_SL g1053 ( .A1(n_744), .A2(n_1054), .B(n_1055), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_744), .A2(n_1191), .B1(n_1193), .B2(n_1217), .Y(n_1190) );
OR2x6_ASAP7_75t_L g815 ( .A(n_752), .B(n_812), .Y(n_815) );
INVx1_ASAP7_75t_L g1009 ( .A(n_754), .Y(n_1009) );
INVx1_ASAP7_75t_L g1059 ( .A(n_754), .Y(n_1059) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx3_ASAP7_75t_L g1307 ( .A(n_770), .Y(n_1307) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g1068 ( .A(n_779), .Y(n_1068) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_1020), .B2(n_1066), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
XNOR2x1_ASAP7_75t_L g781 ( .A(n_782), .B(n_896), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_840), .C(n_850), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_805), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_796), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_792), .B2(n_793), .Y(n_786) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_787), .A2(n_792), .B1(n_857), .B2(n_858), .C(n_859), .Y(n_856) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
AND2x2_ASAP7_75t_L g798 ( .A(n_790), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
OR2x6_ASAP7_75t_L g794 ( .A(n_791), .B(n_795), .Y(n_794) );
OR2x6_ASAP7_75t_L g803 ( .A(n_791), .B(n_804), .Y(n_803) );
CKINVDCx6p67_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B1(n_801), .B2(n_802), .Y(n_796) );
INVx2_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g918 ( .A(n_800), .Y(n_918) );
CKINVDCx6p67_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
BUFx3_ASAP7_75t_L g1173 ( .A(n_804), .Y(n_1173) );
INVx1_ASAP7_75t_L g1392 ( .A(n_804), .Y(n_1392) );
NAND3xp33_ASAP7_75t_SL g805 ( .A(n_806), .B(n_816), .C(n_836), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_813), .B2(n_814), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_807), .A2(n_813), .B1(n_866), .B2(n_868), .Y(n_865) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND2x1p5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx2_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g839 ( .A(n_812), .Y(n_839) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI33xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_820), .A3(n_825), .B1(n_828), .B2(n_831), .B3(n_835), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g1303 ( .A(n_818), .Y(n_1303) );
INVx1_ASAP7_75t_L g1012 ( .A(n_819), .Y(n_1012) );
BUFx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_824), .B(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_824), .Y(n_1264) );
BUFx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g1713 ( .A1(n_834), .A2(n_1339), .B1(n_1714), .B2(n_1715), .Y(n_1713) );
BUFx4f_ASAP7_75t_L g1313 ( .A(n_835), .Y(n_1313) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NOR2xp67_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx2_ASAP7_75t_L g1192 ( .A(n_844), .Y(n_1192) );
AOI211xp5_ASAP7_75t_L g1376 ( .A1(n_844), .A2(n_1377), .B(n_1395), .C(n_1402), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx8_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
AND2x4_ASAP7_75t_L g895 ( .A(n_854), .B(n_887), .Y(n_895) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVxp67_ASAP7_75t_L g1370 ( .A(n_858), .Y(n_1370) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
CKINVDCx11_ASAP7_75t_R g868 ( .A(n_869), .Y(n_868) );
CKINVDCx6p67_ASAP7_75t_R g871 ( .A(n_872), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g1039 ( .A1(n_875), .A2(n_1040), .B1(n_1041), .B2(n_1042), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1236 ( .A(n_875), .Y(n_1236) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_883), .B1(n_884), .B2(n_889), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx3_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
AO22x2_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_959), .B1(n_1018), .B2(n_1019), .Y(n_896) );
INVx1_ASAP7_75t_L g1019 ( .A(n_897), .Y(n_1019) );
XOR2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_958), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_926), .Y(n_898) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_913), .C(n_922), .Y(n_901) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_904), .Y(n_1010) );
INVxp67_ASAP7_75t_L g1210 ( .A(n_908), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_910), .A2(n_924), .B1(n_948), .B2(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1212 ( .A(n_919), .Y(n_1212) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g1310 ( .A(n_920), .Y(n_1310) );
INVx1_ASAP7_75t_L g1352 ( .A(n_920), .Y(n_1352) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_921), .A2(n_923), .B1(n_942), .B2(n_956), .Y(n_955) );
NOR3xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_935), .C(n_939), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_932), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B1(n_944), .B2(n_945), .Y(n_940) );
BUFx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_943), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_984) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_943), .A2(n_1051), .B1(n_1343), .B2(n_1366), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_943), .A2(n_1051), .B1(n_1372), .B2(n_1373), .Y(n_1371) );
INVx1_ASAP7_75t_L g1430 ( .A(n_943), .Y(n_1430) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g1037 ( .A(n_949), .Y(n_1037) );
INVx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
BUFx2_ASAP7_75t_L g1439 ( .A(n_950), .Y(n_1439) );
CKINVDCx5p33_ASAP7_75t_R g953 ( .A(n_954), .Y(n_953) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g1018 ( .A(n_959), .Y(n_1018) );
XNOR2xp5_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_989), .Y(n_961) );
NOR3xp33_ASAP7_75t_SL g962 ( .A(n_963), .B(n_970), .C(n_971), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_967), .Y(n_963) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_976), .A2(n_1049), .B1(n_1050), .B2(n_1052), .Y(n_1048) );
INVx3_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
AOI21xp5_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
AOI31xp33_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_1000), .A3(n_1002), .B(n_1003), .Y(n_995) );
INVx1_ASAP7_75t_L g1097 ( .A(n_997), .Y(n_1097) );
INVx1_ASAP7_75t_L g1340 ( .A(n_998), .Y(n_1340) );
BUFx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1181 ( .A(n_999), .Y(n_1181) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
BUFx2_ASAP7_75t_SL g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1022), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1053), .Y(n_1023) );
NOR3xp33_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1032), .C(n_1034), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1029), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_1037), .A2(n_1044), .B1(n_1045), .B2(n_1047), .Y(n_1043) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1045), .Y(n_1131) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1046), .Y(n_1122) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1046), .Y(n_1364) );
INVx2_ASAP7_75t_L g1790 ( .A(n_1046), .Y(n_1790) );
OAI22xp33_ASAP7_75t_L g1428 ( .A1(n_1050), .A2(n_1429), .B1(n_1431), .B2(n_1432), .Y(n_1428) );
BUFx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
OAI22xp33_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1074), .B1(n_1183), .B2(n_1184), .Y(n_1072) );
INVxp67_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
XNOR2x1_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1134), .Y(n_1076) );
NOR2x1_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1104), .Y(n_1078) );
AOI21xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1092), .B(n_1103), .Y(n_1079) );
AOI221xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1084), .B1(n_1086), .B2(n_1088), .C(n_1091), .Y(n_1080) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1091), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx2_ASAP7_75t_L g1353 ( .A(n_1100), .Y(n_1353) );
NAND4xp25_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1108), .C(n_1112), .D(n_1115), .Y(n_1104) );
AOI22xp5_ASAP7_75t_L g1399 ( .A1(n_1116), .A2(n_1160), .B1(n_1400), .B2(n_1401), .Y(n_1399) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1122), .Y(n_1734) );
AOI33xp33_ASAP7_75t_L g1140 ( .A1(n_1127), .A2(n_1141), .A3(n_1145), .B1(n_1148), .B2(n_1150), .B3(n_1151), .Y(n_1140) );
AOI33xp33_ASAP7_75t_L g1730 ( .A1(n_1127), .A2(n_1151), .A3(n_1731), .B1(n_1733), .B2(n_1735), .B3(n_1736), .Y(n_1730) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1130), .Y(n_1369) );
NAND3xp33_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1154), .C(n_1163), .Y(n_1135) );
AND3x1_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1140), .C(n_1152), .Y(n_1136) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
BUFx3_ASAP7_75t_L g1319 ( .A(n_1149), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1159), .Y(n_1154) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1156), .Y(n_1396) );
OAI211xp5_ASAP7_75t_L g1172 ( .A1(n_1158), .A2(n_1173), .B(n_1174), .C(n_1175), .Y(n_1172) );
INVx2_ASAP7_75t_L g1742 ( .A(n_1160), .Y(n_1742) );
NAND3xp33_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1172), .C(n_1176), .Y(n_1165) );
OAI211xp5_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1168), .B(n_1169), .C(n_1171), .Y(n_1166) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1170), .Y(n_1457) );
OAI211xp5_ASAP7_75t_L g1385 ( .A1(n_1173), .A2(n_1386), .B(n_1387), .C(n_1388), .Y(n_1385) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_1185), .A2(n_1186), .B1(n_1238), .B2(n_1328), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
XNOR2x1_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1189), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1218), .Y(n_1189) );
OAI31xp33_ASAP7_75t_L g1711 ( .A1(n_1191), .A2(n_1712), .A3(n_1719), .B(n_1728), .Y(n_1711) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AOI31xp33_ASAP7_75t_SL g1336 ( .A1(n_1192), .A2(n_1337), .A3(n_1346), .B(n_1349), .Y(n_1336) );
NAND5xp2_ASAP7_75t_SL g1193 ( .A(n_1194), .B(n_1203), .C(n_1206), .D(n_1209), .E(n_1215), .Y(n_1193) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI22xp33_ASAP7_75t_L g1235 ( .A1(n_1197), .A2(n_1204), .B1(n_1236), .B2(n_1237), .Y(n_1235) );
BUFx3_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
OAI221xp5_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1211), .B1(n_1212), .B2(n_1213), .C(n_1214), .Y(n_1209) );
NOR3xp33_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1224), .C(n_1226), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1222), .Y(n_1219) );
INVxp67_ASAP7_75t_SL g1238 ( .A(n_1239), .Y(n_1238) );
HB1xp67_ASAP7_75t_L g1328 ( .A(n_1239), .Y(n_1328) );
INVx2_ASAP7_75t_L g1327 ( .A(n_1240), .Y(n_1327) );
AO211x2_ASAP7_75t_L g1240 ( .A1(n_1241), .A2(n_1243), .B(n_1275), .C(n_1301), .Y(n_1240) );
NAND4xp25_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1255), .C(n_1262), .D(n_1272), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1246), .B1(n_1251), .B2(n_1252), .Y(n_1244) );
HB1xp67_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
AND2x4_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1250), .Y(n_1247) );
INVx1_ASAP7_75t_SL g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1253), .Y(n_1274) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_1256), .A2(n_1257), .B1(n_1260), .B2(n_1261), .Y(n_1255) );
AOI22xp33_ASAP7_75t_SL g1295 ( .A1(n_1256), .A2(n_1296), .B1(n_1297), .B2(n_1298), .Y(n_1295) );
AND2x4_ASAP7_75t_L g1267 ( .A(n_1258), .B(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
AOI222xp33_ASAP7_75t_L g1262 ( .A1(n_1263), .A2(n_1264), .B1(n_1265), .B2(n_1266), .C1(n_1270), .C2(n_1271), .Y(n_1262) );
BUFx4f_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx5_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
AOI31xp33_ASAP7_75t_L g1275 ( .A1(n_1276), .A2(n_1287), .A3(n_1295), .B(n_1300), .Y(n_1275) );
AOI211xp5_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1278), .B(n_1280), .C(n_1283), .Y(n_1276) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
AOI22xp33_ASAP7_75t_SL g1287 ( .A1(n_1288), .A2(n_1290), .B1(n_1291), .B2(n_1294), .Y(n_1287) );
AND2x4_ASAP7_75t_L g1291 ( .A(n_1289), .B(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1323 ( .A(n_1293), .Y(n_1323) );
INVx4_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1314), .Y(n_1301) );
AOI33xp33_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1304), .A3(n_1308), .B1(n_1311), .B2(n_1312), .B3(n_1313), .Y(n_1302) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
XNOR2xp5_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1412), .Y(n_1330) );
HB1xp67_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
XNOR2x1_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1375), .Y(n_1332) );
XNOR2x1_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1335), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1355), .Y(n_1335) );
AOI22xp5_ASAP7_75t_L g1349 ( .A1(n_1350), .A2(n_1351), .B1(n_1353), .B2(n_1354), .Y(n_1349) );
NAND3xp33_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1367), .C(n_1374), .Y(n_1355) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
NAND4xp25_ASAP7_75t_L g1377 ( .A(n_1378), .B(n_1381), .C(n_1385), .D(n_1389), .Y(n_1377) );
OAI211xp5_ASAP7_75t_L g1389 ( .A1(n_1390), .A2(n_1391), .B(n_1393), .C(n_1394), .Y(n_1389) );
INVx2_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1410), .Y(n_1402) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1409), .Y(n_1743) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
HB1xp67_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
XNOR2x1_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1416), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1445), .Y(n_1416) );
NOR3xp33_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1425), .C(n_1426), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1422), .Y(n_1418) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
BUFx2_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
NAND3xp33_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1451), .C(n_1458), .Y(n_1446) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx2_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
OAI221xp5_ASAP7_75t_L g1465 ( .A1(n_1466), .A2(n_1704), .B1(n_1706), .B2(n_1746), .C(n_1752), .Y(n_1465) );
AOI211xp5_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1615), .B(n_1657), .C(n_1683), .Y(n_1466) );
NAND5xp2_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1577), .C(n_1602), .D(n_1607), .E(n_1612), .Y(n_1467) );
AOI21xp5_ASAP7_75t_L g1468 ( .A1(n_1469), .A2(n_1548), .B(n_1556), .Y(n_1468) );
OAI211xp5_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1508), .B(n_1518), .C(n_1542), .Y(n_1469) );
INVxp67_ASAP7_75t_SL g1470 ( .A(n_1471), .Y(n_1470) );
NOR2xp33_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1496), .Y(n_1471) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
AOI22xp5_ASAP7_75t_L g1638 ( .A1(n_1473), .A2(n_1533), .B1(n_1639), .B2(n_1640), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1493), .Y(n_1473) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1474), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_1474), .B(n_1560), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1474), .B(n_1497), .Y(n_1600) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1474), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1474), .B(n_1549), .Y(n_1645) );
AOI221xp5_ASAP7_75t_L g1646 ( .A1(n_1474), .A2(n_1619), .B1(n_1647), .B2(n_1650), .C(n_1654), .Y(n_1646) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1474), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1487), .Y(n_1474) );
AND2x4_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1482), .Y(n_1476) );
OAI21xp33_ASAP7_75t_SL g1798 ( .A1(n_1477), .A2(n_1756), .B(n_1799), .Y(n_1798) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_1478), .B(n_1483), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1481), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1481), .Y(n_1490) );
AND2x4_ASAP7_75t_L g1484 ( .A(n_1482), .B(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1483), .B(n_1486), .Y(n_1507) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
BUFx3_ASAP7_75t_L g1523 ( .A(n_1488), .Y(n_1523) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1488), .Y(n_1553) );
AND2x4_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1491), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1489), .B(n_1491), .Y(n_1514) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
AND2x4_ASAP7_75t_L g1492 ( .A(n_1490), .B(n_1491), .Y(n_1492) );
INVx2_ASAP7_75t_L g1500 ( .A(n_1492), .Y(n_1500) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1493), .Y(n_1541) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1493), .Y(n_1560) );
BUFx6f_ASAP7_75t_L g1598 ( .A(n_1493), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1493), .B(n_1544), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1493), .B(n_1550), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1495), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1496), .B(n_1576), .Y(n_1627) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1496), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1496), .B(n_1587), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1703 ( .A(n_1496), .B(n_1559), .Y(n_1703) );
BUFx3_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
INVx2_ASAP7_75t_SL g1532 ( .A(n_1497), .Y(n_1532) );
NOR2xp33_ASAP7_75t_L g1543 ( .A(n_1497), .B(n_1544), .Y(n_1543) );
BUFx2_ASAP7_75t_L g1584 ( .A(n_1497), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1497), .B(n_1515), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1497), .B(n_1619), .Y(n_1618) );
INVx2_ASAP7_75t_SL g1497 ( .A(n_1498), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1498), .B(n_1564), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1498), .B(n_1544), .Y(n_1697) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1500), .Y(n_1524) );
OAI22xp5_ASAP7_75t_SL g1552 ( .A1(n_1500), .A2(n_1553), .B1(n_1554), .B2(n_1555), .Y(n_1552) );
OAI22xp33_ASAP7_75t_L g1501 ( .A1(n_1502), .A2(n_1503), .B1(n_1505), .B2(n_1506), .Y(n_1501) );
BUFx3_ASAP7_75t_L g1527 ( .A(n_1503), .Y(n_1527) );
BUFx6f_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
HB1xp67_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1507), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1508), .B(n_1579), .Y(n_1578) );
NOR2xp33_ASAP7_75t_L g1654 ( .A(n_1508), .B(n_1655), .Y(n_1654) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
AOI221xp5_ASAP7_75t_L g1617 ( .A1(n_1509), .A2(n_1566), .B1(n_1592), .B2(n_1618), .C(n_1620), .Y(n_1617) );
A2O1A1Ixp33_ASAP7_75t_SL g1634 ( .A1(n_1509), .A2(n_1573), .B(n_1635), .C(n_1636), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1515), .Y(n_1509) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1510), .Y(n_1568) );
OR2x2_ASAP7_75t_L g1641 ( .A(n_1510), .B(n_1515), .Y(n_1641) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1511), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1511), .B(n_1536), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1511), .B(n_1537), .Y(n_1588) );
INVxp67_ASAP7_75t_SL g1594 ( .A(n_1511), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1511), .B(n_1515), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1513), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1515), .B(n_1534), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1515), .B(n_1546), .Y(n_1545) );
CKINVDCx5p33_ASAP7_75t_R g1564 ( .A(n_1515), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1515), .B(n_1593), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1515), .B(n_1588), .Y(n_1614) );
NOR2xp33_ASAP7_75t_L g1625 ( .A(n_1515), .B(n_1535), .Y(n_1625) );
NOR2xp33_ASAP7_75t_L g1632 ( .A(n_1515), .B(n_1568), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1515), .B(n_1571), .Y(n_1643) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1515), .B(n_1535), .Y(n_1674) );
HB1xp67_ASAP7_75t_L g1686 ( .A(n_1515), .Y(n_1686) );
AND2x4_ASAP7_75t_SL g1515 ( .A(n_1516), .B(n_1517), .Y(n_1515) );
OAI21xp5_ASAP7_75t_SL g1518 ( .A1(n_1519), .A2(n_1531), .B(n_1540), .Y(n_1518) );
OAI221xp5_ASAP7_75t_L g1637 ( .A1(n_1519), .A2(n_1550), .B1(n_1638), .B2(n_1642), .C(n_1644), .Y(n_1637) );
INVx2_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1520), .B(n_1541), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1520), .B(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
OAI22xp33_ASAP7_75t_L g1525 ( .A1(n_1526), .A2(n_1527), .B1(n_1528), .B2(n_1529), .Y(n_1525) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1527), .Y(n_1705) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
OAI31xp33_ASAP7_75t_L g1659 ( .A1(n_1531), .A2(n_1603), .A3(n_1660), .B(n_1662), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1533), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1532), .B(n_1571), .Y(n_1570) );
HB1xp67_ASAP7_75t_L g1575 ( .A(n_1532), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1532), .B(n_1625), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1532), .B(n_1559), .Y(n_1656) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1536), .B(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1537), .B(n_1594), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1539), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1541), .B(n_1550), .Y(n_1581) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1541), .Y(n_1596) );
OAI32xp33_ASAP7_75t_L g1620 ( .A1(n_1541), .A2(n_1571), .A3(n_1598), .B1(n_1621), .B2(n_1623), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1666 ( .A(n_1541), .B(n_1550), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1670 ( .A(n_1541), .B(n_1549), .Y(n_1670) );
NAND2xp5_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1545), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1544), .B(n_1560), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1544), .B(n_1549), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1546), .B(n_1564), .Y(n_1576) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1546), .Y(n_1690) );
NAND2xp5_ASAP7_75t_SL g1558 ( .A(n_1549), .B(n_1559), .Y(n_1558) );
AOI32xp33_ASAP7_75t_L g1561 ( .A1(n_1549), .A2(n_1550), .A3(n_1562), .B1(n_1567), .B2(n_1569), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1549), .B(n_1606), .Y(n_1693) );
CKINVDCx6p67_ASAP7_75t_R g1549 ( .A(n_1550), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1611 ( .A(n_1550), .B(n_1566), .Y(n_1611) );
CKINVDCx5p33_ASAP7_75t_R g1616 ( .A(n_1550), .Y(n_1616) );
NAND2xp5_ASAP7_75t_L g1696 ( .A(n_1550), .B(n_1697), .Y(n_1696) );
OR2x6_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1552), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1556 ( .A1(n_1557), .A2(n_1561), .B1(n_1572), .B2(n_1574), .Y(n_1556) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1559), .Y(n_1589) );
AOI211xp5_ASAP7_75t_L g1626 ( .A1(n_1559), .A2(n_1627), .B(n_1628), .C(n_1637), .Y(n_1626) );
INVxp67_ASAP7_75t_SL g1562 ( .A(n_1563), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1564), .B(n_1571), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1564), .B(n_1588), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1564), .B(n_1593), .Y(n_1603) );
OR2x2_ASAP7_75t_L g1653 ( .A(n_1564), .B(n_1570), .Y(n_1653) );
OR2x2_ASAP7_75t_L g1691 ( .A(n_1564), .B(n_1648), .Y(n_1691) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
OAI21xp5_ASAP7_75t_SL g1602 ( .A1(n_1571), .A2(n_1603), .B(n_1604), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1571), .B(n_1595), .Y(n_1672) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
NAND2xp5_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1576), .Y(n_1574) );
AOI311xp33_ASAP7_75t_L g1577 ( .A1(n_1578), .A2(n_1581), .A3(n_1582), .B(n_1585), .C(n_1590), .Y(n_1577) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1581), .B(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1581), .Y(n_1675) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1583), .B(n_1614), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1583), .B(n_1632), .Y(n_1631) );
INVx2_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1584), .B(n_1606), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1636 ( .A(n_1584), .B(n_1588), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1584), .B(n_1596), .Y(n_1639) );
OR2x2_ASAP7_75t_L g1648 ( .A(n_1584), .B(n_1649), .Y(n_1648) );
NAND2xp5_ASAP7_75t_L g1652 ( .A(n_1584), .B(n_1632), .Y(n_1652) );
OR2x2_ASAP7_75t_L g1661 ( .A(n_1584), .B(n_1601), .Y(n_1661) );
NOR2xp33_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1589), .Y(n_1585) );
OAI22xp5_ASAP7_75t_L g1701 ( .A1(n_1586), .A2(n_1598), .B1(n_1702), .B2(n_1703), .Y(n_1701) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
OAI21xp33_ASAP7_75t_L g1630 ( .A1(n_1587), .A2(n_1631), .B(n_1633), .Y(n_1630) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1588), .Y(n_1689) );
OAI21xp33_ASAP7_75t_SL g1590 ( .A1(n_1591), .A2(n_1596), .B(n_1597), .Y(n_1590) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
NAND2xp67_ASAP7_75t_L g1682 ( .A(n_1592), .B(n_1619), .Y(n_1682) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1592), .B(n_1664), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1595), .Y(n_1592) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1593), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1593), .B(n_1622), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1599), .Y(n_1597) );
CKINVDCx14_ASAP7_75t_R g1651 ( .A(n_1598), .Y(n_1651) );
NOR2xp33_ASAP7_75t_SL g1681 ( .A(n_1599), .B(n_1643), .Y(n_1681) );
NOR2xp33_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1601), .Y(n_1599) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1603), .Y(n_1699) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1606), .Y(n_1629) );
INVxp67_ASAP7_75t_SL g1607 ( .A(n_1608), .Y(n_1607) );
NOR2xp33_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1611), .Y(n_1608) );
OAI211xp5_ASAP7_75t_L g1628 ( .A1(n_1609), .A2(n_1629), .B(n_1630), .C(n_1634), .Y(n_1628) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1611), .Y(n_1633) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1614), .Y(n_1700) );
OAI211xp5_ASAP7_75t_L g1615 ( .A1(n_1616), .A2(n_1617), .B(n_1626), .C(n_1646), .Y(n_1615) );
AOI221xp5_ASAP7_75t_L g1667 ( .A1(n_1616), .A2(n_1619), .B1(n_1668), .B2(n_1676), .C(n_1678), .Y(n_1667) );
OAI22xp33_ASAP7_75t_SL g1678 ( .A1(n_1616), .A2(n_1679), .B1(n_1681), .B2(n_1682), .Y(n_1678) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
CKINVDCx5p33_ASAP7_75t_R g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
OAI21xp33_ASAP7_75t_L g1650 ( .A1(n_1651), .A2(n_1652), .B(n_1653), .Y(n_1650) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
O2A1O1Ixp33_ASAP7_75t_L g1694 ( .A1(n_1656), .A2(n_1695), .B(n_1698), .C(n_1701), .Y(n_1694) );
A2O1A1Ixp33_ASAP7_75t_L g1657 ( .A1(n_1658), .A2(n_1659), .B(n_1666), .C(n_1667), .Y(n_1657) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1664), .B(n_1677), .Y(n_1676) );
INVx3_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
OAI22xp5_ASAP7_75t_L g1668 ( .A1(n_1669), .A2(n_1671), .B1(n_1673), .B2(n_1675), .Y(n_1668) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
A2O1A1Ixp33_ASAP7_75t_L g1683 ( .A1(n_1684), .A2(n_1691), .B(n_1692), .C(n_1694), .Y(n_1683) );
INVxp67_ASAP7_75t_SL g1684 ( .A(n_1685), .Y(n_1684) );
NOR2xp33_ASAP7_75t_L g1685 ( .A(n_1686), .B(n_1687), .Y(n_1685) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1690), .Y(n_1688) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVxp67_ASAP7_75t_SL g1695 ( .A(n_1696), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1700), .Y(n_1698) );
CKINVDCx5p33_ASAP7_75t_R g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
HB1xp67_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1709), .Y(n_1745) );
NAND4xp75_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1711), .C(n_1729), .D(n_1738), .Y(n_1709) );
OAI211xp5_ASAP7_75t_L g1723 ( .A1(n_1724), .A2(n_1725), .B(n_1726), .C(n_1727), .Y(n_1723) );
AND2x2_ASAP7_75t_SL g1729 ( .A(n_1730), .B(n_1737), .Y(n_1729) );
INVx1_ASAP7_75t_SL g1746 ( .A(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
CKINVDCx5p33_ASAP7_75t_R g1754 ( .A(n_1755), .Y(n_1754) );
INVxp33_ASAP7_75t_SL g1757 ( .A(n_1758), .Y(n_1757) );
AND2x2_ASAP7_75t_L g1759 ( .A(n_1760), .B(n_1780), .Y(n_1759) );
NAND3xp33_ASAP7_75t_SL g1761 ( .A(n_1762), .B(n_1771), .C(n_1776), .Y(n_1761) );
INVx2_ASAP7_75t_SL g1765 ( .A(n_1766), .Y(n_1765) );
AND4x1_ASAP7_75t_L g1780 ( .A(n_1781), .B(n_1784), .C(n_1792), .D(n_1794), .Y(n_1780) );
INVx2_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
HB1xp67_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
endmodule