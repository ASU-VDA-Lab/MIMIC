module fake_jpeg_6713_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_32),
.B(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_3),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_43),
.Y(n_61)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx12_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_46),
.B1(n_22),
.B2(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_21),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_38),
.C(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_26),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_39),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_72),
.B(n_73),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_25),
.B1(n_40),
.B2(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_25),
.Y(n_85)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_87),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_4),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_66),
.A3(n_75),
.B1(n_70),
.B2(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_42),
.B1(n_47),
.B2(n_54),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_96),
.B1(n_65),
.B2(n_17),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_63),
.A3(n_67),
.B1(n_56),
.B2(n_24),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_56),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_26),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_100),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_23),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_109),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_26),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_117),
.B(n_83),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_116),
.B1(n_82),
.B2(n_87),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_24),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_24),
.B(n_15),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

XOR2x2_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_88),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_117),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_91),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_132),
.C(n_129),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_113),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_133),
.B1(n_110),
.B2(n_97),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_81),
.B1(n_98),
.B2(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_136),
.Y(n_152)
);

NOR2xp67_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_98),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_81),
.B1(n_96),
.B2(n_99),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_112),
.B1(n_111),
.B2(n_113),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_115),
.B1(n_102),
.B2(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_151),
.B1(n_153),
.B2(n_125),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_114),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_126),
.B(n_120),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_105),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_150),
.C(n_132),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_110),
.B(n_104),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_104),
.B1(n_93),
.B2(n_105),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_159),
.C(n_163),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_161),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_145),
.A3(n_149),
.B1(n_138),
.B2(n_139),
.C(n_147),
.Y(n_169)
);

AOI211xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_126),
.B(n_130),
.C(n_128),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_158),
.B(n_142),
.C(n_77),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_80),
.C(n_125),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_20),
.B1(n_23),
.B2(n_17),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_136),
.C(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_108),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_172),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_163),
.B(n_118),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_153),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_176),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_175),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_77),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_53),
.C(n_50),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_65),
.B1(n_20),
.B2(n_50),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_160),
.C(n_158),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_184),
.B(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_157),
.B1(n_165),
.B2(n_14),
.Y(n_182)
);

OAI21x1_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_6),
.B(n_7),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_186),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_65),
.B1(n_53),
.B2(n_50),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_171),
.A3(n_167),
.B1(n_14),
.B2(n_19),
.C1(n_15),
.C2(n_11),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_190),
.B(n_193),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_192),
.B(n_8),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_179),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_15),
.B(n_19),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_182),
.B(n_6),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_19),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_181),
.B1(n_10),
.B2(n_11),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_19),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.C(n_202),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_9),
.C(n_10),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_9),
.C(n_12),
.Y(n_204)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_12),
.B1(n_13),
.B2(n_19),
.C(n_203),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_12),
.Y(n_206)
);


endmodule