module fake_netlist_1_12387_n_1006 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1006);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1006;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_667;
wire n_496;
wire n_311;
wire n_988;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_505;
wire n_823;
wire n_822;
wire n_970;
wire n_706;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_875;
wire n_339;
wire n_657;
wire n_583;
wire n_728;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_84), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_266), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_104), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_138), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_246), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_275), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_241), .Y(n_295) );
XOR2x2_ASAP7_75t_L g296 ( .A(n_37), .B(n_10), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_117), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_0), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_51), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_189), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_66), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_2), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_68), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_90), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_201), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_121), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_248), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_235), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_204), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_252), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_264), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_93), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_162), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_98), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_236), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_85), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_4), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_247), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_265), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_129), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_118), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_176), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_31), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_263), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_4), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_178), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_77), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_135), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_258), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_231), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g333 ( .A(n_260), .B(n_242), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_127), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_159), .Y(n_335) );
NOR2xp67_ASAP7_75t_L g336 ( .A(n_243), .B(n_177), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_268), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_140), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_11), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_78), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_226), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_249), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_259), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_46), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_202), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_57), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_134), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_1), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_33), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_7), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_16), .Y(n_351) );
NOR2xp67_ASAP7_75t_L g352 ( .A(n_44), .B(n_28), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_13), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_167), .Y(n_354) );
BUFx10_ASAP7_75t_L g355 ( .A(n_19), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_12), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_244), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_279), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_262), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_184), .Y(n_360) );
CKINVDCx14_ASAP7_75t_R g361 ( .A(n_211), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_30), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_154), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_130), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_111), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_180), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_116), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_120), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_141), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_163), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_232), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_239), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_192), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_59), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_257), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_224), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_112), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_196), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_255), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_277), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_250), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_221), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_72), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_71), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_24), .Y(n_385) );
BUFx10_ASAP7_75t_L g386 ( .A(n_70), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_213), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_283), .B(n_151), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_254), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_181), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_101), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_170), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_26), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_62), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_55), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_234), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_233), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_76), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_198), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_270), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_110), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_91), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_146), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_36), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_245), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_61), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_237), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_97), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_256), .Y(n_409) );
BUFx8_ASAP7_75t_SL g410 ( .A(n_238), .Y(n_410) );
XNOR2xp5_ASAP7_75t_L g411 ( .A(n_253), .B(n_267), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_190), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_153), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_240), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_175), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_230), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_188), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_22), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_19), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_79), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_169), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_50), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_408), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_310), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_355), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_341), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_310), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_350), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_355), .Y(n_429) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_391), .B(n_21), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_315), .B(n_3), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_380), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_293), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_327), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_294), .Y(n_435) );
NOR2xp33_ASAP7_75t_SL g436 ( .A(n_288), .B(n_23), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_307), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_298), .A2(n_6), .B1(n_3), .B2(n_5), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_353), .Y(n_439) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_291), .A2(n_27), .B(n_25), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_302), .B(n_5), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_318), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_356), .B(n_6), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_289), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_386), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_433), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_424), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_433), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_432), .B(n_373), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_434), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_427), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_431), .Y(n_453) );
INVx2_ASAP7_75t_SL g454 ( .A(n_434), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_446), .B(n_386), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_435), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_446), .B(n_300), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_431), .Y(n_458) );
AOI21x1_ASAP7_75t_L g459 ( .A1(n_440), .A2(n_304), .B(n_292), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_437), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_439), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_442), .B(n_395), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_444), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_445), .B(n_306), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_445), .B(n_312), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_429), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_453), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_458), .B(n_423), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_463), .A2(n_443), .B1(n_441), .B2(n_426), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_448), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_464), .B(n_429), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_466), .B(n_425), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_464), .B(n_430), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_466), .B(n_436), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_452), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_454), .B(n_436), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_455), .B(n_438), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_451), .B(n_443), .Y(n_478) );
O2A1O1Ixp5_ASAP7_75t_L g479 ( .A1(n_459), .A2(n_316), .B(n_319), .C(n_313), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_465), .B(n_290), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_462), .A2(n_323), .B(n_324), .C(n_321), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_457), .B(n_379), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_456), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_449), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_465), .B(n_361), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_461), .A2(n_428), .B1(n_347), .B2(n_362), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_460), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_447), .B(n_297), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_450), .B(n_384), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_450), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_453), .B(n_299), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_491), .A2(n_440), .B(n_330), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_467), .B(n_301), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_468), .A2(n_334), .B(n_326), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_490), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_485), .A2(n_344), .B(n_340), .Y(n_496) );
INVx4_ASAP7_75t_L g497 ( .A(n_484), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_478), .B(n_296), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_469), .B(n_339), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_471), .A2(n_366), .B(n_359), .Y(n_500) );
AO32x1_ASAP7_75t_L g501 ( .A1(n_486), .A2(n_428), .A3(n_369), .B1(n_370), .B2(n_368), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_484), .Y(n_502) );
OAI21xp33_ASAP7_75t_L g503 ( .A1(n_472), .A2(n_351), .B(n_348), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_473), .A2(n_374), .B(n_367), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_489), .B(n_332), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_486), .A2(n_394), .B1(n_403), .B2(n_385), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_479), .A2(n_381), .B(n_377), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_470), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_481), .A2(n_390), .B(n_397), .C(n_383), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g510 ( .A(n_477), .B(n_411), .Y(n_510) );
AOI22x1_ASAP7_75t_SL g511 ( .A1(n_475), .A2(n_305), .B1(n_308), .B2(n_303), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_474), .A2(n_405), .B(n_402), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_483), .A2(n_415), .B(n_409), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_487), .Y(n_514) );
OR2x6_ASAP7_75t_L g515 ( .A(n_477), .B(n_333), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_476), .A2(n_418), .B(n_422), .C(n_420), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_482), .B(n_410), .Y(n_517) );
AOI21x1_ASAP7_75t_L g518 ( .A1(n_492), .A2(n_352), .B(n_336), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_496), .A2(n_480), .B(n_488), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g520 ( .A(n_498), .B(n_7), .Y(n_520) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_507), .A2(n_388), .B(n_314), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_510), .B(n_8), .Y(n_522) );
BUFx4_ASAP7_75t_SL g523 ( .A(n_515), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_508), .B(n_309), .Y(n_524) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_512), .A2(n_314), .B(n_295), .Y(n_525) );
BUFx6f_ASAP7_75t_SL g526 ( .A(n_515), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_500), .A2(n_416), .B(n_317), .Y(n_527) );
AO32x2_ASAP7_75t_L g528 ( .A1(n_497), .A2(n_501), .A3(n_509), .B1(n_513), .B2(n_516), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_504), .A2(n_376), .B(n_393), .C(n_346), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_514), .A2(n_320), .B(n_311), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_499), .B(n_322), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_511), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_501), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_495), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_494), .A2(n_328), .B(n_325), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_505), .B(n_329), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_502), .B(n_295), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_503), .B(n_331), .Y(n_538) );
BUFx10_ASAP7_75t_L g539 ( .A(n_517), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_493), .B(n_335), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_505), .A2(n_338), .B1(n_342), .B2(n_337), .Y(n_541) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_492), .A2(n_314), .B(n_295), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_508), .B(n_8), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_505), .A2(n_345), .B1(n_349), .B2(n_343), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_492), .A2(n_357), .B(n_354), .Y(n_545) );
O2A1O1Ixp5_ASAP7_75t_L g546 ( .A1(n_492), .A2(n_360), .B(n_363), .C(n_358), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_492), .A2(n_365), .B(n_364), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_498), .B(n_9), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_506), .B(n_421), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_498), .B(n_9), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_522), .B(n_10), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_548), .A2(n_412), .B1(n_389), .B2(n_372), .Y(n_552) );
BUFx3_ASAP7_75t_L g553 ( .A(n_532), .Y(n_553) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_542), .A2(n_412), .B(n_389), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_537), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_546), .A2(n_375), .B(n_371), .Y(n_556) );
AOI22x1_ASAP7_75t_L g557 ( .A1(n_545), .A2(n_412), .B1(n_389), .B2(n_382), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_533), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_539), .Y(n_559) );
AOI221x1_ASAP7_75t_L g560 ( .A1(n_547), .A2(n_11), .B1(n_12), .B2(n_13), .C(n_14), .Y(n_560) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_521), .A2(n_387), .B(n_378), .Y(n_561) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_525), .A2(n_32), .B(n_29), .Y(n_562) );
AOI21x1_ASAP7_75t_L g563 ( .A1(n_518), .A2(n_417), .B(n_396), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_543), .A2(n_398), .B1(n_399), .B2(n_392), .Y(n_564) );
O2A1O1Ixp33_ASAP7_75t_SL g565 ( .A1(n_529), .A2(n_35), .B(n_38), .C(n_34), .Y(n_565) );
BUFx2_ASAP7_75t_L g566 ( .A(n_543), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_534), .Y(n_567) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_519), .A2(n_40), .B(n_39), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_550), .A2(n_401), .B1(n_404), .B2(n_400), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_549), .A2(n_16), .B(n_14), .C(n_15), .Y(n_570) );
AND2x2_ASAP7_75t_SL g571 ( .A(n_523), .B(n_15), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_524), .B(n_17), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_526), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_528), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_528), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_527), .A2(n_42), .B(n_41), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_526), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_536), .A2(n_407), .B1(n_413), .B2(n_406), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_531), .A2(n_414), .B(n_45), .Y(n_580) );
BUFx3_ASAP7_75t_L g581 ( .A(n_539), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_528), .Y(n_582) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_530), .A2(n_47), .B(n_43), .Y(n_583) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_538), .A2(n_49), .B(n_48), .Y(n_584) );
BUFx3_ASAP7_75t_L g585 ( .A(n_541), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_540), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_535), .A2(n_18), .B(n_20), .C(n_52), .Y(n_587) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_544), .A2(n_54), .B(n_53), .Y(n_588) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_542), .A2(n_58), .B(n_56), .Y(n_589) );
OR2x6_ASAP7_75t_L g590 ( .A(n_543), .B(n_20), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_548), .B(n_60), .Y(n_591) );
OR2x6_ASAP7_75t_L g592 ( .A(n_543), .B(n_63), .Y(n_592) );
INVx4_ASAP7_75t_SL g593 ( .A(n_526), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_549), .B(n_64), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_543), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_533), .Y(n_596) );
CKINVDCx16_ASAP7_75t_R g597 ( .A(n_526), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_543), .Y(n_598) );
AO21x2_ASAP7_75t_L g599 ( .A1(n_542), .A2(n_65), .B(n_67), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_558), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_596), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_590), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_582), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_590), .B(n_69), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_566), .B(n_73), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_581), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_574), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_567), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_570), .A2(n_74), .B(n_75), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_595), .B(n_287), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_598), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_598), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_592), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_572), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_559), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_553), .Y(n_617) );
BUFx3_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
OAI22xp33_ASAP7_75t_SL g619 ( .A1(n_592), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_555), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_551), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_555), .B(n_83), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_600), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_571), .B(n_86), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_551), .Y(n_625) );
BUFx4f_ASAP7_75t_SL g626 ( .A(n_593), .Y(n_626) );
OR2x6_ASAP7_75t_L g627 ( .A(n_600), .B(n_87), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_585), .B(n_88), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_568), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_564), .B(n_89), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_578), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_597), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_576), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_574), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
OA21x2_ASAP7_75t_L g636 ( .A1(n_575), .A2(n_92), .B(n_94), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_562), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_586), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_561), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_593), .Y(n_640) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_554), .A2(n_589), .B(n_560), .Y(n_641) );
AO21x2_ASAP7_75t_L g642 ( .A1(n_599), .A2(n_95), .B(n_96), .Y(n_642) );
OAI21x1_ASAP7_75t_L g643 ( .A1(n_577), .A2(n_99), .B(n_100), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_569), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_561), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_583), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_588), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_552), .B(n_285), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_591), .B(n_102), .Y(n_649) );
AOI21x1_ASAP7_75t_L g650 ( .A1(n_563), .A2(n_284), .B(n_103), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_560), .B(n_105), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_587), .Y(n_652) );
BUFx12f_ASAP7_75t_L g653 ( .A(n_594), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_584), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_556), .B(n_106), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_565), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_557), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_580), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_579), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_567), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_597), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_567), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_590), .B(n_282), .Y(n_663) );
BUFx5_ASAP7_75t_L g664 ( .A(n_598), .Y(n_664) );
OAI21x1_ASAP7_75t_L g665 ( .A1(n_554), .A2(n_107), .B(n_108), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_590), .A2(n_109), .B1(n_113), .B2(n_114), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_558), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_558), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_558), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_558), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_558), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_558), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_558), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_590), .B(n_115), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_558), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_558), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_555), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_601), .Y(n_678) );
INVx3_ASAP7_75t_SL g679 ( .A(n_632), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_609), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_660), .B(n_119), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_662), .B(n_122), .Y(n_682) );
AO21x2_ASAP7_75t_L g683 ( .A1(n_639), .A2(n_645), .B(n_657), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_614), .B(n_123), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_612), .B(n_124), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_615), .B(n_125), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_607), .B(n_126), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_620), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_624), .B(n_128), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_638), .B(n_131), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_670), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_605), .B(n_132), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_603), .B(n_281), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_621), .B(n_133), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_613), .B(n_280), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_625), .Y(n_696) );
INVx2_ASAP7_75t_SL g697 ( .A(n_626), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_601), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_674), .B(n_136), .Y(n_699) );
AND2x4_ASAP7_75t_L g700 ( .A(n_602), .B(n_137), .Y(n_700) );
BUFx2_ASAP7_75t_SL g701 ( .A(n_617), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_633), .B(n_278), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_627), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_627), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_667), .B(n_276), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_623), .B(n_139), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_667), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_668), .B(n_274), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_623), .B(n_142), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_677), .B(n_143), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_669), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_677), .B(n_144), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_671), .Y(n_713) );
INVxp67_ASAP7_75t_R g714 ( .A(n_606), .Y(n_714) );
INVx3_ASAP7_75t_L g715 ( .A(n_622), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_663), .B(n_145), .Y(n_716) );
INVx4_ASAP7_75t_L g717 ( .A(n_622), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_628), .B(n_147), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_672), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_672), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_673), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_673), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_659), .B(n_148), .Y(n_723) );
INVx3_ASAP7_75t_L g724 ( .A(n_655), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_644), .B(n_149), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_675), .Y(n_726) );
INVx4_ASAP7_75t_L g727 ( .A(n_616), .Y(n_727) );
OR2x2_ASAP7_75t_SL g728 ( .A(n_636), .B(n_150), .Y(n_728) );
BUFx3_ASAP7_75t_L g729 ( .A(n_618), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_676), .Y(n_730) );
INVx3_ASAP7_75t_L g731 ( .A(n_655), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_676), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_630), .B(n_152), .Y(n_733) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_664), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_640), .B(n_155), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_653), .B(n_156), .Y(n_736) );
INVx4_ASAP7_75t_SL g737 ( .A(n_631), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_604), .Y(n_738) );
AND2x4_ASAP7_75t_L g739 ( .A(n_608), .B(n_157), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_604), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_664), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_634), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_661), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_635), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_608), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_664), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_619), .Y(n_747) );
AND2x4_ASAP7_75t_L g748 ( .A(n_647), .B(n_158), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_652), .B(n_160), .Y(n_749) );
OR2x2_ASAP7_75t_L g750 ( .A(n_664), .B(n_273), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_611), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_647), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_651), .B(n_161), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_636), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_651), .B(n_272), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_649), .B(n_164), .Y(n_756) );
INVxp67_ASAP7_75t_SL g757 ( .A(n_637), .Y(n_757) );
INVx1_ASAP7_75t_SL g758 ( .A(n_648), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_650), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_637), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_666), .B(n_165), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_637), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_646), .Y(n_763) );
BUFx3_ASAP7_75t_L g764 ( .A(n_658), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_629), .Y(n_765) );
BUFx3_ASAP7_75t_L g766 ( .A(n_665), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_654), .B(n_271), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_641), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_643), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_641), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_642), .Y(n_771) );
OR2x2_ASAP7_75t_L g772 ( .A(n_720), .B(n_610), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_717), .B(n_656), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_680), .B(n_166), .Y(n_774) );
INVx3_ASAP7_75t_L g775 ( .A(n_717), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_722), .B(n_168), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_698), .B(n_171), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_738), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_688), .B(n_172), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_713), .B(n_173), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_707), .Y(n_781) );
AND2x4_ASAP7_75t_SL g782 ( .A(n_727), .B(n_174), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_738), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_703), .Y(n_784) );
BUFx2_ASAP7_75t_L g785 ( .A(n_704), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_719), .B(n_179), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_711), .Y(n_787) );
NAND4xp25_ASAP7_75t_L g788 ( .A(n_725), .B(n_269), .C(n_183), .D(n_185), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_678), .B(n_182), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_691), .B(n_186), .Y(n_790) );
INVx2_ASAP7_75t_SL g791 ( .A(n_729), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_741), .B(n_187), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_726), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_740), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_732), .B(n_191), .Y(n_795) );
INVxp67_ASAP7_75t_L g796 ( .A(n_701), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_740), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_714), .B(n_193), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_678), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_721), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_721), .B(n_194), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_730), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_745), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_741), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_724), .B(n_195), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_730), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_696), .B(n_197), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_747), .A2(n_199), .B1(n_200), .B2(n_203), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_715), .B(n_205), .Y(n_809) );
INVx3_ASAP7_75t_L g810 ( .A(n_715), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_742), .B(n_206), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_744), .B(n_207), .Y(n_812) );
BUFx2_ASAP7_75t_L g813 ( .A(n_737), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_763), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_686), .B(n_208), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_687), .B(n_209), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_764), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_763), .Y(n_818) );
AND2x4_ASAP7_75t_L g819 ( .A(n_724), .B(n_210), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_727), .B(n_212), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_765), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_734), .Y(n_822) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_731), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_731), .B(n_214), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_751), .B(n_215), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_765), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_739), .B(n_216), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_739), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_758), .B(n_217), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_752), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_700), .Y(n_831) );
OR2x2_ASAP7_75t_L g832 ( .A(n_708), .B(n_218), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_700), .Y(n_833) );
BUFx2_ASAP7_75t_L g834 ( .A(n_737), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_684), .B(n_219), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_692), .B(n_699), .Y(n_836) );
CKINVDCx16_ASAP7_75t_R g837 ( .A(n_697), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_702), .B(n_220), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_768), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_768), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_750), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_681), .B(n_222), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_752), .Y(n_843) );
OR2x2_ASAP7_75t_L g844 ( .A(n_693), .B(n_223), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_770), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_770), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_682), .B(n_225), .Y(n_847) );
INVx2_ASAP7_75t_SL g848 ( .A(n_679), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_784), .B(n_746), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_817), .B(n_757), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_800), .Y(n_851) );
INVxp33_ASAP7_75t_L g852 ( .A(n_813), .Y(n_852) );
AND2x4_ASAP7_75t_L g853 ( .A(n_823), .B(n_760), .Y(n_853) );
BUFx2_ASAP7_75t_L g854 ( .A(n_834), .Y(n_854) );
INVx1_ASAP7_75t_SL g855 ( .A(n_785), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_781), .Y(n_856) );
INVx2_ASAP7_75t_SL g857 ( .A(n_837), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_787), .B(n_760), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_796), .B(n_743), .Y(n_859) );
NOR2xp67_ASAP7_75t_L g860 ( .A(n_775), .B(n_759), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_778), .Y(n_861) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_822), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_778), .Y(n_863) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_793), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_783), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_783), .B(n_723), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_803), .B(n_762), .Y(n_867) );
INVxp67_ASAP7_75t_L g868 ( .A(n_791), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_794), .B(n_771), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_803), .B(n_762), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_794), .B(n_771), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_810), .B(n_736), .Y(n_872) );
OR2x2_ASAP7_75t_L g873 ( .A(n_799), .B(n_767), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_797), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_797), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_802), .B(n_683), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_848), .B(n_837), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_806), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_830), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_810), .B(n_748), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_836), .B(n_748), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_839), .Y(n_882) );
AND2x4_ASAP7_75t_L g883 ( .A(n_804), .B(n_766), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_845), .B(n_754), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_840), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_845), .B(n_754), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_775), .B(n_689), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_841), .B(n_716), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_828), .B(n_685), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_814), .B(n_685), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_831), .B(n_690), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_814), .B(n_753), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_818), .B(n_755), .Y(n_893) );
NOR2x1_ASAP7_75t_L g894 ( .A(n_820), .B(n_695), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_846), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_846), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_833), .B(n_735), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_818), .B(n_769), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_804), .B(n_718), .Y(n_899) );
NAND2x1p5_ASAP7_75t_L g900 ( .A(n_857), .B(n_798), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_864), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_862), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_851), .Y(n_903) );
NAND3xp33_ASAP7_75t_SL g904 ( .A(n_854), .B(n_808), .C(n_827), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_855), .B(n_881), .Y(n_905) );
NOR2x1_ASAP7_75t_L g906 ( .A(n_877), .B(n_788), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_879), .Y(n_907) );
BUFx2_ASAP7_75t_L g908 ( .A(n_868), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_855), .B(n_830), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_861), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_863), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_865), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_874), .B(n_843), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_875), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_878), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_884), .Y(n_916) );
INVx6_ASAP7_75t_L g917 ( .A(n_850), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_895), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_896), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_849), .B(n_843), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_856), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_884), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_888), .B(n_773), .Y(n_923) );
NOR2xp67_ASAP7_75t_R g924 ( .A(n_852), .B(n_782), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_899), .B(n_773), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_886), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_866), .B(n_772), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_883), .B(n_821), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_886), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_867), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_870), .Y(n_931) );
AOI32xp33_ASAP7_75t_L g932 ( .A1(n_906), .A2(n_894), .A3(n_859), .B1(n_887), .B2(n_872), .Y(n_932) );
NOR2x1_ASAP7_75t_L g933 ( .A(n_908), .B(n_860), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_917), .Y(n_934) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_900), .A2(n_890), .B1(n_825), .B2(n_893), .C(n_892), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_927), .B(n_882), .Y(n_936) );
NAND3xp33_ASAP7_75t_L g937 ( .A(n_901), .B(n_869), .C(n_871), .Y(n_937) );
INVxp67_ASAP7_75t_L g938 ( .A(n_902), .Y(n_938) );
OAI21xp5_ASAP7_75t_L g939 ( .A1(n_904), .A2(n_860), .B(n_779), .Y(n_939) );
NAND2x1p5_ASAP7_75t_L g940 ( .A(n_924), .B(n_805), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_917), .A2(n_897), .B1(n_889), .B2(n_891), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_905), .B(n_880), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_923), .B(n_853), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_909), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_916), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_925), .A2(n_728), .B1(n_853), .B2(n_819), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_930), .B(n_885), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_931), .B(n_916), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_920), .B(n_883), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_922), .B(n_858), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_921), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_951), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_948), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_945), .B(n_926), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_936), .Y(n_955) );
NOR2x1p5_ASAP7_75t_L g956 ( .A(n_934), .B(n_903), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_946), .A2(n_928), .B1(n_929), .B2(n_915), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_938), .B(n_928), .Y(n_958) );
AOI21xp5_ASAP7_75t_SL g959 ( .A1(n_940), .A2(n_805), .B(n_819), .Y(n_959) );
INVx1_ASAP7_75t_SL g960 ( .A(n_943), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_945), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_947), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_935), .B(n_907), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_933), .A2(n_914), .B1(n_912), .B2(n_911), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_950), .Y(n_965) );
O2A1O1Ixp33_ASAP7_75t_SL g966 ( .A1(n_964), .A2(n_939), .B(n_932), .C(n_937), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_959), .A2(n_949), .B(n_913), .Y(n_967) );
A2O1A1O1Ixp25_ASAP7_75t_L g968 ( .A1(n_964), .A2(n_910), .B(n_919), .C(n_918), .D(n_941), .Y(n_968) );
NAND3xp33_ASAP7_75t_SL g969 ( .A(n_957), .B(n_844), .C(n_838), .Y(n_969) );
O2A1O1Ixp33_ASAP7_75t_L g970 ( .A1(n_963), .A2(n_829), .B(n_835), .C(n_824), .Y(n_970) );
AOI211xp5_ASAP7_75t_L g971 ( .A1(n_958), .A2(n_942), .B(n_816), .C(n_733), .Y(n_971) );
AOI211xp5_ASAP7_75t_L g972 ( .A1(n_960), .A2(n_944), .B(n_807), .C(n_774), .Y(n_972) );
AOI21xp33_ASAP7_75t_L g973 ( .A1(n_965), .A2(n_869), .B(n_871), .Y(n_973) );
NAND3xp33_ASAP7_75t_SL g974 ( .A(n_953), .B(n_832), .C(n_776), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_973), .B(n_955), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_971), .B(n_962), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_966), .B(n_954), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_969), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_974), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_970), .B(n_961), .Y(n_980) );
NOR3xp33_ASAP7_75t_L g981 ( .A(n_977), .B(n_968), .C(n_967), .Y(n_981) );
AND3x4_ASAP7_75t_L g982 ( .A(n_978), .B(n_952), .C(n_972), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_979), .B(n_956), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_980), .B(n_873), .Y(n_984) );
NAND4xp75_ASAP7_75t_L g985 ( .A(n_976), .B(n_761), .C(n_809), .D(n_847), .Y(n_985) );
NOR2xp67_ASAP7_75t_L g986 ( .A(n_983), .B(n_975), .Y(n_986) );
NOR3xp33_ASAP7_75t_L g987 ( .A(n_981), .B(n_756), .C(n_694), .Y(n_987) );
NOR2x1_ASAP7_75t_L g988 ( .A(n_982), .B(n_792), .Y(n_988) );
NOR2x1_ASAP7_75t_L g989 ( .A(n_985), .B(n_792), .Y(n_989) );
XOR2xp5_ASAP7_75t_L g990 ( .A(n_988), .B(n_984), .Y(n_990) );
AND2x4_ASAP7_75t_L g991 ( .A(n_986), .B(n_876), .Y(n_991) );
NAND4xp75_ASAP7_75t_L g992 ( .A(n_989), .B(n_842), .C(n_815), .D(n_706), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_991), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_990), .A2(n_987), .B1(n_709), .B2(n_710), .Y(n_994) );
A2O1A1Ixp33_ASAP7_75t_L g995 ( .A1(n_992), .A2(n_712), .B(n_780), .C(n_786), .Y(n_995) );
NAND3x1_ASAP7_75t_L g996 ( .A(n_994), .B(n_777), .C(n_749), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_993), .B(n_995), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_997), .B(n_876), .Y(n_998) );
NOR2xp67_ASAP7_75t_L g999 ( .A(n_996), .B(n_227), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_998), .B(n_898), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_999), .B(n_898), .Y(n_1001) );
OAI221xp5_ASAP7_75t_L g1002 ( .A1(n_1001), .A2(n_789), .B1(n_801), .B2(n_705), .C(n_795), .Y(n_1002) );
AOI21xp33_ASAP7_75t_L g1003 ( .A1(n_1000), .A2(n_228), .B(n_229), .Y(n_1003) );
AOI21xp5_ASAP7_75t_L g1004 ( .A1(n_1003), .A2(n_811), .B(n_812), .Y(n_1004) );
OR2x6_ASAP7_75t_L g1005 ( .A(n_1004), .B(n_1002), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_1005), .A2(n_821), .B1(n_826), .B2(n_790), .Y(n_1006) );
endmodule