module real_jpeg_1777_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_38),
.B1(n_49),
.B2(n_55),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_31),
.B1(n_33),
.B2(n_62),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_5),
.A2(n_49),
.B1(n_55),
.B2(n_62),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_8),
.A2(n_35),
.B1(n_85),
.B2(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_8),
.A2(n_35),
.B1(n_49),
.B2(n_55),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_11),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_11),
.B(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_87),
.B(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_11),
.B(n_24),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_33),
.B(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_11),
.B(n_49),
.C(n_65),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_11),
.B(n_52),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_11),
.B(n_70),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_12),
.A2(n_49),
.B1(n_55),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_12),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_14),
.A2(n_49),
.B1(n_55),
.B2(n_69),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_111),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_110),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_81),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_20),
.B(n_81),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_59),
.C(n_71),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_21),
.B(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_40),
.C(n_58),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_23),
.A2(n_36),
.B1(n_37),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_125),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

AO22x2_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_25),
.A2(n_26),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_25),
.B(n_29),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_26),
.A2(n_28),
.A3(n_33),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_26),
.B(n_135),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_28),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_31),
.B(n_74),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_31),
.B(n_45),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_33),
.A2(n_44),
.A3(n_85),
.B1(n_87),
.B2(n_89),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_47),
.B2(n_58),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_43),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_45),
.B1(n_85),
.B2(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_48),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_52),
.B1(n_56),
.B2(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_48),
.A2(n_52),
.B1(n_79),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_48),
.A2(n_52),
.B1(n_74),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_48),
.A2(n_52),
.B1(n_147),
.B2(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_49),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_49),
.B(n_145),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_51),
.A2(n_77),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_59),
.B(n_71),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_70),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_61),
.A2(n_67),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_68),
.B1(n_70),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_70),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_63),
.A2(n_70),
.B1(n_116),
.B2(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_95),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_94),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_161),
.B(n_165),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_130),
.B(n_160),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_121),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_118),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_124),
.C(n_127),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_141),
.B(n_159),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_153),
.B(n_158),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_148),
.B(n_152),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_150),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_164),
.Y(n_165)
);


endmodule