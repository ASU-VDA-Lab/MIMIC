module fake_jpeg_21534_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_23),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_20),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_19),
.B1(n_32),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_54),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_19),
.B1(n_31),
.B2(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_17),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_40),
.C(n_33),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_26),
.B1(n_22),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_30),
.B1(n_39),
.B2(n_33),
.Y(n_72)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_62),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_21),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_81),
.C(n_49),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_42),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_70),
.B(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_73),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_16),
.B(n_21),
.C(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_58),
.B1(n_52),
.B2(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_77),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_40),
.B(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_56),
.B1(n_57),
.B2(n_43),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_48),
.B1(n_45),
.B2(n_51),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_95),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_43),
.B1(n_52),
.B2(n_58),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_43),
.B1(n_52),
.B2(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_80),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_63),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_67),
.B1(n_58),
.B2(n_52),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_81),
.C(n_68),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_119),
.C(n_130),
.Y(n_134)
);

AO21x2_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_64),
.B(n_70),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_114),
.B(n_105),
.C(n_4),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_68),
.B(n_72),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_120),
.B(n_126),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_123),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_83),
.A3(n_76),
.B1(n_78),
.B2(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_80),
.B(n_22),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_27),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_27),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_88),
.B(n_96),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_55),
.C(n_59),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_71),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_132),
.B(n_105),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_93),
.A3(n_94),
.B1(n_107),
.B2(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_92),
.B1(n_102),
.B2(n_95),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_123),
.B1(n_127),
.B2(n_111),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_119),
.C(n_126),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_118),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_100),
.B1(n_87),
.B2(n_98),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_146),
.B1(n_152),
.B2(n_154),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_131),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_98),
.B1(n_105),
.B2(n_5),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_105),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_3),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_3),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_158),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_114),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_173),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_152),
.C(n_150),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_109),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_147),
.B1(n_151),
.B2(n_138),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_111),
.B1(n_119),
.B2(n_120),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_174),
.B1(n_142),
.B2(n_152),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_111),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_111),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_3),
.B(n_4),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_167),
.C(n_172),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_151),
.B1(n_136),
.B2(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_152),
.B1(n_153),
.B2(n_138),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_157),
.B1(n_166),
.B2(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_165),
.C(n_173),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_148),
.B1(n_140),
.B2(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_148),
.B(n_8),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_156),
.B(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_165),
.C(n_171),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_175),
.C(n_184),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_166),
.C(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_178),
.C(n_179),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_188),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_185),
.B(n_187),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_202),
.C(n_204),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_198),
.A2(n_185),
.B(n_193),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_13),
.B(n_10),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_181),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_207),
.C(n_7),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_176),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_180),
.C(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_214),
.B(n_7),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_206),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_207),
.C(n_201),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_157),
.B1(n_8),
.B2(n_9),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_204),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_205),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_10),
.C(n_12),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_220),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_210),
.C(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_217),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_223),
.B(n_224),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_227),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_216),
.Y(n_229)
);


endmodule