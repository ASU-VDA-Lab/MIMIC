module fake_jpeg_26347_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_28),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_28),
.Y(n_90)
);

BUFx2_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_51),
.B(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_23),
.C(n_17),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_17),
.C(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_35),
.B1(n_32),
.B2(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_26),
.B1(n_19),
.B2(n_20),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_68),
.B(n_76),
.Y(n_122)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_23),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_34),
.B(n_22),
.C(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_86),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_35),
.B1(n_32),
.B2(n_17),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_87),
.B1(n_20),
.B2(n_31),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_77),
.B(n_79),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_32),
.B1(n_35),
.B2(n_18),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_78),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_84),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_21),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_97),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_25),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_31),
.Y(n_131)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_28),
.B1(n_19),
.B2(n_30),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_109),
.B1(n_123),
.B2(n_98),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_27),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_69),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_131),
.C(n_89),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_39),
.B1(n_31),
.B2(n_0),
.Y(n_123)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_134),
.B(n_137),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_80),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_158),
.Y(n_182)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_74),
.B(n_89),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_126),
.B(n_123),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_148),
.B1(n_127),
.B2(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_71),
.B1(n_81),
.B2(n_95),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_159),
.B1(n_107),
.B2(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_149),
.B(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_104),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_150),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_147),
.B(n_151),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_101),
.B1(n_85),
.B2(n_83),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_98),
.B(n_88),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_113),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_68),
.C(n_82),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_158),
.C(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_94),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_79),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_84),
.B1(n_76),
.B2(n_96),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_160),
.B1(n_124),
.B2(n_121),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_109),
.B(n_31),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_39),
.C(n_93),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_108),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_1),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_164),
.A2(n_188),
.B(n_144),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_126),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_182),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_170),
.B1(n_176),
.B2(n_186),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_129),
.B(n_114),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_185),
.B(n_187),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_175),
.B(n_189),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_129),
.B1(n_114),
.B2(n_121),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_136),
.B1(n_8),
.B2(n_9),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_149),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_107),
.B(n_2),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_4),
.B(n_5),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_6),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_160),
.B1(n_157),
.B2(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_181),
.C(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_184),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_198),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_209),
.B1(n_215),
.B2(n_188),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_140),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_173),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_134),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_154),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_214),
.B1(n_197),
.B2(n_165),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_187),
.B(n_7),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_16),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_16),
.B(n_10),
.C(n_12),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_210),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_219),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_202),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_188),
.B1(n_186),
.B2(n_164),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_190),
.B1(n_171),
.B2(n_168),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_168),
.B1(n_163),
.B2(n_187),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_203),
.C(n_192),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_250),
.C(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_240),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_223),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_244),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_242),
.B1(n_249),
.B2(n_216),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_247),
.B1(n_233),
.B2(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_232),
.Y(n_247)
);

FAx1_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_210),
.CI(n_208),
.CON(n_249),
.SN(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_196),
.C(n_207),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_229),
.B(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_222),
.C(n_217),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_255),
.C(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_222),
.C(n_193),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_198),
.B1(n_194),
.B2(n_199),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_213),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_204),
.B1(n_221),
.B2(n_202),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_228),
.B1(n_195),
.B2(n_216),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_246),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_249),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_263),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_264),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_242),
.B1(n_258),
.B2(n_259),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_248),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_256),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_271),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_257),
.B(n_262),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_205),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_252),
.B(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_279),
.C(n_268),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_265),
.B(n_255),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_282),
.B(n_267),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_163),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_285),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_212),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_277),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_287),
.A2(n_284),
.B(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_289),
.B(n_10),
.Y(n_293)
);

AOI332xp33_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_9),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.B3(n_15),
.C1(n_147),
.C2(n_220),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);


endmodule