module fake_netlist_1_11801_n_656 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_656);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_656;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_68), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_76), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_42), .Y(n_79) );
BUFx6f_ASAP7_75t_L g80 ( .A(n_64), .Y(n_80) );
INVx2_ASAP7_75t_SL g81 ( .A(n_18), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_1), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_23), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_15), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_39), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_20), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_40), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_36), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_3), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_9), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_62), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_67), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_5), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_8), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_75), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_24), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
BUFx10_ASAP7_75t_L g99 ( .A(n_61), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_71), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_31), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_74), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_14), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_5), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_56), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_13), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_13), .Y(n_107) );
BUFx5_ASAP7_75t_L g108 ( .A(n_58), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_29), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_6), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_10), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_60), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_19), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_53), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_7), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_116), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_80), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_107), .B(n_0), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_99), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_108), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_81), .B(n_1), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_102), .B(n_2), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_104), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_81), .B(n_3), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_108), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_112), .B(n_4), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_108), .B(n_6), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
CKINVDCx6p67_ASAP7_75t_R g141 ( .A(n_99), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_104), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_114), .B(n_7), .Y(n_143) );
BUFx12f_ASAP7_75t_L g144 ( .A(n_78), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_114), .B(n_9), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_107), .B(n_11), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_93), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_117), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_80), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_119), .B(n_11), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_119), .B(n_12), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_117), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_77), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
BUFx10_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_121), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_127), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_125), .B(n_102), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_122), .B(n_83), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_122), .B(n_83), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_125), .B(n_126), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_125), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_148), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
NAND2xp33_ASAP7_75t_L g172 ( .A(n_125), .B(n_108), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_155), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_131), .Y(n_176) );
INVxp67_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_126), .B(n_78), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_126), .B(n_105), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_153), .A2(n_82), .B1(n_113), .B2(n_84), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_126), .B(n_105), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_141), .B(n_92), .Y(n_183) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_123), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_124), .B(n_118), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_154), .A2(n_90), .B1(n_109), .B2(n_98), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_146), .B(n_106), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_141), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_123), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_130), .B(n_103), .Y(n_194) );
INVx8_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_123), .Y(n_196) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_124), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_130), .B(n_110), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_128), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_156), .B(n_92), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_123), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_176), .B(n_143), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_158), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_161), .B(n_128), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_195), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_161), .B(n_132), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_197), .B(n_144), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_179), .B(n_132), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_199), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_199), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_162), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_195), .A2(n_156), .B1(n_134), .B2(n_129), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_180), .B(n_134), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_197), .B(n_144), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_182), .B(n_120), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_197), .B(n_133), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_195), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_175), .A2(n_139), .B(n_145), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_195), .A2(n_166), .B1(n_167), .B2(n_184), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_163), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_195), .B(n_137), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_175), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_168), .B(n_152), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_191), .B(n_152), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_163), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_183), .B(n_138), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_157), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_166), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_178), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_178), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_158), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_186), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_186), .Y(n_237) );
BUFx4f_ASAP7_75t_L g238 ( .A(n_166), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_189), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_191), .B(n_138), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_191), .B(n_140), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_158), .Y(n_242) );
NOR2xp33_ASAP7_75t_R g243 ( .A(n_192), .B(n_94), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_191), .B(n_140), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_166), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_194), .B(n_147), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_166), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_166), .A2(n_147), .B1(n_150), .B2(n_149), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_194), .B(n_149), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_184), .B(n_97), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_184), .B(n_96), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_157), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_198), .B(n_150), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_169), .B(n_95), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_198), .B(n_12), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_160), .Y(n_256) );
OR2x6_ASAP7_75t_L g257 ( .A(n_206), .B(n_165), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_211), .A2(n_165), .B(n_173), .C(n_185), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_202), .A2(n_170), .B1(n_174), .B2(n_94), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_211), .A2(n_165), .B(n_185), .C(n_173), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_212), .A2(n_215), .B(n_210), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_228), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_206), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_206), .B(n_173), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_220), .B(n_158), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_220), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_255), .A2(n_189), .B(n_188), .C(n_200), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_256), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_208), .B(n_181), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_243), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_228), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_212), .A2(n_160), .B(n_190), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_220), .B(n_185), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_214), .A2(n_169), .B1(n_79), .B2(n_85), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_205), .A2(n_172), .B(n_88), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_228), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_214), .B(n_166), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_218), .B(n_167), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_246), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_253), .A2(n_91), .B1(n_101), .B2(n_111), .C(n_100), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_253), .B(n_167), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_223), .A2(n_100), .B1(n_167), .B2(n_80), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_202), .Y(n_284) );
NAND2x1_ASAP7_75t_SL g285 ( .A(n_235), .B(n_167), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_232), .B(n_167), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_218), .A2(n_201), .B(n_196), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_256), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_249), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_255), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_209), .B(n_167), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_232), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_240), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_241), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_244), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_207), .A2(n_187), .B(n_196), .Y(n_296) );
NOR2x1_ASAP7_75t_L g297 ( .A(n_216), .B(n_201), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_232), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_221), .A2(n_135), .B(n_121), .C(n_151), .Y(n_299) );
INVx3_ASAP7_75t_SL g300 ( .A(n_245), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_225), .A2(n_187), .B(n_196), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_221), .B(n_108), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_226), .A2(n_201), .B(n_193), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_226), .B(n_108), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_280), .B(n_245), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_303), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_287), .A2(n_233), .B(n_236), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_284), .B(n_230), .Y(n_310) );
OR2x6_ASAP7_75t_L g311 ( .A(n_286), .B(n_247), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_262), .A2(n_238), .B(n_219), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_259), .A2(n_217), .B(n_248), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_304), .A2(n_234), .B(n_236), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_257), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_284), .B(n_233), .Y(n_317) );
AO21x1_ASAP7_75t_L g318 ( .A1(n_283), .A2(n_234), .B(n_237), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_302), .A2(n_237), .B(n_239), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_289), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_258), .A2(n_239), .B(n_252), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_290), .B(n_231), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_305), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_286), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_270), .B(n_231), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_267), .B(n_245), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_305), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_293), .B(n_252), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_260), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_296), .A2(n_254), .B(n_227), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_279), .A2(n_238), .B(n_250), .Y(n_333) );
AO21x2_ASAP7_75t_L g334 ( .A1(n_261), .A2(n_222), .B(n_251), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_299), .A2(n_229), .B(n_203), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_294), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_279), .A2(n_229), .B(n_203), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_320), .A2(n_271), .B1(n_278), .B2(n_286), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_306), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_310), .B(n_275), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
AOI22xp33_ASAP7_75t_SL g343 ( .A1(n_316), .A2(n_275), .B1(n_298), .B2(n_278), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_330), .A2(n_282), .B1(n_257), .B2(n_283), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
AO21x2_ASAP7_75t_L g346 ( .A1(n_318), .A2(n_276), .B(n_222), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_337), .B(n_295), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_330), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_337), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_309), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_327), .B(n_272), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_327), .B(n_277), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_326), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_316), .A2(n_247), .B1(n_291), .B2(n_257), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_313), .B(n_229), .Y(n_355) );
OAI321xp33_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_281), .A3(n_268), .B1(n_151), .B2(n_135), .C(n_121), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_314), .A2(n_291), .B1(n_265), .B2(n_264), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
OAI211xp5_ASAP7_75t_L g359 ( .A1(n_317), .A2(n_297), .B(n_285), .C(n_274), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_326), .B(n_267), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_324), .A2(n_265), .B1(n_264), .B2(n_247), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_331), .B(n_267), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_324), .A2(n_222), .B1(n_238), .B2(n_292), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_325), .A2(n_245), .B1(n_204), .B2(n_242), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_321), .A2(n_301), .B(n_235), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_342), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g367 ( .A1(n_341), .A2(n_325), .B1(n_329), .B2(n_313), .C(n_335), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_350), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_342), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_345), .B(n_318), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_350), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_353), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_358), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_340), .B(n_326), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_348), .B(n_309), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_345), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_348), .B(n_331), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_353), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_341), .B(n_321), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_355), .B(n_335), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_365), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_353), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_355), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_349), .B(n_329), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_360), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_349), .B(n_334), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_340), .B(n_334), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_362), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_347), .B(n_334), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_353), .Y(n_391) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_360), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_340), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_360), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_346), .Y(n_396) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_392), .B(n_346), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_383), .B(n_346), .Y(n_398) );
NAND4xp25_ASAP7_75t_L g399 ( .A(n_367), .B(n_343), .C(n_357), .D(n_354), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_383), .B(n_108), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
AOI33xp33_ASAP7_75t_L g402 ( .A1(n_366), .A2(n_339), .A3(n_363), .B1(n_361), .B2(n_16), .B3(n_15), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_373), .A2(n_352), .B1(n_351), .B2(n_359), .C(n_344), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_379), .B(n_360), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_366), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_387), .B(n_326), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_369), .B(n_319), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_376), .B(n_319), .Y(n_410) );
AND2x4_ASAP7_75t_SL g411 ( .A(n_374), .B(n_311), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_380), .Y(n_414) );
INVx4_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_368), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_386), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_389), .A2(n_326), .B1(n_311), .B2(n_306), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_368), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_387), .B(n_336), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_378), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_382), .B(n_356), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_371), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g426 ( .A(n_367), .B(n_312), .C(n_333), .D(n_16), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_370), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_371), .B(n_375), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_371), .B(n_336), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_377), .B(n_326), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_375), .B(n_336), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_370), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_377), .B(n_336), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_384), .A2(n_311), .B1(n_306), .B2(n_364), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_379), .B(n_332), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_384), .A2(n_311), .B1(n_306), .B2(n_338), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_390), .B(n_14), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_413), .B(n_393), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_398), .B(n_396), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_403), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_414), .B(n_393), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_398), .B(n_396), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_419), .B(n_385), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_397), .B(n_395), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_405), .B(n_385), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_436), .B(n_388), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_437), .B(n_395), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_409), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_437), .B(n_395), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_409), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_412), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_439), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_428), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_439), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_400), .B(n_395), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_408), .Y(n_463) );
OAI211xp5_ASAP7_75t_L g464 ( .A1(n_399), .A2(n_382), .B(n_372), .C(n_395), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_434), .B(n_395), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_424), .A2(n_356), .B(n_394), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_434), .B(n_395), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_408), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_422), .B(n_394), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_422), .B(n_394), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_436), .B(n_392), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_432), .B(n_381), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_401), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g474 ( .A1(n_399), .A2(n_382), .B1(n_372), .B2(n_391), .C(n_381), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_415), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_410), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_430), .Y(n_477) );
OAI31xp33_ASAP7_75t_L g478 ( .A1(n_426), .A2(n_374), .A3(n_391), .B(n_372), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_432), .B(n_417), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_430), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_427), .B(n_374), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_417), .B(n_381), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_410), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_430), .Y(n_484) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_435), .A2(n_374), .B(n_372), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_420), .B(n_391), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_405), .B(n_332), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_420), .B(n_151), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_401), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_427), .B(n_151), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_426), .A2(n_311), .B1(n_151), .B2(n_135), .C(n_121), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_397), .B(n_135), .Y(n_493) );
INVx4_ASAP7_75t_L g494 ( .A(n_415), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_415), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_458), .B(n_423), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_457), .B(n_433), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_444), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_475), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_473), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_459), .B(n_433), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_460), .B(n_423), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_452), .Y(n_505) );
OAI21xp33_ASAP7_75t_L g506 ( .A1(n_464), .A2(n_402), .B(n_135), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_479), .B(n_407), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_465), .B(n_429), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_492), .A2(n_418), .B1(n_415), .B2(n_404), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_447), .B(n_438), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_485), .B(n_431), .C(n_407), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_473), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_477), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_479), .B(n_429), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_463), .B(n_421), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_468), .B(n_421), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_476), .B(n_425), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_455), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_456), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_475), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_483), .B(n_425), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_441), .B(n_416), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_494), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_494), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_489), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_441), .B(n_407), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_494), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_446), .B(n_407), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_450), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_465), .B(n_467), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_446), .B(n_411), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_475), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_450), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_440), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_461), .B(n_411), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_445), .B(n_411), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_467), .B(n_451), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_481), .B(n_135), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_482), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_491), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_495), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_482), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_469), .B(n_121), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_486), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_486), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_480), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_471), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_471), .B(n_121), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_542), .B(n_469), .Y(n_552) );
OAI22xp33_ASAP7_75t_L g553 ( .A1(n_524), .A2(n_495), .B1(n_484), .B2(n_487), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_510), .A2(n_478), .B1(n_451), .B2(n_453), .Y(n_554) );
NOR3xp33_ASAP7_75t_SL g555 ( .A(n_509), .B(n_474), .C(n_466), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_502), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_497), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_525), .A2(n_495), .B1(n_453), .B2(n_493), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g559 ( .A1(n_511), .A2(n_462), .B1(n_449), .B2(n_488), .C(n_470), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_498), .Y(n_560) );
OAI32xp33_ASAP7_75t_L g561 ( .A1(n_511), .A2(n_470), .A3(n_472), .B1(n_488), .B2(n_448), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_539), .B(n_472), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_506), .A2(n_493), .B(n_448), .C(n_328), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_500), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_515), .B(n_448), .Y(n_565) );
OAI211xp5_ASAP7_75t_SL g566 ( .A1(n_535), .A2(n_171), .B(n_193), .C(n_201), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_545), .B(n_493), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_549), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_523), .B(n_315), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_505), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_512), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_520), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_519), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_530), .B(n_315), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_531), .B(n_17), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_507), .B(n_21), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_534), .B(n_519), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_514), .B(n_22), .Y(n_578) );
INVx3_ASAP7_75t_L g579 ( .A(n_501), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_525), .A2(n_235), .B(n_266), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_540), .B(n_171), .C(n_193), .Y(n_581) );
AOI221xp5_ASAP7_75t_SL g582 ( .A1(n_510), .A2(n_171), .B1(n_159), .B2(n_27), .C(n_28), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_549), .B(n_25), .Y(n_583) );
NAND3x2_ASAP7_75t_L g584 ( .A(n_504), .B(n_26), .C(n_30), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_499), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_496), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_503), .B(n_308), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_526), .B(n_543), .Y(n_588) );
AOI221x1_ASAP7_75t_L g589 ( .A1(n_540), .A2(n_159), .B1(n_224), .B2(n_213), .C(n_35), .Y(n_589) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_528), .B(n_245), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_547), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_528), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_554), .A2(n_537), .B1(n_550), .B2(n_548), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_592), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_585), .B(n_508), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_577), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_555), .A2(n_521), .B(n_501), .C(n_544), .Y(n_597) );
XNOR2xp5_ASAP7_75t_L g598 ( .A(n_586), .B(n_529), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_561), .A2(n_527), .B(n_532), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_557), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_591), .B(n_508), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_552), .B(n_518), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_577), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_562), .B(n_544), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_568), .Y(n_605) );
XOR2xp5_ASAP7_75t_L g606 ( .A(n_575), .B(n_536), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_588), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_559), .A2(n_533), .B1(n_551), .B2(n_537), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_558), .A2(n_533), .B1(n_538), .B2(n_541), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_552), .B(n_502), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_553), .A2(n_546), .B1(n_517), .B2(n_522), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_579), .B(n_526), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_560), .A2(n_516), .B1(n_543), .B2(n_513), .C(n_159), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_564), .B(n_513), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_584), .A2(n_245), .B1(n_300), .B2(n_235), .Y(n_616) );
OAI322xp33_ASAP7_75t_L g617 ( .A1(n_565), .A2(n_159), .A3(n_224), .B1(n_213), .B2(n_37), .C1(n_38), .C2(n_41), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_596), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_603), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_594), .B(n_571), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_609), .B(n_579), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_599), .A2(n_576), .B1(n_581), .B2(n_567), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_597), .A2(n_563), .B(n_578), .C(n_582), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_608), .A2(n_567), .B(n_556), .Y(n_624) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_616), .B(n_583), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_594), .A2(n_570), .B(n_572), .C(n_580), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_610), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_605), .A2(n_566), .B(n_590), .C(n_574), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g629 ( .A1(n_600), .A2(n_573), .B1(n_574), .B2(n_587), .C1(n_569), .C2(n_589), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_615), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_616), .A2(n_587), .B(n_590), .Y(n_631) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_617), .B(n_32), .Y(n_632) );
OAI311xp33_ASAP7_75t_L g633 ( .A1(n_629), .A2(n_593), .A3(n_611), .B1(n_613), .C1(n_595), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_621), .A2(n_606), .B(n_598), .Y(n_634) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_622), .A2(n_602), .B1(n_601), .B2(n_604), .C(n_607), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_618), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_626), .A2(n_614), .B1(n_612), .B2(n_159), .C(n_44), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_632), .B(n_308), .C(n_242), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_625), .B(n_33), .Y(n_639) );
AOI321xp33_ASAP7_75t_L g640 ( .A1(n_622), .A2(n_34), .A3(n_43), .B1(n_45), .B2(n_46), .C(n_47), .Y(n_640) );
NAND3xp33_ASAP7_75t_SL g641 ( .A(n_623), .B(n_48), .C(n_49), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_634), .B(n_627), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_636), .B(n_630), .Y(n_643) );
INVx4_ASAP7_75t_L g644 ( .A(n_640), .Y(n_644) );
XNOR2x1_ASAP7_75t_L g645 ( .A(n_639), .B(n_619), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_633), .A2(n_624), .B1(n_628), .B2(n_620), .C(n_631), .Y(n_646) );
OAI31xp33_ASAP7_75t_L g647 ( .A1(n_642), .A2(n_638), .A3(n_635), .B(n_641), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_645), .B(n_637), .Y(n_648) );
OAI222xp33_ASAP7_75t_L g649 ( .A1(n_644), .A2(n_50), .B1(n_51), .B2(n_52), .C1(n_54), .C2(n_55), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_647), .A2(n_646), .B(n_643), .Y(n_650) );
OAI31xp33_ASAP7_75t_SL g651 ( .A1(n_648), .A2(n_57), .A3(n_59), .B(n_63), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_650), .Y(n_652) );
AOI222xp33_ASAP7_75t_SL g653 ( .A1(n_652), .A2(n_647), .B1(n_651), .B2(n_648), .C1(n_649), .C2(n_73), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_653), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_204), .B1(n_66), .B2(n_70), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_65), .B(n_72), .Y(n_656) );
endmodule