module fake_jpeg_28038_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_33),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_20),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_55),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_31),
.B1(n_27),
.B2(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_56),
.B1(n_61),
.B2(n_44),
.Y(n_73)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_24),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_31),
.B1(n_27),
.B2(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_62),
.Y(n_86)
);

AO22x1_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_28),
.B1(n_32),
.B2(n_19),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_62),
.B1(n_49),
.B2(n_58),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.C(n_19),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_28),
.Y(n_63)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_39),
.A3(n_36),
.B1(n_17),
.B2(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_45),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_82),
.Y(n_108)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_76),
.Y(n_104)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_75),
.Y(n_90)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_26),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_88),
.CON(n_103),
.SN(n_103)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_45),
.B1(n_19),
.B2(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_49),
.B1(n_54),
.B2(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_87),
.B1(n_78),
.B2(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_30),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_22),
.B1(n_23),
.B2(n_16),
.Y(n_87)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_39),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_47),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_66),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_25),
.Y(n_124)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_97),
.CON(n_127),
.SN(n_127)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_48),
.B1(n_25),
.B2(n_16),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_53),
.B(n_25),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_108),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_80),
.C(n_85),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_132),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_80),
.C(n_89),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_92),
.C(n_4),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_72),
.B1(n_75),
.B2(n_69),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_98),
.B(n_111),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_125),
.B(n_101),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_79),
.B1(n_48),
.B2(n_22),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_126),
.B1(n_134),
.B2(n_113),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_21),
.B1(n_29),
.B2(n_2),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_1),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_109),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_112),
.B(n_106),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_107),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_144),
.B(n_155),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_94),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_147),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_121),
.B1(n_134),
.B2(n_5),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_123),
.B1(n_126),
.B2(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_96),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_156),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_128),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_96),
.B(n_92),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_116),
.C(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_157),
.B(n_158),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_133),
.C(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_151),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_124),
.C(n_119),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_166),
.B1(n_168),
.B2(n_171),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_170),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_127),
.B(n_122),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_161),
.C(n_156),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_140),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_160),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_145),
.B1(n_136),
.B2(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_152),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_148),
.B(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_150),
.B1(n_137),
.B2(n_144),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_187),
.A2(n_169),
.B1(n_168),
.B2(n_153),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_165),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_191),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_195),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_156),
.C(n_154),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_179),
.C(n_184),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_171),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_196),
.A2(n_177),
.B(n_185),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_176),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_198),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_14),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_205),
.B(n_186),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_191),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_183),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_189),
.B1(n_205),
.B2(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_208),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_210),
.A2(n_5),
.B(n_6),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_190),
.C(n_148),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_212),
.B(n_213),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_148),
.C(n_147),
.Y(n_212)
);

AOI21x1_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_13),
.B(n_6),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_217),
.C(n_9),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_13),
.B(n_6),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_211),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_221),
.B(n_218),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_9),
.B(n_10),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_222),
.B(n_10),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_11),
.Y(n_226)
);


endmodule