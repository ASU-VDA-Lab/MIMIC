module fake_jpeg_9329_n_61 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_61);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_61;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_7),
.C(n_6),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_34),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_23),
.B1(n_10),
.B2(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_26),
.B1(n_25),
.B2(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_0),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_37),
.B(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_2),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_30),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_25),
.C(n_29),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_49),
.C(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_12),
.B1(n_19),
.B2(n_18),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_13),
.C(n_20),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_53),
.B(n_46),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_50),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_54),
.B2(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_57),
.B(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_40),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_44),
.B(n_47),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_41),
.Y(n_61)
);


endmodule