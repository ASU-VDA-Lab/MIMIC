module fake_jpeg_10208_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_181;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_21),
.Y(n_66)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_20),
.C(n_23),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_22),
.B1(n_34),
.B2(n_18),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_5),
.B(n_6),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_18),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_61),
.B(n_24),
.Y(n_73)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_22),
.B1(n_20),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_30),
.B1(n_31),
.B2(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_66),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_34),
.B1(n_18),
.B2(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_82)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_70),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_31),
.B(n_28),
.C(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_34),
.B1(n_30),
.B2(n_21),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_76),
.B1(n_89),
.B2(n_91),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_64),
.B(n_47),
.C(n_59),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_5),
.Y(n_118)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_30),
.B1(n_24),
.B2(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_36),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_101),
.B1(n_5),
.B2(n_6),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_96),
.B1(n_56),
.B2(n_54),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_88),
.Y(n_120)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_36),
.B(n_32),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_45),
.C(n_47),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_32),
.B1(n_37),
.B2(n_3),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_7),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_85),
.B(n_83),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_46),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_126),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_60),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_84),
.C(n_77),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_54),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_94),
.B1(n_75),
.B2(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_127),
.B1(n_99),
.B2(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_16),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_85),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_70),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_14),
.B1(n_9),
.B2(n_10),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_111),
.B(n_109),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_144),
.B(n_148),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_95),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_153),
.C(n_105),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_125),
.A2(n_87),
.B1(n_69),
.B2(n_94),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_136),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_141),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_98),
.B(n_86),
.C(n_81),
.D(n_68),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_145),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_83),
.B(n_100),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_106),
.B(n_108),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_154),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_145),
.B(n_126),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_119),
.B(n_108),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_127),
.B(n_96),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_166),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_116),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_167),
.C(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_176),
.B1(n_143),
.B2(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_154),
.B1(n_148),
.B2(n_105),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_192),
.B1(n_162),
.B2(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_181),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_149),
.A3(n_129),
.B1(n_131),
.B2(n_141),
.C1(n_128),
.C2(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_194),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_106),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_191),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_128),
.B1(n_110),
.B2(n_69),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_125),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_187),
.C(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_107),
.C(n_114),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_107),
.C(n_140),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_173),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_110),
.B1(n_69),
.B2(n_140),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_171),
.B(n_161),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_97),
.A3(n_134),
.B1(n_14),
.B2(n_12),
.C1(n_8),
.C2(n_11),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_161),
.CI(n_159),
.CON(n_198),
.SN(n_198)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_202),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_210),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_174),
.B1(n_155),
.B2(n_158),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_204),
.B1(n_189),
.B2(n_165),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_205),
.B(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_174),
.B1(n_168),
.B2(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_156),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_187),
.C(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_220),
.C(n_222),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_204),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_223),
.B(n_205),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_221),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_193),
.B1(n_181),
.B2(n_184),
.Y(n_217)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_192),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_183),
.B(n_169),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_211),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_183),
.B(n_12),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_207),
.C(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_217),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_198),
.C(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_233),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_218),
.B1(n_219),
.B2(n_223),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_235),
.A2(n_230),
.B(n_231),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_238),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_241),
.A2(n_239),
.B1(n_234),
.B2(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_13),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_198),
.B(n_13),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_247),
.A2(n_248),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_245),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_13),
.Y(n_251)
);


endmodule