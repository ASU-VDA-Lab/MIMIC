module fake_ariane_1889_n_2088 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2088);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2088;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_600;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_1906;
wire n_1899;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1733;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_1789;
wire n_763;
wire n_1986;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_1252;
wire n_1129;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx3_ASAP7_75t_L g547 ( 
.A(n_146),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_77),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_259),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_115),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_514),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_288),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_378),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_456),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_448),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_356),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_382),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_255),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_430),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_160),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_317),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_543),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_272),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_270),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_283),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_312),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_56),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_88),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_284),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_25),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_526),
.Y(n_571)
);

BUFx5_ASAP7_75t_L g572 ( 
.A(n_36),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_322),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_169),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_219),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_426),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_46),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_14),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_238),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_168),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_429),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_85),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_204),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_154),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_340),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_535),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_483),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_221),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_501),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_290),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_394),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_540),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_527),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_386),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_85),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_84),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_266),
.Y(n_598)
);

CKINVDCx14_ASAP7_75t_R g599 ( 
.A(n_61),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_491),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_118),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_189),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_537),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_137),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_218),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_410),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_141),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_330),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_244),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_442),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_24),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_390),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_479),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_90),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_468),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_62),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_464),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_353),
.Y(n_618)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_506),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_342),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_169),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_329),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_305),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_498),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_12),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_380),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_409),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_297),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_517),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_158),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_121),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_338),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_497),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_331),
.Y(n_634)
);

BUFx10_ASAP7_75t_L g635 ( 
.A(n_84),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_231),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_11),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_117),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_391),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_250),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_190),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_110),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_162),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_166),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_105),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_325),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_327),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_267),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_66),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_332),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_421),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_499),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_337),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_128),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_511),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_310),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_70),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_26),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_237),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_196),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_485),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_34),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_293),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_201),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_53),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_120),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_116),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_113),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_437),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_411),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_248),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_157),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_241),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_18),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_67),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_42),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_279),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_217),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_147),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_484),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_211),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_170),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_359),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_98),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_14),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_113),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_323),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_339),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_295),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_404),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_9),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_111),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_181),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_434),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_363),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_400),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_182),
.Y(n_697)
);

CKINVDCx16_ASAP7_75t_R g698 ( 
.A(n_44),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_408),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_423),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_53),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_31),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_6),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_412),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_185),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_350),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_72),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_367),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_21),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_167),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_320),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_528),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_149),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_402),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_173),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_374),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_531),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_276),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_455),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_152),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_472),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_466),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_162),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_541),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_82),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_77),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_64),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_444),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_41),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_64),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_242),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_131),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_107),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_95),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_247),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_40),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_346),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_306),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_301),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_433),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_102),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_333),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_265),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_251),
.Y(n_744)
);

CKINVDCx16_ASAP7_75t_R g745 ( 
.A(n_271),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_533),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_495),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_177),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_281),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_364),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_299),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_120),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_8),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_233),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_507),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_547),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_547),
.Y(n_757)
);

INVxp33_ASAP7_75t_SL g758 ( 
.A(n_548),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_607),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_607),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_698),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_657),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_657),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_572),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_572),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_638),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_572),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_572),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_726),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_668),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_572),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_668),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_668),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_564),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_727),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_572),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_668),
.Y(n_777)
);

INVxp33_ASAP7_75t_SL g778 ( 
.A(n_550),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_732),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_576),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_606),
.Y(n_781)
);

CKINVDCx16_ASAP7_75t_R g782 ( 
.A(n_599),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_596),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_730),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_745),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_596),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_730),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_577),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_601),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_614),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_568),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_615),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_631),
.Y(n_793)
);

CKINVDCx16_ASAP7_75t_R g794 ( 
.A(n_635),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_653),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_730),
.Y(n_797)
);

INVxp33_ASAP7_75t_SL g798 ( 
.A(n_570),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_733),
.Y(n_799)
);

INVxp33_ASAP7_75t_SL g800 ( 
.A(n_574),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_616),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_677),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_681),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_621),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_630),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_662),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_573),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_665),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_666),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_635),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_573),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_667),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_728),
.Y(n_813)
);

INVxp33_ASAP7_75t_SL g814 ( 
.A(n_578),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_733),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_738),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_742),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_672),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_679),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_682),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_691),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_734),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_741),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_751),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_752),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_581),
.Y(n_826)
);

CKINVDCx14_ASAP7_75t_R g827 ( 
.A(n_623),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_567),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_560),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_583),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_585),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_683),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_597),
.Y(n_833)
);

INVxp33_ASAP7_75t_L g834 ( 
.A(n_619),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_623),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_549),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_554),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_604),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_565),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_713),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_575),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_580),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_582),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_611),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_584),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_587),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_793),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_834),
.B(n_683),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_770),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_SL g850 ( 
.A1(n_766),
.A2(n_775),
.B1(n_769),
.B2(n_813),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_772),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_773),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_763),
.B(n_592),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_784),
.Y(n_854)
);

OA21x2_ASAP7_75t_L g855 ( 
.A1(n_764),
.A2(n_608),
.B(n_593),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_807),
.B(n_609),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_834),
.B(n_553),
.Y(n_857)
);

NAND2xp33_ASAP7_75t_L g858 ( 
.A(n_836),
.B(n_598),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_784),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_777),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_785),
.A2(n_625),
.B1(n_654),
.B2(n_645),
.Y(n_861)
);

OA21x2_ASAP7_75t_L g862 ( 
.A1(n_765),
.A2(n_622),
.B(n_620),
.Y(n_862)
);

OA21x2_ASAP7_75t_L g863 ( 
.A1(n_767),
.A2(n_771),
.B(n_768),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_787),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_807),
.B(n_632),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_761),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_787),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_811),
.B(n_553),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_811),
.B(n_618),
.Y(n_869)
);

BUFx8_ASAP7_75t_L g870 ( 
.A(n_835),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_776),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_774),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_795),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_795),
.Y(n_874)
);

BUFx8_ASAP7_75t_SL g875 ( 
.A(n_766),
.Y(n_875)
);

INVx5_ASAP7_75t_L g876 ( 
.A(n_777),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_782),
.Y(n_877)
);

OAI22x1_ASAP7_75t_L g878 ( 
.A1(n_779),
.A2(n_642),
.B1(n_643),
.B2(n_637),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_832),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_788),
.Y(n_880)
);

OA21x2_ASAP7_75t_L g881 ( 
.A1(n_837),
.A2(n_641),
.B(n_636),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_789),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_790),
.Y(n_883)
);

BUFx8_ASAP7_75t_L g884 ( 
.A(n_832),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_801),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_797),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_804),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_805),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_830),
.B(n_556),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_797),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_839),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_841),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_842),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_843),
.Y(n_894)
);

AND2x2_ASAP7_75t_SL g895 ( 
.A(n_786),
.B(n_618),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_845),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_806),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_826),
.Y(n_898)
);

AND2x6_ASAP7_75t_L g899 ( 
.A(n_846),
.B(n_626),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_808),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_791),
.Y(n_901)
);

OA21x2_ASAP7_75t_L g902 ( 
.A1(n_809),
.A2(n_651),
.B(n_650),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_827),
.B(n_652),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_812),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_879),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_903),
.B(n_758),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_863),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_863),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_863),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_879),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_880),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_859),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_895),
.B(n_626),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_895),
.B(n_891),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_882),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_859),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_886),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_883),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_872),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_849),
.B(n_778),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_L g921 ( 
.A(n_871),
.B(n_844),
.Y(n_921)
);

CKINVDCx6p67_ASAP7_75t_R g922 ( 
.A(n_847),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_891),
.B(n_798),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_848),
.B(n_827),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_885),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_887),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_864),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_877),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_851),
.B(n_800),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_852),
.B(n_833),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_901),
.B(n_794),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_L g932 ( 
.A(n_899),
.B(n_831),
.Y(n_932)
);

INVx6_ASAP7_75t_L g933 ( 
.A(n_884),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_867),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_891),
.B(n_893),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_L g936 ( 
.A(n_899),
.B(n_598),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_877),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_898),
.B(n_838),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_867),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_891),
.B(n_798),
.Y(n_940)
);

INVxp33_ASAP7_75t_SL g941 ( 
.A(n_872),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_SL g942 ( 
.A(n_893),
.B(n_644),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_888),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_886),
.Y(n_944)
);

INVxp33_ASAP7_75t_L g945 ( 
.A(n_866),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_873),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_873),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_874),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_874),
.Y(n_949)
);

AO21x2_ASAP7_75t_L g950 ( 
.A1(n_857),
.A2(n_669),
.B(n_655),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_889),
.B(n_814),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_L g952 ( 
.A(n_899),
.B(n_598),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_886),
.Y(n_953)
);

BUFx6f_ASAP7_75t_SL g954 ( 
.A(n_868),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_897),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_854),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_875),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_889),
.B(n_814),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_855),
.A2(n_688),
.B(n_670),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_893),
.B(n_689),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_854),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_877),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_900),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_857),
.A2(n_697),
.B(n_695),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_854),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_884),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_890),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_893),
.B(n_699),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_892),
.B(n_815),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_899),
.Y(n_970)
);

OA22x2_ASAP7_75t_L g971 ( 
.A1(n_878),
.A2(n_757),
.B1(n_759),
.B2(n_756),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_892),
.B(n_700),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_890),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_892),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_890),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_875),
.Y(n_976)
);

INVx8_ASAP7_75t_L g977 ( 
.A(n_899),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_886),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_L g979 ( 
.A(n_904),
.B(n_598),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_894),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_894),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_855),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_855),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_896),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_974),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_958),
.B(n_780),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_937),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_938),
.B(n_781),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_911),
.Y(n_989)
);

XNOR2x2_ASAP7_75t_L g990 ( 
.A(n_971),
.B(n_878),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_951),
.B(n_853),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_915),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_918),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_925),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_926),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_907),
.B(n_881),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_937),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_943),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_955),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_963),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_922),
.B(n_792),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_956),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_956),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_919),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_931),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_961),
.Y(n_1006)
);

XNOR2x2_ASAP7_75t_L g1007 ( 
.A(n_971),
.B(n_861),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_961),
.Y(n_1008)
);

INVx3_ASAP7_75t_R g1009 ( 
.A(n_957),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_907),
.B(n_881),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_965),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_928),
.B(n_896),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_965),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_962),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_967),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_908),
.B(n_909),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_973),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_912),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_973),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_975),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_966),
.B(n_799),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_975),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_908),
.B(n_881),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_945),
.B(n_796),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_906),
.B(n_884),
.Y(n_1025)
);

INVxp33_ASAP7_75t_L g1026 ( 
.A(n_945),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_980),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_930),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_913),
.B(n_802),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_981),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_984),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_959),
.A2(n_862),
.B(n_902),
.Y(n_1032)
);

XOR2xp5_ASAP7_75t_L g1033 ( 
.A(n_941),
.B(n_813),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_SL g1034 ( 
.A(n_913),
.B(n_870),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_905),
.Y(n_1035)
);

BUFx8_ASAP7_75t_L g1036 ( 
.A(n_976),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_910),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_924),
.B(n_803),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_912),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_923),
.B(n_940),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_916),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_916),
.Y(n_1042)
);

INVxp33_ASAP7_75t_L g1043 ( 
.A(n_920),
.Y(n_1043)
);

XOR2xp5_ASAP7_75t_L g1044 ( 
.A(n_914),
.B(n_816),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_929),
.B(n_824),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_927),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_927),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_953),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_934),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_923),
.B(n_850),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_934),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_909),
.B(n_902),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_939),
.Y(n_1053)
);

XNOR2xp5_ASAP7_75t_L g1054 ( 
.A(n_940),
.B(n_816),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_933),
.B(n_840),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_939),
.Y(n_1056)
);

XOR2xp5_ASAP7_75t_L g1057 ( 
.A(n_914),
.B(n_817),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_933),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_946),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_946),
.Y(n_1060)
);

XNOR2xp5_ASAP7_75t_L g1061 ( 
.A(n_942),
.B(n_817),
.Y(n_1061)
);

NAND2xp33_ASAP7_75t_R g1062 ( 
.A(n_982),
.B(n_862),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_947),
.Y(n_1063)
);

XNOR2xp5_ASAP7_75t_L g1064 ( 
.A(n_942),
.B(n_769),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_948),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_948),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_933),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_949),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_L g1069 ( 
.A(n_970),
.B(n_865),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_949),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_969),
.Y(n_1071)
);

INVxp33_ASAP7_75t_L g1072 ( 
.A(n_972),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_935),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_978),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_954),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_950),
.Y(n_1076)
);

XOR2x2_ASAP7_75t_L g1077 ( 
.A(n_950),
.B(n_775),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_935),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_972),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_960),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_960),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_968),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_964),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_921),
.B(n_856),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_968),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_921),
.B(n_783),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_L g1087 ( 
.A(n_970),
.B(n_868),
.Y(n_1087)
);

XOR2xp5_ASAP7_75t_L g1088 ( 
.A(n_953),
.B(n_783),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_964),
.Y(n_1089)
);

XNOR2x2_ASAP7_75t_L g1090 ( 
.A(n_954),
.B(n_810),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_917),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_917),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_917),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_944),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_944),
.Y(n_1095)
);

INVxp33_ASAP7_75t_SL g1096 ( 
.A(n_978),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_944),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_982),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_932),
.B(n_810),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_932),
.B(n_829),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_983),
.Y(n_1101)
);

XNOR2xp5_ASAP7_75t_L g1102 ( 
.A(n_983),
.B(n_870),
.Y(n_1102)
);

XOR2xp5_ASAP7_75t_L g1103 ( 
.A(n_953),
.B(n_868),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_953),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_979),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_979),
.Y(n_1106)
);

XOR2xp5_ASAP7_75t_L g1107 ( 
.A(n_977),
.B(n_869),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_977),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_936),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_936),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_991),
.B(n_869),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_991),
.B(n_869),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1018),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1028),
.B(n_977),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1004),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_986),
.B(n_977),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1046),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1084),
.B(n_902),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1007),
.A2(n_862),
.B1(n_970),
.B2(n_952),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_989),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_992),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1036),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_993),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1084),
.B(n_649),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_1001),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1058),
.Y(n_1126)
);

AND2x4_ASAP7_75t_SL g1127 ( 
.A(n_1067),
.B(n_818),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1050),
.A2(n_970),
.B1(n_952),
.B2(n_658),
.Y(n_1128)
);

AO221x1_ASAP7_75t_L g1129 ( 
.A1(n_1086),
.A2(n_627),
.B1(n_646),
.B2(n_664),
.C(n_708),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_SL g1130 ( 
.A(n_1034),
.B(n_970),
.Y(n_1130)
);

INVx8_ASAP7_75t_L g1131 ( 
.A(n_1108),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1040),
.B(n_674),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1040),
.B(n_675),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_990),
.A2(n_676),
.B1(n_685),
.B2(n_684),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1071),
.B(n_686),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1043),
.A2(n_985),
.B1(n_995),
.B2(n_994),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1100),
.B(n_692),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_998),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1056),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1002),
.A2(n_716),
.B(n_714),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1079),
.A2(n_731),
.B(n_747),
.C(n_724),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1055),
.B(n_999),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_997),
.B(n_820),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1000),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1027),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1016),
.A2(n_552),
.B(n_551),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1024),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1039),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1045),
.B(n_701),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1005),
.B(n_702),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1021),
.B(n_1038),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_987),
.B(n_988),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1029),
.A2(n_703),
.B1(n_709),
.B2(n_707),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1048),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1026),
.B(n_710),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1021),
.B(n_1012),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1012),
.B(n_715),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1036),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1072),
.B(n_720),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1048),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1041),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1091),
.A2(n_725),
.B1(n_729),
.B2(n_723),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1030),
.B(n_736),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1092),
.A2(n_753),
.B1(n_748),
.B2(n_755),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1033),
.Y(n_1165)
);

O2A1O1Ixp5_ASAP7_75t_L g1166 ( 
.A1(n_1093),
.A2(n_1094),
.B(n_1097),
.C(n_1095),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_1099),
.B(n_822),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1031),
.B(n_760),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1034),
.B(n_762),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1035),
.B(n_819),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_1103),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1014),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1037),
.B(n_821),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1042),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_1109),
.B(n_860),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1096),
.B(n_823),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1080),
.B(n_825),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1003),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1081),
.B(n_600),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1082),
.B(n_696),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1085),
.B(n_706),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_1054),
.B(n_1008),
.C(n_1006),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1025),
.B(n_754),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1073),
.A2(n_858),
.B1(n_640),
.B2(n_746),
.Y(n_1184)
);

AND2x6_ASAP7_75t_SL g1185 ( 
.A(n_1009),
.B(n_828),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1078),
.A2(n_740),
.B1(n_633),
.B2(n_557),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1048),
.B(n_860),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1011),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1013),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1098),
.B(n_860),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1101),
.B(n_1016),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1044),
.B(n_555),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1075),
.B(n_1087),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1015),
.B(n_860),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1017),
.B(n_876),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1104),
.B(n_876),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1019),
.A2(n_1022),
.B(n_1020),
.C(n_1110),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1102),
.B(n_876),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1061),
.B(n_1105),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1047),
.B(n_876),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1057),
.A2(n_858),
.B1(n_559),
.B2(n_561),
.Y(n_1201)
);

AND2x6_ASAP7_75t_L g1202 ( 
.A(n_1083),
.B(n_646),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1106),
.B(n_1064),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1077),
.A2(n_562),
.B1(n_563),
.B2(n_558),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1049),
.B(n_566),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1051),
.B(n_569),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1053),
.B(n_571),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1059),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1074),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1107),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1088),
.B(n_0),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1060),
.B(n_579),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1090),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_996),
.A2(n_588),
.B(n_586),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1063),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1065),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1066),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1068),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1070),
.B(n_589),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1089),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1076),
.A2(n_591),
.B1(n_594),
.B2(n_590),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_996),
.B(n_595),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1010),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1023),
.A2(n_603),
.B1(n_605),
.B2(n_602),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1062),
.A2(n_612),
.B1(n_613),
.B2(n_610),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1023),
.B(n_750),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1052),
.A2(n_624),
.B1(n_628),
.B2(n_617),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1052),
.B(n_0),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1032),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1069),
.B(n_629),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1069),
.B(n_634),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_R g1232 ( 
.A(n_1004),
.B(n_639),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_988),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_991),
.B(n_647),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_997),
.B(n_1),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_988),
.B(n_1),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_988),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1007),
.A2(n_648),
.B1(n_659),
.B2(n_656),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_991),
.B(n_660),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_991),
.B(n_661),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_991),
.B(n_663),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1004),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1004),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1084),
.B(n_671),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1084),
.B(n_673),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_991),
.B(n_678),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_989),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_989),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_986),
.B(n_680),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_989),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_991),
.B(n_687),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_989),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_991),
.B(n_690),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_989),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1018),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1007),
.A2(n_694),
.B1(n_704),
.B2(n_693),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_989),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_986),
.A2(n_711),
.B1(n_712),
.B2(n_705),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1018),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1024),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1018),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1018),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_991),
.A2(n_718),
.B(n_717),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_988),
.B(n_2),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1001),
.Y(n_1265)
);

NOR3xp33_ASAP7_75t_L g1266 ( 
.A(n_986),
.B(n_721),
.C(n_719),
.Y(n_1266)
);

O2A1O1Ixp5_ASAP7_75t_L g1267 ( 
.A1(n_986),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_SL g1268 ( 
.A(n_986),
.B(n_735),
.C(n_722),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1018),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1004),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_986),
.B(n_737),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1001),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1007),
.A2(n_743),
.B1(n_744),
.B2(n_739),
.Y(n_1273)
);

INVxp67_ASAP7_75t_L g1274 ( 
.A(n_988),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_986),
.B(n_749),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1048),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_L g1277 ( 
.A(n_986),
.B(n_664),
.C(n_646),
.Y(n_1277)
);

NAND2x1_ASAP7_75t_L g1278 ( 
.A(n_1048),
.B(n_664),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_991),
.B(n_5),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_989),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1024),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_988),
.B(n_6),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1018),
.Y(n_1283)
);

AND2x6_ASAP7_75t_SL g1284 ( 
.A(n_986),
.B(n_7),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1084),
.B(n_7),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_991),
.B(n_8),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_1058),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_SL g1288 ( 
.A1(n_991),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1048),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1033),
.B(n_10),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_991),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1084),
.B(n_13),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_989),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1120),
.Y(n_1294)
);

NOR3xp33_ASAP7_75t_SL g1295 ( 
.A(n_1242),
.B(n_1270),
.C(n_1243),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1121),
.Y(n_1296)
);

OR2x6_ASAP7_75t_L g1297 ( 
.A(n_1131),
.B(n_16),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1123),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1293),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1151),
.B(n_17),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1143),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1138),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1249),
.B(n_19),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1144),
.Y(n_1304)
);

AND2x2_ASAP7_75t_SL g1305 ( 
.A(n_1204),
.B(n_19),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1116),
.A2(n_184),
.B(n_183),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1193),
.B(n_20),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1271),
.B(n_20),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1247),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1115),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1148),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1158),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1248),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1275),
.B(n_21),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1142),
.B(n_22),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1250),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1111),
.B(n_22),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1126),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1232),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1122),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1112),
.B(n_23),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1143),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1260),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1131),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1252),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_SL g1326 ( 
.A(n_1279),
.B(n_23),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1143),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1165),
.B(n_24),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1161),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1254),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1160),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1174),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1257),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1185),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1234),
.B(n_1239),
.Y(n_1335)
);

NOR3xp33_ASAP7_75t_SL g1336 ( 
.A(n_1149),
.B(n_25),
.C(n_26),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1208),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1167),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1280),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1145),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_1156),
.Y(n_1341)
);

BUFx4f_ASAP7_75t_SL g1342 ( 
.A(n_1126),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1167),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1160),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1217),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1287),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1160),
.Y(n_1347)
);

AND3x1_ASAP7_75t_SL g1348 ( 
.A(n_1284),
.B(n_27),
.C(n_28),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1167),
.Y(n_1349)
);

OR2x2_ASAP7_75t_SL g1350 ( 
.A(n_1290),
.B(n_27),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1233),
.B(n_28),
.Y(n_1351)
);

NOR3xp33_ASAP7_75t_SL g1352 ( 
.A(n_1268),
.B(n_29),
.C(n_30),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1281),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1260),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1178),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1131),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1240),
.B(n_29),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1188),
.Y(n_1358)
);

BUFx8_ASAP7_75t_L g1359 ( 
.A(n_1235),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1154),
.Y(n_1360)
);

NOR3xp33_ASAP7_75t_SL g1361 ( 
.A(n_1150),
.B(n_31),
.C(n_32),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1241),
.B(n_32),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1127),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1218),
.Y(n_1364)
);

INVx3_ASAP7_75t_SL g1365 ( 
.A(n_1287),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1189),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1193),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1113),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1235),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1154),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_R g1371 ( 
.A(n_1125),
.B(n_186),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1246),
.B(n_33),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1147),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1117),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1276),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1265),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1192),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1276),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1237),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1182),
.B(n_37),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1155),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1289),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1215),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1172),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1134),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_SL g1386 ( 
.A(n_1162),
.B(n_38),
.C(n_39),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1139),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1171),
.B(n_41),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1289),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_R g1390 ( 
.A(n_1272),
.B(n_1274),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1251),
.B(n_42),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1213),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1253),
.B(n_43),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1137),
.B(n_43),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_SL g1395 ( 
.A(n_1152),
.B(n_44),
.C(n_45),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_R g1396 ( 
.A(n_1176),
.B(n_1286),
.Y(n_1396)
);

INVx5_ASAP7_75t_L g1397 ( 
.A(n_1202),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1255),
.Y(n_1398)
);

CKINVDCx8_ASAP7_75t_R g1399 ( 
.A(n_1159),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1132),
.B(n_45),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1210),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1278),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1220),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1216),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1199),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1259),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1263),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1133),
.B(n_49),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1261),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1266),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1136),
.Y(n_1411)
);

INVxp67_ASAP7_75t_L g1412 ( 
.A(n_1236),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1262),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1124),
.B(n_1169),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1269),
.Y(n_1415)
);

BUFx4f_ASAP7_75t_L g1416 ( 
.A(n_1264),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1283),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1211),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1291),
.B(n_50),
.C(n_51),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1282),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1153),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1114),
.B(n_52),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1177),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1153),
.B(n_54),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1170),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1203),
.B(n_54),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1183),
.B(n_55),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1209),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1223),
.B(n_55),
.Y(n_1429)
);

INVx5_ASAP7_75t_L g1430 ( 
.A(n_1202),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1196),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1209),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1238),
.B(n_1256),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1157),
.B(n_56),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1198),
.B(n_187),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1173),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1168),
.Y(n_1437)
);

NOR3xp33_ASAP7_75t_SL g1438 ( 
.A(n_1164),
.B(n_57),
.C(n_58),
.Y(n_1438)
);

INVx6_ASAP7_75t_L g1439 ( 
.A(n_1228),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1135),
.B(n_1258),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1273),
.B(n_57),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1202),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1163),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1166),
.Y(n_1444)
);

NOR3xp33_ASAP7_75t_SL g1445 ( 
.A(n_1285),
.B(n_58),
.C(n_59),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1197),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1179),
.B(n_59),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1191),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1140),
.B(n_60),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1292),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_1291),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1180),
.B(n_1181),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1225),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1225),
.B(n_60),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1244),
.B(n_61),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1187),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1222),
.B(n_62),
.Y(n_1457)
);

NAND2x2_ASAP7_75t_L g1458 ( 
.A(n_1288),
.B(n_63),
.Y(n_1458)
);

AND2x6_ASAP7_75t_L g1459 ( 
.A(n_1130),
.B(n_188),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1202),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1205),
.Y(n_1461)
);

BUFx8_ASAP7_75t_L g1462 ( 
.A(n_1267),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1201),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1206),
.Y(n_1464)
);

BUFx10_ASAP7_75t_L g1465 ( 
.A(n_1219),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1207),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1226),
.B(n_63),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1212),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_1118),
.Y(n_1469)
);

INVx4_ASAP7_75t_L g1470 ( 
.A(n_1229),
.Y(n_1470)
);

NOR3xp33_ASAP7_75t_SL g1471 ( 
.A(n_1245),
.B(n_65),
.C(n_66),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1194),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1141),
.B(n_65),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1195),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1190),
.Y(n_1475)
);

AND3x1_ASAP7_75t_SL g1476 ( 
.A(n_1129),
.B(n_67),
.C(n_68),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1200),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1214),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1186),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1230),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1231),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1128),
.A2(n_74),
.B1(n_71),
.B2(n_73),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1184),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1221),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1184),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1403),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1342),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1469),
.A2(n_1277),
.B(n_1119),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1444),
.A2(n_1175),
.B(n_1146),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1306),
.A2(n_1227),
.B(n_1224),
.Y(n_1490)
);

OAI22x1_ASAP7_75t_L g1491 ( 
.A1(n_1421),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1320),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1335),
.A2(n_192),
.B(n_191),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1414),
.A2(n_194),
.B(n_193),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1451),
.B(n_75),
.Y(n_1495)
);

AOI221x1_ASAP7_75t_L g1496 ( 
.A1(n_1303),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.C(n_80),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1446),
.A2(n_197),
.B(n_195),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1355),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1358),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1448),
.B(n_76),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1338),
.B(n_78),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1453),
.B(n_79),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1331),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1319),
.B(n_198),
.Y(n_1504)
);

AOI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1457),
.A2(n_200),
.B(n_199),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1314),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1331),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1308),
.A2(n_81),
.B(n_83),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1472),
.A2(n_203),
.B(n_202),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1475),
.A2(n_206),
.B(n_205),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1477),
.A2(n_208),
.B(n_207),
.Y(n_1511)
);

BUFx4f_ASAP7_75t_L g1512 ( 
.A(n_1320),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1359),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1338),
.B(n_83),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1343),
.B(n_86),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1425),
.B(n_86),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1310),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1440),
.A2(n_87),
.B(n_88),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1467),
.A2(n_1321),
.B(n_1317),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1411),
.A2(n_210),
.B(n_209),
.Y(n_1520)
);

O2A1O1Ixp5_ASAP7_75t_L g1521 ( 
.A1(n_1454),
.A2(n_90),
.B(n_87),
.C(n_89),
.Y(n_1521)
);

OA22x2_ASAP7_75t_L g1522 ( 
.A1(n_1388),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1305),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1357),
.A2(n_213),
.B(n_212),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1436),
.B(n_93),
.Y(n_1525)
);

NOR2x1_ASAP7_75t_SL g1526 ( 
.A(n_1397),
.B(n_94),
.Y(n_1526)
);

NOR2x1_ASAP7_75t_L g1527 ( 
.A(n_1323),
.B(n_214),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1362),
.A2(n_216),
.B(n_215),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1442),
.A2(n_222),
.B(n_220),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1372),
.A2(n_224),
.B(n_223),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1381),
.A2(n_96),
.B(n_97),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1300),
.A2(n_96),
.B(n_97),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1365),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1359),
.Y(n_1534)
);

NOR2xp67_ASAP7_75t_SL g1535 ( 
.A(n_1312),
.B(n_98),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1311),
.Y(n_1536)
);

O2A1O1Ixp5_ASAP7_75t_L g1537 ( 
.A1(n_1455),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1474),
.A2(n_226),
.B(n_225),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1391),
.A2(n_1393),
.B(n_1429),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1423),
.B(n_99),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1363),
.B(n_100),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1450),
.A2(n_228),
.B(n_227),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1369),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1437),
.B(n_101),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1400),
.A2(n_1408),
.B(n_1452),
.Y(n_1545)
);

NOR2xp67_ASAP7_75t_L g1546 ( 
.A(n_1318),
.B(n_229),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1396),
.B(n_102),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1353),
.B(n_1341),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1384),
.B(n_1443),
.Y(n_1549)
);

INVx4_ASAP7_75t_L g1550 ( 
.A(n_1331),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1367),
.B(n_546),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1470),
.A2(n_232),
.B(n_230),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1428),
.B(n_234),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1384),
.B(n_103),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1329),
.Y(n_1555)
);

AOI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1422),
.A2(n_236),
.B(n_235),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1466),
.A2(n_240),
.B(n_239),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1427),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1399),
.B(n_104),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1435),
.A2(n_245),
.B(n_243),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_SL g1561 ( 
.A1(n_1407),
.A2(n_106),
.B(n_107),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1295),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1468),
.A2(n_106),
.B(n_108),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1332),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1366),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1343),
.B(n_108),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1344),
.Y(n_1567)
);

NOR4xp25_ASAP7_75t_L g1568 ( 
.A(n_1419),
.B(n_111),
.C(n_109),
.D(n_110),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1416),
.A2(n_249),
.B(n_246),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1349),
.B(n_109),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1390),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1354),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1349),
.B(n_1424),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1449),
.A2(n_115),
.B(n_112),
.C(n_114),
.Y(n_1574)
);

AO31x2_ASAP7_75t_L g1575 ( 
.A1(n_1483),
.A2(n_253),
.A3(n_254),
.B(n_252),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1404),
.B(n_114),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1481),
.B(n_116),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1376),
.B(n_117),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1461),
.B(n_118),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1485),
.B(n_1464),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1294),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1337),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1351),
.Y(n_1583)
);

CKINVDCx6p67_ASAP7_75t_R g1584 ( 
.A(n_1334),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1447),
.A2(n_257),
.B(n_256),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1315),
.A2(n_260),
.B(n_258),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1296),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1298),
.B(n_119),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1299),
.B(n_119),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1394),
.A2(n_262),
.B(n_261),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1388),
.B(n_121),
.Y(n_1591)
);

AO21x1_ASAP7_75t_L g1592 ( 
.A1(n_1449),
.A2(n_122),
.B(n_123),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1301),
.B(n_122),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1302),
.A2(n_264),
.B(n_263),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1392),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1344),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1412),
.A2(n_1433),
.B1(n_1439),
.B2(n_1478),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1397),
.A2(n_269),
.B(n_268),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1380),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1599)
);

AOI221x1_ASAP7_75t_L g1600 ( 
.A1(n_1326),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.C(n_127),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1304),
.B(n_126),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1420),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1354),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1309),
.B(n_129),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1313),
.A2(n_274),
.B(n_273),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1397),
.A2(n_277),
.B(n_275),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1484),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1344),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1482),
.A2(n_130),
.B(n_132),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1316),
.A2(n_280),
.B(n_278),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1441),
.A2(n_132),
.B(n_133),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1325),
.B(n_133),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1330),
.B(n_134),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1301),
.B(n_134),
.Y(n_1614)
);

AOI21x1_ASAP7_75t_SL g1615 ( 
.A1(n_1434),
.A2(n_135),
.B(n_136),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1439),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1460),
.A2(n_285),
.B(n_282),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1333),
.B(n_138),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1339),
.B(n_139),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_L g1620 ( 
.A(n_1438),
.B(n_140),
.C(n_141),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1340),
.B(n_140),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1465),
.B(n_1322),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1479),
.A2(n_142),
.B(n_143),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_SL g1624 ( 
.A1(n_1410),
.A2(n_142),
.B(n_143),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1432),
.A2(n_287),
.B(n_286),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1327),
.B(n_144),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_SL g1627 ( 
.A1(n_1375),
.A2(n_144),
.B(n_145),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1430),
.A2(n_291),
.B(n_289),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1430),
.A2(n_294),
.B(n_292),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1345),
.A2(n_298),
.B(n_296),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1430),
.A2(n_302),
.B(n_300),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1426),
.A2(n_1385),
.B1(n_1380),
.B2(n_1463),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1364),
.A2(n_304),
.B(n_303),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1406),
.A2(n_308),
.B(n_307),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1409),
.A2(n_311),
.B(n_309),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1415),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1480),
.A2(n_314),
.B(n_313),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1368),
.A2(n_316),
.B(n_315),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1383),
.B(n_146),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1307),
.B(n_147),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1307),
.B(n_148),
.Y(n_1641)
);

AO31x2_ASAP7_75t_L g1642 ( 
.A1(n_1374),
.A2(n_1398),
.A3(n_1413),
.B(n_1387),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1417),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1458),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1426),
.B(n_1297),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1473),
.A2(n_1386),
.B(n_1445),
.C(n_1471),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1480),
.A2(n_319),
.B(n_318),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1459),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1346),
.A2(n_324),
.B(n_321),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1480),
.B(n_148),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1405),
.A2(n_328),
.B(n_326),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1377),
.A2(n_149),
.B(n_150),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1379),
.A2(n_335),
.B(n_334),
.Y(n_1653)
);

AO21x1_ASAP7_75t_L g1654 ( 
.A1(n_1382),
.A2(n_150),
.B(n_151),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1373),
.B(n_151),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1297),
.B(n_153),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1395),
.A2(n_154),
.B(n_155),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1462),
.A2(n_341),
.B(n_336),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_SL g1659 ( 
.A(n_1324),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1519),
.A2(n_1460),
.B(n_1347),
.Y(n_1660)
);

AO31x2_ASAP7_75t_L g1661 ( 
.A1(n_1539),
.A2(n_1462),
.A3(n_1476),
.B(n_1459),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1489),
.A2(n_1402),
.B(n_1328),
.Y(n_1662)
);

AO32x2_ASAP7_75t_L g1663 ( 
.A1(n_1597),
.A2(n_1356),
.A3(n_1348),
.B1(n_1350),
.B2(n_1336),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_SL g1664 ( 
.A1(n_1506),
.A2(n_1352),
.B(n_1361),
.C(n_1371),
.Y(n_1664)
);

O2A1O1Ixp33_ASAP7_75t_SL g1665 ( 
.A1(n_1646),
.A2(n_155),
.B(n_156),
.C(n_157),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1523),
.A2(n_1401),
.B1(n_1418),
.B2(n_1456),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1502),
.A2(n_1431),
.B1(n_1456),
.B2(n_1378),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1545),
.A2(n_1347),
.B(n_1360),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1486),
.Y(n_1669)
);

AO31x2_ASAP7_75t_L g1670 ( 
.A1(n_1648),
.A2(n_1402),
.A3(n_1389),
.B(n_1378),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1632),
.A2(n_1431),
.B1(n_1389),
.B2(n_1378),
.Y(n_1671)
);

OAI21x1_ASAP7_75t_SL g1672 ( 
.A1(n_1518),
.A2(n_1389),
.B(n_1370),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1562),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1580),
.B(n_1347),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1652),
.A2(n_1431),
.B(n_1370),
.C(n_1402),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1495),
.A2(n_1370),
.B1(n_158),
.B2(n_159),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1532),
.A2(n_1609),
.B(n_1623),
.Y(n_1677)
);

O2A1O1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1558),
.A2(n_156),
.B(n_159),
.C(n_160),
.Y(n_1678)
);

AO31x2_ASAP7_75t_L g1679 ( 
.A1(n_1648),
.A2(n_427),
.A3(n_544),
.B(n_542),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1584),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1494),
.A2(n_161),
.B(n_163),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1548),
.B(n_161),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1520),
.A2(n_344),
.B(n_343),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1490),
.A2(n_164),
.B(n_165),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1571),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1549),
.B(n_1573),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1493),
.A2(n_166),
.B(n_167),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1552),
.A2(n_168),
.B(n_170),
.Y(n_1688)
);

AND2x2_ASAP7_75t_SL g1689 ( 
.A(n_1568),
.B(n_171),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1498),
.Y(n_1690)
);

AO22x1_ASAP7_75t_L g1691 ( 
.A1(n_1527),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1508),
.A2(n_172),
.B(n_174),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1620),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_1693)
);

BUFx10_ASAP7_75t_L g1694 ( 
.A(n_1659),
.Y(n_1694)
);

O2A1O1Ixp5_ASAP7_75t_SL g1695 ( 
.A1(n_1650),
.A2(n_175),
.B(n_176),
.C(n_177),
.Y(n_1695)
);

O2A1O1Ixp5_ASAP7_75t_SL g1696 ( 
.A1(n_1499),
.A2(n_1581),
.B(n_1587),
.C(n_1565),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1497),
.A2(n_347),
.B(n_345),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1611),
.A2(n_178),
.B(n_179),
.Y(n_1698)
);

AOI221x1_ASAP7_75t_L g1699 ( 
.A1(n_1531),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.C(n_348),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1599),
.A2(n_180),
.B1(n_349),
.B2(n_351),
.Y(n_1700)
);

AO31x2_ASAP7_75t_L g1701 ( 
.A1(n_1636),
.A2(n_352),
.A3(n_354),
.B(n_355),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1586),
.A2(n_357),
.B(n_358),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1499),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1487),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_SL g1705 ( 
.A1(n_1574),
.A2(n_360),
.B(n_361),
.C(n_362),
.Y(n_1705)
);

BUFx4_ASAP7_75t_SL g1706 ( 
.A(n_1595),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1533),
.Y(n_1707)
);

AO21x1_ASAP7_75t_L g1708 ( 
.A1(n_1563),
.A2(n_545),
.B(n_365),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1547),
.A2(n_366),
.B1(n_368),
.B2(n_369),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1572),
.Y(n_1710)
);

OA21x2_ASAP7_75t_L g1711 ( 
.A1(n_1653),
.A2(n_370),
.B(n_371),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1528),
.A2(n_372),
.B(n_373),
.Y(n_1712)
);

CKINVDCx11_ASAP7_75t_R g1713 ( 
.A(n_1492),
.Y(n_1713)
);

AO31x2_ASAP7_75t_L g1714 ( 
.A1(n_1636),
.A2(n_375),
.A3(n_376),
.B(n_377),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1512),
.Y(n_1715)
);

AO21x2_ASAP7_75t_L g1716 ( 
.A1(n_1565),
.A2(n_379),
.B(n_381),
.Y(n_1716)
);

AND2x6_ASAP7_75t_SL g1717 ( 
.A(n_1559),
.B(n_383),
.Y(n_1717)
);

AO21x2_ASAP7_75t_L g1718 ( 
.A1(n_1581),
.A2(n_384),
.B(n_385),
.Y(n_1718)
);

AO31x2_ASAP7_75t_L g1719 ( 
.A1(n_1587),
.A2(n_387),
.A3(n_388),
.B(n_389),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1512),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1542),
.A2(n_392),
.B(n_393),
.Y(n_1721)
);

AO31x2_ASAP7_75t_L g1722 ( 
.A1(n_1643),
.A2(n_395),
.A3(n_396),
.B(n_397),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1533),
.Y(n_1723)
);

O2A1O1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1607),
.A2(n_398),
.B(n_399),
.C(n_401),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1517),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1503),
.Y(n_1726)
);

NAND2x1p5_ASAP7_75t_L g1727 ( 
.A(n_1543),
.B(n_403),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1602),
.Y(n_1728)
);

AO31x2_ASAP7_75t_L g1729 ( 
.A1(n_1592),
.A2(n_405),
.A3(n_406),
.B(n_407),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1536),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1521),
.A2(n_413),
.B(n_414),
.C(n_415),
.Y(n_1731)
);

NOR4xp25_ASAP7_75t_L g1732 ( 
.A(n_1657),
.B(n_416),
.C(n_417),
.D(n_418),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1496),
.A2(n_419),
.B(n_420),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1513),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1516),
.B(n_422),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1491),
.A2(n_424),
.B1(n_425),
.B2(n_428),
.C(n_431),
.Y(n_1736)
);

O2A1O1Ixp5_ASAP7_75t_L g1737 ( 
.A1(n_1537),
.A2(n_432),
.B(n_435),
.C(n_436),
.Y(n_1737)
);

A2O1A1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1579),
.A2(n_438),
.B(n_439),
.C(n_440),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1522),
.A2(n_441),
.B1(n_443),
.B2(n_445),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1555),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1600),
.A2(n_446),
.B(n_447),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1583),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_SL g1743 ( 
.A1(n_1526),
.A2(n_452),
.B(n_453),
.Y(n_1743)
);

AOI221x1_ASAP7_75t_L g1744 ( 
.A1(n_1624),
.A2(n_454),
.B1(n_457),
.B2(n_458),
.C(n_459),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1530),
.A2(n_460),
.B(n_461),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1538),
.A2(n_462),
.B(n_463),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_SL g1747 ( 
.A(n_1622),
.B(n_465),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1590),
.A2(n_467),
.B(n_469),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1564),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1503),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1543),
.Y(n_1751)
);

AOI31xp67_ASAP7_75t_L g1752 ( 
.A1(n_1588),
.A2(n_470),
.A3(n_471),
.B(n_473),
.Y(n_1752)
);

NAND3x1_ASAP7_75t_L g1753 ( 
.A(n_1645),
.B(n_474),
.C(n_475),
.Y(n_1753)
);

BUFx2_ASAP7_75t_R g1754 ( 
.A(n_1641),
.Y(n_1754)
);

INVx4_ASAP7_75t_L g1755 ( 
.A(n_1541),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_SL g1756 ( 
.A1(n_1655),
.A2(n_476),
.B(n_477),
.C(n_478),
.Y(n_1756)
);

AO31x2_ASAP7_75t_L g1757 ( 
.A1(n_1582),
.A2(n_480),
.A3(n_481),
.B(n_482),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1525),
.B(n_539),
.Y(n_1758)
);

OAI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1509),
.A2(n_486),
.B(n_487),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1585),
.A2(n_488),
.B(n_489),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1577),
.B(n_490),
.C(n_492),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1510),
.A2(n_493),
.B(n_494),
.Y(n_1762)
);

INVx5_ASAP7_75t_L g1763 ( 
.A(n_1503),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1659),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1585),
.A2(n_496),
.B(n_500),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1534),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1540),
.A2(n_502),
.B(n_503),
.Y(n_1767)
);

CKINVDCx20_ASAP7_75t_R g1768 ( 
.A(n_1603),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1608),
.B(n_504),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1608),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1608),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1553),
.B(n_505),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1553),
.A2(n_508),
.B(n_509),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1541),
.B(n_510),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1511),
.A2(n_512),
.B(n_513),
.Y(n_1775)
);

CKINVDCx11_ASAP7_75t_R g1776 ( 
.A(n_1550),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1557),
.A2(n_538),
.B(n_516),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1640),
.A2(n_515),
.B1(n_518),
.B2(n_519),
.Y(n_1778)
);

NOR4xp25_ASAP7_75t_L g1779 ( 
.A(n_1616),
.B(n_521),
.C(n_522),
.D(n_523),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1569),
.A2(n_524),
.B(n_525),
.Y(n_1780)
);

AO32x2_ASAP7_75t_L g1781 ( 
.A1(n_1550),
.A2(n_529),
.A3(n_530),
.B1(n_532),
.B2(n_534),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1488),
.A2(n_536),
.B(n_1649),
.Y(n_1782)
);

O2A1O1Ixp33_ASAP7_75t_SL g1783 ( 
.A1(n_1554),
.A2(n_1639),
.B(n_1578),
.C(n_1644),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1488),
.A2(n_1610),
.B(n_1594),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1634),
.A2(n_1635),
.B(n_1605),
.Y(n_1785)
);

AOI21xp33_ASAP7_75t_L g1786 ( 
.A1(n_1500),
.A2(n_1544),
.B(n_1561),
.Y(n_1786)
);

AOI221x1_ASAP7_75t_L g1787 ( 
.A1(n_1644),
.A2(n_1627),
.B1(n_1566),
.B2(n_1647),
.C(n_1637),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1501),
.B(n_1570),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1514),
.B(n_1515),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1598),
.A2(n_1606),
.B(n_1631),
.Y(n_1790)
);

O2A1O1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1576),
.A2(n_1612),
.B(n_1613),
.C(n_1589),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1642),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1601),
.A2(n_1621),
.B1(n_1619),
.B2(n_1618),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1604),
.Y(n_1794)
);

AO32x2_ASAP7_75t_L g1795 ( 
.A1(n_1615),
.A2(n_1654),
.A3(n_1575),
.B1(n_1614),
.B2(n_1593),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1626),
.B(n_1591),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1651),
.A2(n_1560),
.B(n_1546),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1551),
.B(n_1596),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1551),
.B(n_1596),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1677),
.A2(n_1656),
.B1(n_1658),
.B2(n_1504),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1689),
.A2(n_1535),
.B1(n_1507),
.B2(n_1567),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1739),
.A2(n_1567),
.B1(n_1628),
.B2(n_1629),
.Y(n_1802)
);

INVx6_ASAP7_75t_L g1803 ( 
.A(n_1720),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1692),
.A2(n_1698),
.B1(n_1736),
.B2(n_1793),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1670),
.Y(n_1805)
);

BUFx12f_ASAP7_75t_L g1806 ( 
.A(n_1713),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1733),
.A2(n_1633),
.B1(n_1630),
.B2(n_1638),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1700),
.A2(n_1666),
.B1(n_1664),
.B2(n_1676),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1774),
.A2(n_1529),
.B1(n_1625),
.B2(n_1617),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_SL g1810 ( 
.A1(n_1741),
.A2(n_1575),
.B1(n_1505),
.B2(n_1524),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1786),
.A2(n_1556),
.B1(n_1575),
.B2(n_1708),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1685),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1794),
.A2(n_1749),
.B1(n_1740),
.B2(n_1730),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_SL g1814 ( 
.A1(n_1747),
.A2(n_1767),
.B1(n_1772),
.B2(n_1789),
.Y(n_1814)
);

BUFx8_ASAP7_75t_SL g1815 ( 
.A(n_1680),
.Y(n_1815)
);

CKINVDCx6p67_ASAP7_75t_R g1816 ( 
.A(n_1715),
.Y(n_1816)
);

BUFx8_ASAP7_75t_L g1817 ( 
.A(n_1720),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_1776),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1690),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1755),
.A2(n_1691),
.B1(n_1693),
.B2(n_1671),
.Y(n_1820)
);

INVx4_ASAP7_75t_L g1821 ( 
.A(n_1763),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1686),
.B(n_1788),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1703),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1768),
.A2(n_1678),
.B1(n_1682),
.B2(n_1791),
.Y(n_1824)
);

CKINVDCx20_ASAP7_75t_R g1825 ( 
.A(n_1725),
.Y(n_1825)
);

BUFx12f_ASAP7_75t_L g1826 ( 
.A(n_1710),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1726),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1778),
.A2(n_1731),
.B1(n_1681),
.B2(n_1687),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1706),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1728),
.Y(n_1830)
);

INVx6_ASAP7_75t_L g1831 ( 
.A(n_1694),
.Y(n_1831)
);

INVx2_ASAP7_75t_SL g1832 ( 
.A(n_1707),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1667),
.A2(n_1753),
.B1(n_1665),
.B2(n_1783),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1704),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1796),
.A2(n_1761),
.B1(n_1672),
.B2(n_1735),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1758),
.A2(n_1734),
.B1(n_1688),
.B2(n_1709),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1798),
.A2(n_1799),
.B1(n_1674),
.B2(n_1675),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1742),
.A2(n_1738),
.B1(n_1732),
.B2(n_1766),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1792),
.A2(n_1684),
.B1(n_1662),
.B2(n_1718),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1716),
.A2(n_1760),
.B1(n_1765),
.B2(n_1721),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1750),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1795),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1754),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1743),
.A2(n_1797),
.B1(n_1668),
.B2(n_1777),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1795),
.Y(n_1845)
);

BUFx8_ASAP7_75t_L g1846 ( 
.A(n_1663),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1705),
.A2(n_1779),
.B1(n_1764),
.B2(n_1673),
.Y(n_1847)
);

BUFx12f_ASAP7_75t_L g1848 ( 
.A(n_1717),
.Y(n_1848)
);

BUFx12f_ASAP7_75t_L g1849 ( 
.A(n_1723),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1726),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1660),
.A2(n_1727),
.B1(n_1771),
.B2(n_1702),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1712),
.A2(n_1745),
.B1(n_1748),
.B2(n_1769),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1711),
.A2(n_1782),
.B1(n_1770),
.B2(n_1721),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1724),
.A2(n_1751),
.B1(n_1773),
.B2(n_1663),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1697),
.A2(n_1784),
.B1(n_1790),
.B2(n_1699),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1763),
.Y(n_1856)
);

BUFx10_ASAP7_75t_L g1857 ( 
.A(n_1756),
.Y(n_1857)
);

INVx6_ASAP7_75t_L g1858 ( 
.A(n_1696),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1661),
.B(n_1781),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1679),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1787),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1701),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_SL g1863 ( 
.A1(n_1781),
.A2(n_1683),
.B1(n_1746),
.B2(n_1661),
.Y(n_1863)
);

BUFx12f_ASAP7_75t_L g1864 ( 
.A(n_1780),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1719),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1701),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1722),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1759),
.A2(n_1775),
.B1(n_1762),
.B2(n_1785),
.Y(n_1868)
);

INVx6_ASAP7_75t_L g1869 ( 
.A(n_1752),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1714),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1719),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1744),
.A2(n_1695),
.B1(n_1729),
.B2(n_1737),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1757),
.A2(n_1451),
.B1(n_1204),
.B2(n_1305),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1677),
.A2(n_1451),
.B1(n_1303),
.B2(n_1314),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1677),
.A2(n_1451),
.B1(n_1204),
.B2(n_1305),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1669),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1686),
.B(n_1486),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1685),
.Y(n_1878)
);

CKINVDCx11_ASAP7_75t_R g1879 ( 
.A(n_1715),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1706),
.Y(n_1880)
);

INVx4_ASAP7_75t_L g1881 ( 
.A(n_1763),
.Y(n_1881)
);

CKINVDCx11_ASAP7_75t_R g1882 ( 
.A(n_1715),
.Y(n_1882)
);

OAI21xp33_ASAP7_75t_L g1883 ( 
.A1(n_1804),
.A2(n_1874),
.B(n_1808),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1861),
.Y(n_1884)
);

BUFx2_ASAP7_75t_L g1885 ( 
.A(n_1841),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1842),
.B(n_1845),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1805),
.B(n_1859),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1812),
.Y(n_1888)
);

BUFx3_ASAP7_75t_L g1889 ( 
.A(n_1856),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1878),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1819),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1823),
.Y(n_1892)
);

AO31x2_ASAP7_75t_L g1893 ( 
.A1(n_1862),
.A2(n_1866),
.A3(n_1871),
.B(n_1870),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1876),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1822),
.B(n_1861),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1869),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1860),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1867),
.B(n_1805),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1877),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1827),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1827),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1864),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1827),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1834),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1865),
.B(n_1855),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1832),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1858),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1858),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1846),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1846),
.Y(n_1910)
);

OAI21x1_ASAP7_75t_L g1911 ( 
.A1(n_1844),
.A2(n_1839),
.B(n_1853),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1857),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1875),
.A2(n_1838),
.B1(n_1814),
.B2(n_1873),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1868),
.A2(n_1811),
.B(n_1828),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1863),
.B(n_1835),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1837),
.Y(n_1916)
);

AO21x2_ASAP7_75t_L g1917 ( 
.A1(n_1809),
.A2(n_1833),
.B(n_1802),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1857),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1879),
.Y(n_1919)
);

NOR2x1_ASAP7_75t_SL g1920 ( 
.A(n_1854),
.B(n_1881),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1850),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1895),
.B(n_1887),
.Y(n_1922)
);

AO21x2_ASAP7_75t_L g1923 ( 
.A1(n_1908),
.A2(n_1824),
.B(n_1820),
.Y(n_1923)
);

AO21x2_ASAP7_75t_L g1924 ( 
.A1(n_1908),
.A2(n_1847),
.B(n_1810),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1893),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1893),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1896),
.Y(n_1927)
);

AO21x2_ASAP7_75t_L g1928 ( 
.A1(n_1914),
.A2(n_1840),
.B(n_1872),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1895),
.B(n_1830),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1891),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1891),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1885),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1887),
.B(n_1816),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1899),
.B(n_1813),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1894),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1893),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1894),
.Y(n_1937)
);

OA21x2_ASAP7_75t_L g1938 ( 
.A1(n_1914),
.A2(n_1800),
.B(n_1851),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1897),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1886),
.B(n_1843),
.Y(n_1940)
);

BUFx3_ASAP7_75t_L g1941 ( 
.A(n_1889),
.Y(n_1941)
);

OR2x6_ASAP7_75t_L g1942 ( 
.A(n_1898),
.B(n_1806),
.Y(n_1942)
);

INVxp33_ASAP7_75t_L g1943 ( 
.A(n_1921),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1892),
.B(n_1836),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1889),
.Y(n_1945)
);

AO21x2_ASAP7_75t_L g1946 ( 
.A1(n_1911),
.A2(n_1807),
.B(n_1801),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1893),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1887),
.B(n_1831),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1887),
.B(n_1831),
.Y(n_1949)
);

AO21x2_ASAP7_75t_L g1950 ( 
.A1(n_1911),
.A2(n_1852),
.B(n_1848),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1922),
.B(n_1890),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1930),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1932),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1930),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1922),
.B(n_1890),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1942),
.B(n_1884),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1942),
.B(n_1888),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1931),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1944),
.B(n_1885),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1931),
.B(n_1888),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1940),
.B(n_1886),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1935),
.B(n_1892),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1939),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1942),
.B(n_1884),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1924),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1935),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1941),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1937),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1924),
.Y(n_1969)
);

OAI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1929),
.A2(n_1883),
.B(n_1915),
.C(n_1913),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1948),
.B(n_1906),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1952),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1957),
.Y(n_1973)
);

NAND3xp33_ASAP7_75t_L g1974 ( 
.A(n_1965),
.B(n_1883),
.C(n_1915),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1951),
.B(n_1933),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1954),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1955),
.B(n_1957),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1963),
.Y(n_1978)
);

AND2x4_ASAP7_75t_SL g1979 ( 
.A(n_1971),
.B(n_1942),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1958),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1976),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1979),
.B(n_1967),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1972),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1980),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1978),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1977),
.B(n_1933),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1982),
.B(n_1986),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1981),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1982),
.B(n_1973),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1985),
.B(n_1979),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1984),
.B(n_1975),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1983),
.B(n_1970),
.Y(n_1992)
);

INVxp67_ASAP7_75t_SL g1993 ( 
.A(n_1983),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1982),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1981),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1989),
.B(n_1919),
.Y(n_1996)
);

AO221x2_ASAP7_75t_L g1997 ( 
.A1(n_1988),
.A2(n_1995),
.B1(n_1974),
.B2(n_1992),
.C(n_1994),
.Y(n_1997)
);

INVxp33_ASAP7_75t_SL g1998 ( 
.A(n_1989),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1993),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1991),
.B(n_1978),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1991),
.Y(n_2001)
);

OAI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1994),
.A2(n_1969),
.B1(n_1965),
.B2(n_1938),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1994),
.B(n_1972),
.Y(n_2003)
);

OAI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_1990),
.A2(n_1969),
.B1(n_1940),
.B2(n_1938),
.C(n_1916),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1987),
.B(n_1959),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1990),
.B(n_1818),
.Y(n_2006)
);

AOI21xp33_ASAP7_75t_L g2007 ( 
.A1(n_1999),
.A2(n_2002),
.B(n_2003),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1997),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_2001),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1996),
.B(n_1829),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_2006),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1997),
.B(n_1961),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_2005),
.B(n_1880),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_2000),
.B(n_1960),
.Y(n_2014)
);

AOI222xp33_ASAP7_75t_L g2015 ( 
.A1(n_2008),
.A2(n_2004),
.B1(n_1998),
.B2(n_1916),
.C1(n_1925),
.C2(n_1926),
.Y(n_2015)
);

O2A1O1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_2008),
.A2(n_1923),
.B(n_1924),
.C(n_1904),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_2012),
.A2(n_1923),
.B1(n_1924),
.B2(n_1946),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_2011),
.B(n_1826),
.Y(n_2018)
);

OAI21xp33_ASAP7_75t_L g2019 ( 
.A1(n_2017),
.A2(n_2007),
.B(n_2014),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_2018),
.B(n_2009),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_2015),
.B(n_2013),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_2016),
.B(n_2010),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_2020),
.B(n_1815),
.Y(n_2023)
);

AOI211xp5_ASAP7_75t_L g2024 ( 
.A1(n_2019),
.A2(n_1943),
.B(n_1902),
.C(n_1918),
.Y(n_2024)
);

OAI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_2022),
.A2(n_1825),
.B(n_1918),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_2021),
.Y(n_2026)
);

OAI32xp33_ASAP7_75t_L g2027 ( 
.A1(n_2022),
.A2(n_1953),
.A3(n_1884),
.B1(n_1941),
.B2(n_1945),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_2026),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2024),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_2023),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_2025),
.Y(n_2031)
);

INVxp33_ASAP7_75t_SL g2032 ( 
.A(n_2027),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2026),
.Y(n_2033)
);

BUFx4_ASAP7_75t_SL g2034 ( 
.A(n_2023),
.Y(n_2034)
);

BUFx4_ASAP7_75t_SL g2035 ( 
.A(n_2023),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2026),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2026),
.Y(n_2037)
);

NOR3xp33_ASAP7_75t_L g2038 ( 
.A(n_2033),
.B(n_1882),
.C(n_1817),
.Y(n_2038)
);

NOR2x1_ASAP7_75t_L g2039 ( 
.A(n_2028),
.B(n_1923),
.Y(n_2039)
);

INVxp67_ASAP7_75t_L g2040 ( 
.A(n_2037),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2036),
.Y(n_2041)
);

NOR2x1_ASAP7_75t_L g2042 ( 
.A(n_2030),
.B(n_1923),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_2032),
.B(n_1817),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_L g2044 ( 
.A(n_2029),
.B(n_1907),
.C(n_1934),
.Y(n_2044)
);

NOR3x1_ASAP7_75t_L g2045 ( 
.A(n_2035),
.B(n_1849),
.C(n_1962),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2031),
.A2(n_1953),
.B(n_1963),
.Y(n_2046)
);

INVxp67_ASAP7_75t_L g2047 ( 
.A(n_2035),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2047),
.Y(n_2048)
);

NAND3xp33_ASAP7_75t_L g2049 ( 
.A(n_2040),
.B(n_2034),
.C(n_1912),
.Y(n_2049)
);

NOR3xp33_ASAP7_75t_L g2050 ( 
.A(n_2041),
.B(n_2043),
.C(n_2038),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_2046),
.B(n_1803),
.Y(n_2051)
);

AOI222xp33_ASAP7_75t_L g2052 ( 
.A1(n_2039),
.A2(n_1925),
.B1(n_1947),
.B2(n_1936),
.C1(n_1926),
.C2(n_1905),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2044),
.B(n_1946),
.Y(n_2053)
);

NAND4xp25_ASAP7_75t_SL g2054 ( 
.A(n_2045),
.B(n_1948),
.C(n_1949),
.D(n_1968),
.Y(n_2054)
);

NOR3xp33_ASAP7_75t_SL g2055 ( 
.A(n_2042),
.B(n_1803),
.C(n_1966),
.Y(n_2055)
);

A2O1A1Ixp33_ASAP7_75t_L g2056 ( 
.A1(n_2051),
.A2(n_1907),
.B(n_1902),
.C(n_1949),
.Y(n_2056)
);

NOR2x1p5_ASAP7_75t_L g2057 ( 
.A(n_2049),
.B(n_1945),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2048),
.B(n_1946),
.Y(n_2058)
);

BUFx2_ASAP7_75t_L g2059 ( 
.A(n_2055),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_SL g2060 ( 
.A(n_2050),
.B(n_1910),
.C(n_1909),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_2053),
.B(n_1907),
.C(n_1934),
.Y(n_2061)
);

AOI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_2059),
.A2(n_2054),
.B1(n_2052),
.B2(n_1907),
.C(n_1950),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_2058),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_R g2064 ( 
.A(n_2060),
.B(n_1912),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2057),
.B(n_1946),
.Y(n_2065)
);

OAI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_2061),
.A2(n_1942),
.B1(n_1910),
.B2(n_1909),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2063),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_2064),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2065),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_2067),
.Y(n_2070)
);

NOR4xp25_ASAP7_75t_L g2071 ( 
.A(n_2068),
.B(n_2062),
.C(n_2056),
.D(n_2066),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_2070),
.A2(n_2069),
.B1(n_1950),
.B2(n_1902),
.Y(n_2072)
);

OAI22x1_ASAP7_75t_L g2073 ( 
.A1(n_2071),
.A2(n_1964),
.B1(n_1956),
.B2(n_1881),
.Y(n_2073)
);

AO21x2_ASAP7_75t_L g2074 ( 
.A1(n_2073),
.A2(n_1920),
.B(n_1950),
.Y(n_2074)
);

OA22x2_ASAP7_75t_L g2075 ( 
.A1(n_2072),
.A2(n_1964),
.B1(n_1956),
.B2(n_1937),
.Y(n_2075)
);

AOI221x1_ASAP7_75t_L g2076 ( 
.A1(n_2073),
.A2(n_1964),
.B1(n_1956),
.B2(n_1912),
.C(n_1927),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2075),
.B(n_1950),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2074),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2078),
.B(n_2076),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2077),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_2079),
.A2(n_1902),
.B1(n_1928),
.B2(n_1917),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2081),
.A2(n_2080),
.B1(n_1902),
.B2(n_1912),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2081),
.A2(n_1902),
.B1(n_1912),
.B2(n_1941),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2082),
.A2(n_1920),
.B(n_1928),
.Y(n_2084)
);

NOR2xp67_ASAP7_75t_L g2085 ( 
.A(n_2083),
.B(n_1821),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_2085),
.Y(n_2086)
);

AOI221xp5_ASAP7_75t_L g2087 ( 
.A1(n_2086),
.A2(n_2084),
.B1(n_1912),
.B2(n_1945),
.C(n_1889),
.Y(n_2087)
);

AOI211xp5_ASAP7_75t_L g2088 ( 
.A1(n_2087),
.A2(n_1903),
.B(n_1901),
.C(n_1900),
.Y(n_2088)
);


endmodule