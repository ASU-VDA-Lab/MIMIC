module fake_jpeg_5668_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_44),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_8),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_52),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_17),
.B1(n_27),
.B2(n_18),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_51),
.B1(n_17),
.B2(n_18),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_24),
.B1(n_17),
.B2(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_22),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_35),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_21),
.C(n_34),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_52),
.C(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_35),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_47),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_83),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_17),
.B1(n_27),
.B2(n_18),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_94),
.B1(n_99),
.B2(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_26),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_92),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_21),
.C(n_26),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_91),
.C(n_25),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_26),
.C(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_33),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_18),
.B1(n_27),
.B2(n_34),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_20),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_27),
.B(n_28),
.C(n_32),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_98),
.B(n_22),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_49),
.B1(n_58),
.B2(n_65),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_53),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_107),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_114),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_32),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_67),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_119),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_70),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_128),
.B(n_91),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_68),
.C(n_70),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_129),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_70),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_77),
.B(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_26),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_71),
.B1(n_53),
.B2(n_63),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_87),
.B1(n_95),
.B2(n_92),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_94),
.B1(n_76),
.B2(n_95),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_122),
.B1(n_112),
.B2(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_137),
.B(n_139),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_143),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_89),
.C(n_88),
.Y(n_144)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_146),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_151),
.B1(n_107),
.B2(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_113),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_124),
.B1(n_126),
.B2(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_81),
.B1(n_87),
.B2(n_90),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_60),
.B1(n_84),
.B2(n_28),
.Y(n_153)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_158),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_86),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_31),
.B(n_30),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_167),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_166),
.A2(n_196),
.B(n_84),
.Y(n_209)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_113),
.C(n_105),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_178),
.C(n_132),
.Y(n_203)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_175),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_110),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_176),
.Y(n_210)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_151),
.C(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_187),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_193),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_148),
.B1(n_145),
.B2(n_143),
.Y(n_201)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_185),
.Y(n_211)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_161),
.Y(n_191)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_135),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_114),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_212),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_132),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_203),
.C(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_186),
.B1(n_171),
.B2(n_187),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_202),
.B(n_217),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_136),
.B1(n_140),
.B2(n_134),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_214),
.B1(n_220),
.B2(n_172),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_163),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_86),
.C(n_79),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_168),
.C(n_184),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_175),
.A2(n_78),
.B1(n_30),
.B2(n_69),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_26),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_224),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_30),
.B1(n_69),
.B2(n_29),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_165),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_0),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_69),
.C(n_33),
.Y(n_224)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_231),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_244),
.C(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_173),
.B1(n_192),
.B2(n_181),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_243),
.B1(n_248),
.B2(n_222),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_189),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_232),
.A2(n_246),
.B1(n_215),
.B2(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_234),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

FAx1_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_189),
.CI(n_196),
.CON(n_235),
.SN(n_235)
);

XNOR2x1_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

NOR4xp25_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_194),
.C(n_174),
.D(n_195),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_240),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_170),
.C(n_196),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_176),
.B1(n_180),
.B2(n_179),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_177),
.B(n_33),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_177),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_252),
.A2(n_254),
.B(n_228),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_218),
.B(n_221),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_1),
.C(n_2),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_225),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_19),
.Y(n_288)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_265),
.A2(n_268),
.B1(n_270),
.B2(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_207),
.B1(n_210),
.B2(n_217),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_229),
.C(n_244),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_227),
.C(n_226),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_202),
.B1(n_205),
.B2(n_213),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_283),
.C(n_285),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_282),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_248),
.B1(n_235),
.B2(n_19),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_284),
.B1(n_252),
.B2(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_248),
.C(n_29),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_19),
.B1(n_29),
.B2(n_0),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_29),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_19),
.C(n_1),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_288),
.A2(n_253),
.B1(n_259),
.B2(n_260),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_11),
.B(n_3),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_1),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_258),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

AO221x1_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_263),
.B1(n_268),
.B2(n_259),
.C(n_257),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_288),
.Y(n_299)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_1),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_277),
.B1(n_283),
.B2(n_289),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_296),
.B1(n_294),
.B2(n_291),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_285),
.C(n_275),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_307),
.C(n_298),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_9),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_9),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_313),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_295),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_311),
.Y(n_320)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_303),
.A3(n_7),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_6),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_324),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_319),
.B(n_322),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_308),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_320),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_300),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_294),
.C(n_301),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_309),
.B(n_314),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_306),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_327),
.B(n_328),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_305),
.B(n_15),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_330),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_319),
.B(n_15),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_325),
.C(n_15),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_14),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_333),
.C(n_331),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_16),
.Y(n_337)
);


endmodule