module fake_jpeg_7170_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_36),
.B(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_21),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_1),
.B(n_2),
.Y(n_44)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_45),
.B1(n_31),
.B2(n_2),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_48),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_32),
.B1(n_33),
.B2(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_52),
.B1(n_60),
.B2(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_33),
.B1(n_29),
.B2(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_26),
.B1(n_34),
.B2(n_21),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_34),
.B1(n_20),
.B2(n_27),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_71),
.Y(n_81)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_80),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_82),
.B1(n_65),
.B2(n_48),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_41),
.B1(n_38),
.B2(n_46),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_64),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_47),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_66),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_103),
.B1(n_109),
.B2(n_27),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_64),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_71),
.B1(n_68),
.B2(n_59),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_110),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_24),
.B(n_25),
.Y(n_137)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_81),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_66),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_36),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_69),
.CI(n_42),
.CON(n_119),
.SN(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_46),
.B(n_56),
.C(n_30),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_73),
.B(n_20),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_84),
.B(n_88),
.C(n_38),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_137),
.B(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_99),
.B(n_30),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_139),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_78),
.B(n_24),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_56),
.A3(n_77),
.B1(n_83),
.B2(n_35),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_94),
.B1(n_50),
.B2(n_54),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_147),
.B1(n_152),
.B2(n_104),
.Y(n_177)
);

AO21x2_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_58),
.B(n_53),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_42),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_42),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_153),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_42),
.B1(n_40),
.B2(n_35),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_139),
.B(n_129),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_98),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_164),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_106),
.B(n_119),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_162),
.B(n_166),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_161),
.B(n_167),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_112),
.B(n_126),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_168),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_124),
.B(n_114),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_28),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_16),
.C(n_15),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_176),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_150),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_181),
.B1(n_183),
.B2(n_150),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_138),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_122),
.C(n_40),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_142),
.C(n_149),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_1),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_130),
.B(n_137),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_131),
.B1(n_129),
.B2(n_143),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_104),
.B1(n_125),
.B2(n_58),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_141),
.B1(n_134),
.B2(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_40),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_190),
.C(n_191),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_192),
.B(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_201),
.B1(n_183),
.B2(n_181),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_163),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_131),
.C(n_127),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_198),
.Y(n_232)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_127),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_203),
.Y(n_234)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_161),
.C(n_171),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_17),
.B1(n_19),
.B2(n_23),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_172),
.B1(n_164),
.B2(n_170),
.Y(n_219)
);

AOI22x1_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_28),
.B1(n_30),
.B2(n_22),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_40),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_210),
.A2(n_178),
.B1(n_175),
.B2(n_177),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_212),
.A2(n_217),
.B(n_224),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_209),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_214),
.B(n_220),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_160),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_185),
.C(n_191),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_196),
.B(n_192),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_218),
.B(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_205),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_222),
.B(n_229),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_173),
.B(n_179),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_1),
.B(n_2),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_227),
.B(n_24),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_194),
.B1(n_203),
.B2(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_243),
.C(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_190),
.C(n_199),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_247),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_193),
.C(n_35),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_254),
.C(n_257),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_227),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_24),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_28),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_30),
.C(n_23),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_30),
.C(n_19),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

BUFx4f_ASAP7_75t_SL g262 ( 
.A(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_269),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_278),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_238),
.A2(n_223),
.B1(n_225),
.B2(n_236),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_270),
.A2(n_242),
.B1(n_245),
.B2(n_240),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_224),
.B(n_217),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_275),
.B(n_251),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_272),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_245),
.A2(n_212),
.B1(n_214),
.B2(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

OAI321xp33_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_252),
.A3(n_233),
.B1(n_254),
.B2(n_249),
.C(n_215),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_265),
.C(n_243),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_286),
.C(n_287),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_288),
.B(n_290),
.Y(n_297)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_285),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_241),
.C(n_257),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_291),
.Y(n_298)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_233),
.B(n_4),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_275),
.B1(n_267),
.B2(n_277),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_300),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_269),
.B1(n_266),
.B2(n_272),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_299),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_261),
.B1(n_265),
.B2(n_7),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_307),
.B(n_16),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_3),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_284),
.C(n_10),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_283),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_292),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_7),
.B(n_8),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_8),
.B(n_9),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_11),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_286),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_309),
.B(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_9),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_317),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_303),
.B1(n_299),
.B2(n_302),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_10),
.Y(n_317)
);

OAI21x1_ASAP7_75t_SL g319 ( 
.A1(n_312),
.A2(n_298),
.B(n_304),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_326),
.B(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_313),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_298),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.C(n_331),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_325),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_330),
.A2(n_323),
.B(n_12),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_311),
.B(n_12),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_R g334 ( 
.A(n_332),
.B(n_11),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_333),
.B1(n_327),
.B2(n_16),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);


endmodule