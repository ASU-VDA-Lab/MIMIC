module fake_netlist_1_2684_n_1106 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1106);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1106;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_928;
wire n_813;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_1041;
wire n_578;
wire n_926;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_1060;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_1042;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_1043;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_919;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_1104;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g242 ( .A(n_89), .Y(n_242) );
NOR2xp67_ASAP7_75t_L g243 ( .A(n_195), .B(n_46), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_90), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_54), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_42), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_0), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_186), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_182), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_226), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_127), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_58), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_99), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_133), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_4), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_77), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_87), .Y(n_257) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_26), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_158), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_128), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_76), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_97), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_78), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_213), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_136), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_37), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_21), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_63), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_157), .B(n_149), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_144), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_155), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_55), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_209), .Y(n_275) );
CKINVDCx16_ASAP7_75t_R g276 ( .A(n_113), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_221), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_138), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_217), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_159), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_80), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_53), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_126), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_98), .Y(n_284) );
CKINVDCx16_ASAP7_75t_R g285 ( .A(n_119), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_34), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_201), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_66), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_160), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_110), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_139), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_21), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_60), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_183), .Y(n_294) );
INVxp33_ASAP7_75t_L g295 ( .A(n_227), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_70), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_3), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_58), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_142), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_23), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_120), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_5), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_101), .Y(n_303) );
CKINVDCx16_ASAP7_75t_R g304 ( .A(n_241), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_178), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_184), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_75), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_41), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_84), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_220), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_185), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_37), .B(n_69), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_104), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_18), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_85), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_180), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_190), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_73), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_100), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_79), .Y(n_320) );
INVxp33_ASAP7_75t_L g321 ( .A(n_81), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_93), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_35), .Y(n_323) );
NOR2xp67_ASAP7_75t_L g324 ( .A(n_103), .B(n_117), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_123), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_141), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_131), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_173), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_165), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_222), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_210), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_147), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_164), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_109), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_82), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_35), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_74), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_102), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_169), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_56), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_236), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_203), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_86), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_111), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_26), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_166), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_71), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_11), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_42), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_219), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_8), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_24), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_23), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_137), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_235), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_193), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_207), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_12), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_72), .B(n_181), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_170), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_202), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_132), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_204), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_36), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_40), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_148), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_31), .Y(n_367) );
CKINVDCx14_ASAP7_75t_R g368 ( .A(n_41), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_27), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_234), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_43), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_114), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_30), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_368), .Y(n_374) );
INVx6_ASAP7_75t_L g375 ( .A(n_277), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_245), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_295), .B(n_0), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_344), .B(n_1), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_245), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_277), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_296), .B(n_2), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_263), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_370), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
OAI22xp5_ASAP7_75t_SL g386 ( .A1(n_269), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_311), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_340), .B(n_351), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_340), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
AND2x2_ASAP7_75t_SL g391 ( .A(n_327), .B(n_64), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_263), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_311), .A2(n_67), .B(n_65), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_247), .B(n_5), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_368), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_326), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_263), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_336), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_352), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_295), .B(n_7), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_289), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_352), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_276), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_289), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_290), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_326), .Y(n_407) );
NAND2xp33_ASAP7_75t_L g408 ( .A(n_321), .B(n_68), .Y(n_408) );
AND2x6_ASAP7_75t_L g409 ( .A(n_379), .B(n_377), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
OR2x6_ASAP7_75t_L g411 ( .A(n_398), .B(n_371), .Y(n_411) );
BUFx4f_ASAP7_75t_L g412 ( .A(n_391), .Y(n_412) );
INVx5_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_384), .B(n_252), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_379), .B(n_360), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_391), .A2(n_258), .B1(n_306), .B2(n_261), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_398), .B(n_285), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_404), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_377), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_379), .B(n_360), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_391), .B(n_304), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_391), .B(n_256), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_400), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_400), .B(n_256), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_381), .B(n_337), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_381), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_388), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_383), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_387), .A2(n_255), .B1(n_274), .B2(n_268), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_378), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_374), .A2(n_261), .B1(n_318), .B2(n_306), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_406), .Y(n_434) );
INVx4_ASAP7_75t_L g435 ( .A(n_375), .Y(n_435) );
OR2x6_ASAP7_75t_L g436 ( .A(n_386), .B(n_282), .Y(n_436) );
OR2x6_ASAP7_75t_L g437 ( .A(n_386), .B(n_297), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_378), .B(n_242), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_388), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_378), .B(n_244), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_388), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_388), .Y(n_443) );
AND2x6_ASAP7_75t_L g444 ( .A(n_406), .B(n_290), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_388), .B(n_249), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_376), .B(n_337), .Y(n_446) );
INVx4_ASAP7_75t_L g447 ( .A(n_375), .Y(n_447) );
OR2x6_ASAP7_75t_L g448 ( .A(n_382), .B(n_300), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_376), .B(n_248), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_380), .B(n_293), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_433), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_422), .A2(n_382), .B1(n_395), .B2(n_333), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_411), .B(n_394), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_411), .B(n_298), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_411), .B(n_395), .Y(n_455) );
NAND2xp33_ASAP7_75t_L g456 ( .A(n_409), .B(n_264), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_428), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_428), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_423), .B(n_408), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_SL g460 ( .A1(n_449), .A2(n_396), .B(n_407), .C(n_387), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_434), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_424), .B(n_380), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_412), .A2(n_396), .B1(n_407), .B2(n_387), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_439), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_413), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_415), .A2(n_393), .B(n_343), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_414), .B(n_314), .Y(n_467) );
AND2x6_ASAP7_75t_SL g468 ( .A(n_436), .B(n_302), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_413), .B(n_250), .Y(n_469) );
NAND3xp33_ASAP7_75t_SL g470 ( .A(n_432), .B(n_333), .C(n_318), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_439), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_448), .B(n_335), .Y(n_472) );
BUFx4f_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_441), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_409), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_421), .A2(n_341), .B1(n_342), .B2(n_335), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_443), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_442), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_409), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_425), .B(n_389), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_448), .B(n_323), .Y(n_482) );
INVx5_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_413), .B(n_251), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_409), .B(n_387), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_446), .B(n_396), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_412), .A2(n_341), .B1(n_361), .B2(n_342), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_450), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_426), .B(n_396), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_449), .B(n_361), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_415), .B(n_253), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_418), .B(n_292), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_445), .B(n_407), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_420), .B(n_396), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_420), .A2(n_390), .B1(n_399), .B2(n_389), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_438), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_427), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_444), .B(n_390), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_438), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_440), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_444), .B(n_399), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_430), .A2(n_373), .B1(n_345), .B2(n_348), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_435), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_435), .B(n_402), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_447), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_436), .A2(n_349), .B1(n_353), .B2(n_308), .Y(n_510) );
NAND2xp33_ASAP7_75t_SL g511 ( .A(n_447), .B(n_269), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_436), .B(n_402), .Y(n_512) );
BUFx12f_ASAP7_75t_SL g513 ( .A(n_437), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_437), .B(n_403), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_437), .B(n_403), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_429), .A2(n_365), .B1(n_367), .B2(n_358), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_429), .B(n_254), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_429), .B(n_257), .Y(n_518) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_429), .B(n_369), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_513), .Y(n_520) );
BUFx3_ASAP7_75t_L g521 ( .A(n_472), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_479), .B(n_375), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_466), .A2(n_393), .B(n_338), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_473), .A2(n_472), .B1(n_475), .B2(n_452), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_243), .B(n_260), .C(n_259), .Y(n_525) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_501), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_492), .B(n_286), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_453), .B(n_286), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_457), .Y(n_529) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_519), .A2(n_393), .B(n_312), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_478), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_510), .A2(n_364), .B(n_262), .C(n_270), .Y(n_532) );
AO22x1_ASAP7_75t_L g533 ( .A1(n_492), .A2(n_364), .B1(n_265), .B2(n_278), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_475), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_473), .A2(n_375), .B1(n_246), .B2(n_272), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_475), .B(n_266), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_474), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_457), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_511), .Y(n_539) );
BUFx3_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_482), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_454), .Y(n_542) );
INVxp67_ASAP7_75t_L g543 ( .A(n_467), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_512), .A2(n_267), .B(n_275), .C(n_273), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_455), .A2(n_279), .B1(n_281), .B2(n_280), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_480), .B(n_284), .Y(n_547) );
NOR2xp33_ASAP7_75t_R g548 ( .A(n_470), .B(n_283), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_459), .A2(n_393), .B(n_288), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_SL g550 ( .A1(n_462), .A2(n_271), .B(n_359), .C(n_392), .Y(n_550) );
INVx4_ASAP7_75t_L g551 ( .A(n_475), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_488), .A2(n_393), .B(n_291), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_483), .B(n_480), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_506), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_494), .B(n_310), .Y(n_555) );
INVx4_ASAP7_75t_L g556 ( .A(n_483), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_481), .A2(n_294), .B(n_301), .C(n_287), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_465), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_486), .Y(n_560) );
BUFx8_ASAP7_75t_L g561 ( .A(n_455), .Y(n_561) );
AND2x6_ASAP7_75t_L g562 ( .A(n_485), .B(n_303), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_477), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_514), .B(n_305), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_515), .B(n_309), .Y(n_565) );
XOR2xp5_ASAP7_75t_L g566 ( .A(n_489), .B(n_9), .Y(n_566) );
NOR3xp33_ASAP7_75t_SL g567 ( .A(n_462), .B(n_322), .C(n_307), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_476), .A2(n_246), .B1(n_315), .B2(n_313), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_491), .A2(n_317), .B(n_316), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_487), .A2(n_320), .B(n_319), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_460), .A2(n_328), .B(n_329), .C(n_325), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_498), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_458), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_463), .B(n_505), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_463), .A2(n_246), .B1(n_331), .B2(n_330), .Y(n_575) );
BUFx4f_ASAP7_75t_SL g576 ( .A(n_493), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_SL g577 ( .A1(n_460), .A2(n_332), .B(n_339), .C(n_334), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_508), .A2(n_496), .B(n_471), .C(n_464), .Y(n_578) );
BUFx12f_ASAP7_75t_L g579 ( .A(n_468), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_456), .A2(n_246), .B1(n_356), .B2(n_357), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_495), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_469), .A2(n_347), .B(n_346), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_508), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_500), .A2(n_362), .B(n_372), .C(n_350), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_497), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_502), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_465), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_503), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_507), .B(n_354), .Y(n_589) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_509), .B(n_324), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_504), .A2(n_363), .B1(n_366), .B2(n_271), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_499), .B(n_9), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_516), .B(n_359), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_516), .B(n_289), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_469), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_451), .B(n_10), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_484), .Y(n_597) );
INVx4_ASAP7_75t_L g598 ( .A(n_461), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_517), .A2(n_355), .B1(n_299), .B2(n_401), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_518), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_472), .B(n_10), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_490), .A2(n_355), .B(n_299), .C(n_385), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_473), .A2(n_355), .B1(n_397), .B2(n_385), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_475), .B(n_355), .Y(n_604) );
INVx4_ASAP7_75t_L g605 ( .A(n_475), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_466), .A2(n_385), .B(n_383), .Y(n_606) );
OR2x6_ASAP7_75t_L g607 ( .A(n_472), .B(n_12), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_549), .A2(n_385), .B(n_383), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_539), .B(n_383), .Y(n_609) );
AOI221x1_ASAP7_75t_L g610 ( .A1(n_606), .A2(n_405), .B1(n_397), .B2(n_385), .C(n_383), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_574), .B(n_13), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_578), .A2(n_405), .B(n_397), .C(n_383), .Y(n_612) );
NOR2xp33_ASAP7_75t_SL g613 ( .A(n_579), .B(n_383), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_546), .B(n_13), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_586), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_561), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_546), .B(n_14), .Y(n_617) );
INVx4_ASAP7_75t_L g618 ( .A(n_607), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_552), .A2(n_405), .B(n_397), .Y(n_619) );
AO31x2_ASAP7_75t_L g620 ( .A1(n_602), .A2(n_397), .A3(n_405), .B(n_16), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_560), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_523), .A2(n_405), .B(n_397), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_527), .B(n_14), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_588), .Y(n_624) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_530), .A2(n_405), .B(n_397), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_544), .A2(n_405), .B(n_16), .C(n_17), .Y(n_626) );
O2A1O1Ixp5_ASAP7_75t_L g627 ( .A1(n_550), .A2(n_129), .B(n_239), .C(n_237), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_607), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_537), .B(n_15), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_521), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_534), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_571), .A2(n_15), .B(n_17), .C(n_18), .Y(n_632) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_520), .B(n_19), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_554), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_563), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_531), .B(n_19), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_528), .A2(n_20), .B1(n_22), .B2(n_24), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_542), .A2(n_20), .B1(n_22), .B2(n_25), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_573), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_540), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_557), .A2(n_25), .B(n_27), .C(n_28), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_565), .B(n_28), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_524), .B(n_29), .C(n_30), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_583), .A2(n_29), .B(n_32), .C(n_33), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_601), .B(n_32), .Y(n_645) );
BUFx12f_ASAP7_75t_L g646 ( .A(n_561), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_585), .A2(n_33), .B1(n_34), .B2(n_36), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_525), .B(n_38), .C(n_39), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_584), .A2(n_38), .B(n_39), .C(n_40), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_548), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_SL g652 ( .A1(n_596), .A2(n_593), .B(n_553), .C(n_604), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_589), .A2(n_88), .B(n_83), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_541), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_654) );
NAND2xp33_ASAP7_75t_L g655 ( .A(n_526), .B(n_91), .Y(n_655) );
AO31x2_ASAP7_75t_L g656 ( .A1(n_575), .A2(n_47), .A3(n_48), .B(n_49), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_543), .B(n_47), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_532), .A2(n_48), .B1(n_49), .B2(n_50), .C(n_51), .Y(n_658) );
INVx2_ASAP7_75t_SL g659 ( .A(n_576), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_568), .A2(n_50), .B(n_51), .C(n_52), .Y(n_660) );
AO32x2_ASAP7_75t_L g661 ( .A1(n_535), .A2(n_52), .A3(n_53), .B1(n_54), .B2(n_55), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_533), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_572), .A2(n_162), .B(n_233), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_570), .A2(n_56), .B(n_57), .C(n_59), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_569), .A2(n_59), .B(n_60), .C(n_61), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_522), .A2(n_163), .B(n_232), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_598), .B(n_61), .Y(n_667) );
AOI221x1_ASAP7_75t_L g668 ( .A1(n_592), .A2(n_62), .B1(n_92), .B2(n_94), .C(n_95), .Y(n_668) );
OA21x2_ASAP7_75t_L g669 ( .A1(n_582), .A2(n_168), .B(n_96), .Y(n_669) );
CKINVDCx6p67_ASAP7_75t_R g670 ( .A(n_547), .Y(n_670) );
BUFx10_ASAP7_75t_L g671 ( .A(n_547), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_555), .B(n_62), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_566), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_581), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_562), .A2(n_105), .B1(n_106), .B2(n_107), .Y(n_675) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_526), .Y(n_676) );
AO31x2_ASAP7_75t_L g677 ( .A1(n_603), .A2(n_108), .A3(n_112), .B(n_115), .Y(n_677) );
AO31x2_ASAP7_75t_L g678 ( .A1(n_598), .A2(n_116), .A3(n_118), .B(n_121), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_567), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_534), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_600), .A2(n_122), .B(n_124), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_564), .B(n_125), .C(n_130), .Y(n_682) );
BUFx12f_ASAP7_75t_L g683 ( .A(n_595), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_529), .Y(n_684) );
AOI31xp67_ASAP7_75t_L g685 ( .A1(n_599), .A2(n_134), .A3(n_135), .B(n_140), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_562), .A2(n_143), .B1(n_145), .B2(n_146), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_577), .A2(n_150), .B(n_151), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_558), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_580), .A2(n_152), .B1(n_153), .B2(n_154), .Y(n_689) );
INVx3_ASAP7_75t_SL g690 ( .A(n_551), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_551), .B(n_156), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_538), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_562), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_591), .A2(n_161), .B(n_167), .C(n_171), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_597), .A2(n_172), .B(n_174), .C(n_175), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_562), .A2(n_176), .B1(n_177), .B2(n_179), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_590), .A2(n_187), .B(n_188), .C(n_189), .Y(n_697) );
OAI21xp5_ASAP7_75t_L g698 ( .A1(n_594), .A2(n_191), .B(n_192), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_SL g699 ( .A1(n_536), .A2(n_556), .B(n_545), .C(n_526), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_587), .A2(n_196), .B1(n_197), .B2(n_198), .C(n_199), .Y(n_700) );
OR2x6_ASAP7_75t_L g701 ( .A(n_605), .B(n_200), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_587), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_618), .A2(n_605), .B1(n_545), .B2(n_556), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_635), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_621), .Y(n_705) );
OA21x2_ASAP7_75t_L g706 ( .A1(n_622), .A2(n_559), .B(n_545), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_674), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_608), .A2(n_559), .B(n_206), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_639), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_701), .A2(n_559), .B1(n_208), .B2(n_211), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_615), .B(n_205), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_618), .A2(n_212), .B1(n_214), .B2(n_215), .Y(n_712) );
OA21x2_ASAP7_75t_L g713 ( .A1(n_610), .A2(n_216), .B(n_218), .Y(n_713) );
INVxp67_ASAP7_75t_L g714 ( .A(n_657), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_624), .B(n_223), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_634), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_672), .A2(n_224), .B(n_225), .C(n_228), .Y(n_717) );
BUFx3_ASAP7_75t_L g718 ( .A(n_646), .Y(n_718) );
OA21x2_ASAP7_75t_L g719 ( .A1(n_619), .A2(n_229), .B(n_230), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_670), .B(n_231), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_629), .Y(n_721) );
OR2x6_ASAP7_75t_L g722 ( .A(n_701), .B(n_240), .Y(n_722) );
OA21x2_ASAP7_75t_L g723 ( .A1(n_625), .A2(n_612), .B(n_668), .Y(n_723) );
NOR2xp33_ASAP7_75t_SL g724 ( .A(n_662), .B(n_613), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_676), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_636), .Y(n_726) );
AO21x1_ASAP7_75t_L g727 ( .A1(n_667), .A2(n_643), .B(n_687), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_654), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_616), .Y(n_729) );
AO21x2_ASAP7_75t_L g730 ( .A1(n_611), .A2(n_652), .B(n_632), .Y(n_730) );
OAI211xp5_ASAP7_75t_L g731 ( .A1(n_651), .A2(n_637), .B(n_658), .C(n_648), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_645), .B(n_623), .Y(n_732) );
OR2x6_ASAP7_75t_L g733 ( .A(n_659), .B(n_628), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_642), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_630), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_645), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_684), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_692), .Y(n_738) );
AO31x2_ASAP7_75t_L g739 ( .A1(n_626), .A2(n_694), .A3(n_695), .B(n_650), .Y(n_739) );
OR2x6_ASAP7_75t_L g740 ( .A(n_683), .B(n_691), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_614), .B(n_617), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_649), .A2(n_693), .B1(n_691), .B2(n_644), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_671), .B(n_640), .Y(n_743) );
INVx4_ASAP7_75t_SL g744 ( .A(n_690), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_656), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_620), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_679), .A2(n_673), .B1(n_671), .B2(n_638), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_676), .B(n_633), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_647), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_641), .A2(n_665), .B1(n_664), .B2(n_660), .C(n_682), .Y(n_750) );
AND2x6_ASAP7_75t_L g751 ( .A(n_676), .B(n_631), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_631), .B(n_680), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_656), .Y(n_753) );
INVx1_ASAP7_75t_SL g754 ( .A(n_702), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_688), .A2(n_609), .B1(n_689), .B2(n_655), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_653), .A2(n_700), .B1(n_696), .B2(n_675), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_656), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_699), .B(n_666), .Y(n_758) );
BUFx3_ASAP7_75t_L g759 ( .A(n_620), .Y(n_759) );
OR2x2_ASAP7_75t_L g760 ( .A(n_620), .B(n_678), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_669), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_686), .A2(n_698), .B1(n_663), .B2(n_681), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_661), .A2(n_685), .B1(n_678), .B2(n_677), .Y(n_763) );
INVxp67_ASAP7_75t_L g764 ( .A(n_697), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_661), .A2(n_412), .B(n_672), .C(n_641), .Y(n_765) );
OAI21x1_ASAP7_75t_L g766 ( .A1(n_678), .A2(n_677), .B(n_661), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_677), .B(n_674), .Y(n_767) );
OA21x2_ASAP7_75t_L g768 ( .A1(n_622), .A2(n_610), .B(n_619), .Y(n_768) );
OA21x2_ASAP7_75t_L g769 ( .A1(n_622), .A2(n_610), .B(n_619), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_608), .A2(n_606), .B(n_622), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_646), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_646), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_618), .A2(n_455), .B1(n_412), .B2(n_607), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_657), .A2(n_510), .B1(n_532), .B2(n_543), .C(n_455), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_608), .A2(n_606), .B(n_622), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_674), .B(n_419), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_674), .B(n_618), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_635), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_608), .A2(n_606), .B(n_622), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_674), .B(n_419), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_674), .B(n_419), .Y(n_781) );
AND2x4_ASAP7_75t_L g782 ( .A(n_674), .B(n_618), .Y(n_782) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_618), .B(n_472), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_635), .Y(n_784) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_657), .A2(n_510), .B1(n_532), .B2(n_543), .C(n_455), .Y(n_785) );
AOI21xp33_ASAP7_75t_L g786 ( .A1(n_611), .A2(n_550), .B(n_571), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_614), .A2(n_416), .B1(n_472), .B2(n_412), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_627), .A2(n_552), .B(n_611), .Y(n_788) );
AO31x2_ASAP7_75t_L g789 ( .A1(n_612), .A2(n_668), .A3(n_610), .B(n_608), .Y(n_789) );
OA21x2_ASAP7_75t_L g790 ( .A1(n_622), .A2(n_610), .B(n_619), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_608), .A2(n_606), .B(n_622), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_674), .B(n_419), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_670), .B(n_455), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_674), .B(n_537), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_674), .B(n_419), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_676), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_635), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_635), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_670), .B(n_455), .Y(n_799) );
AO21x2_ASAP7_75t_L g800 ( .A1(n_622), .A2(n_619), .B(n_608), .Y(n_800) );
AO31x2_ASAP7_75t_L g801 ( .A1(n_612), .A2(n_668), .A3(n_610), .B(n_608), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_616), .Y(n_802) );
AO21x2_ASAP7_75t_L g803 ( .A1(n_622), .A2(n_619), .B(n_608), .Y(n_803) );
BUFx3_ASAP7_75t_L g804 ( .A(n_751), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_705), .B(n_716), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_746), .Y(n_806) );
INVx3_ASAP7_75t_L g807 ( .A(n_751), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_767), .Y(n_808) );
OA21x2_ASAP7_75t_L g809 ( .A1(n_766), .A2(n_763), .B(n_767), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_707), .Y(n_810) );
OA21x2_ASAP7_75t_L g811 ( .A1(n_745), .A2(n_757), .B(n_753), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_741), .B(n_794), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_788), .A2(n_791), .B(n_779), .Y(n_813) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_744), .Y(n_814) );
AND2x4_ASAP7_75t_L g815 ( .A(n_722), .B(n_740), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_704), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_709), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_778), .Y(n_818) );
AOI33xp33_ASAP7_75t_L g819 ( .A1(n_773), .A2(n_732), .A3(n_747), .B1(n_774), .B2(n_785), .B3(n_784), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_797), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_798), .B(n_722), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_722), .B(n_737), .Y(n_822) );
OA21x2_ASAP7_75t_L g823 ( .A1(n_770), .A2(n_775), .B(n_760), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_759), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_738), .B(n_728), .Y(n_825) );
OR2x6_ASAP7_75t_L g826 ( .A(n_740), .B(n_710), .Y(n_826) );
AND2x4_ASAP7_75t_L g827 ( .A(n_740), .B(n_725), .Y(n_827) );
NOR2xp67_ASAP7_75t_L g828 ( .A(n_726), .B(n_771), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_711), .Y(n_829) );
NAND2x1_ASAP7_75t_L g830 ( .A(n_751), .B(n_706), .Y(n_830) );
INVx3_ASAP7_75t_L g831 ( .A(n_751), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_793), .B(n_799), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_734), .B(n_721), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_741), .B(n_736), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_776), .B(n_780), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_711), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_706), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_752), .B(n_735), .Y(n_838) );
AND2x4_ASAP7_75t_L g839 ( .A(n_725), .B(n_796), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_787), .B(n_796), .Y(n_840) );
BUFx3_ASAP7_75t_L g841 ( .A(n_743), .Y(n_841) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_710), .Y(n_842) );
AO21x2_ASAP7_75t_L g843 ( .A1(n_765), .A2(n_786), .B(n_803), .Y(n_843) );
OAI322xp33_ASAP7_75t_L g844 ( .A1(n_714), .A2(n_787), .A3(n_783), .B1(n_795), .B2(n_792), .C1(n_781), .C2(n_750), .Y(n_844) );
OR2x2_ASAP7_75t_L g845 ( .A(n_749), .B(n_782), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_713), .Y(n_846) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_744), .Y(n_847) );
AO21x2_ASAP7_75t_L g848 ( .A1(n_786), .A2(n_803), .B(n_800), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_777), .A2(n_782), .B1(n_742), .B2(n_733), .Y(n_849) );
BUFx2_ASAP7_75t_L g850 ( .A(n_777), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_715), .Y(n_851) );
OA21x2_ASAP7_75t_L g852 ( .A1(n_727), .A2(n_764), .B(n_758), .Y(n_852) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_733), .Y(n_853) );
AO21x2_ASAP7_75t_L g854 ( .A1(n_800), .A2(n_730), .B(n_742), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_733), .Y(n_855) );
OAI21xp5_ASAP7_75t_L g856 ( .A1(n_731), .A2(n_756), .B(n_755), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_754), .B(n_720), .Y(n_857) );
OR2x6_ASAP7_75t_L g858 ( .A(n_748), .B(n_719), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_729), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_768), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_723), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_703), .B(n_739), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_723), .Y(n_863) );
BUFx3_ASAP7_75t_L g864 ( .A(n_718), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_739), .B(n_769), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_769), .B(n_790), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_802), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_724), .B(n_712), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_772), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_719), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_789), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_789), .Y(n_872) );
INVx3_ASAP7_75t_L g873 ( .A(n_761), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_789), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_717), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_801), .Y(n_876) );
AO21x2_ASAP7_75t_L g877 ( .A1(n_708), .A2(n_801), .B(n_762), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_724), .A2(n_412), .B1(n_607), .B2(n_728), .Y(n_878) );
AO21x2_ASAP7_75t_L g879 ( .A1(n_766), .A2(n_767), .B(n_788), .Y(n_879) );
BUFx3_ASAP7_75t_L g880 ( .A(n_751), .Y(n_880) );
INVx3_ASAP7_75t_L g881 ( .A(n_751), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_741), .B(n_767), .Y(n_882) );
BUFx2_ASAP7_75t_L g883 ( .A(n_722), .Y(n_883) );
OR2x6_ASAP7_75t_L g884 ( .A(n_722), .B(n_740), .Y(n_884) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_744), .Y(n_885) );
INVx3_ASAP7_75t_L g886 ( .A(n_751), .Y(n_886) );
OR2x2_ASAP7_75t_L g887 ( .A(n_882), .B(n_812), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_865), .B(n_816), .Y(n_888) );
OR2x2_ASAP7_75t_L g889 ( .A(n_882), .B(n_812), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_816), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_865), .B(n_817), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_860), .Y(n_892) );
NAND2x1_ASAP7_75t_L g893 ( .A(n_826), .B(n_884), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_884), .A2(n_883), .B1(n_815), .B2(n_821), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_838), .Y(n_895) );
BUFx2_ASAP7_75t_L g896 ( .A(n_883), .Y(n_896) );
INVx5_ASAP7_75t_SL g897 ( .A(n_884), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_818), .B(n_820), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_820), .B(n_834), .Y(n_899) );
INVx5_ASAP7_75t_SL g900 ( .A(n_884), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_834), .B(n_805), .Y(n_901) );
OAI22xp5_ASAP7_75t_SL g902 ( .A1(n_815), .A2(n_847), .B1(n_885), .B2(n_814), .Y(n_902) );
BUFx3_ASAP7_75t_L g903 ( .A(n_864), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_810), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_811), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_833), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_833), .Y(n_907) );
INVx2_ASAP7_75t_SL g908 ( .A(n_804), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_825), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_811), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_825), .B(n_835), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_811), .Y(n_912) );
AND2x4_ASAP7_75t_L g913 ( .A(n_840), .B(n_826), .Y(n_913) );
INVxp67_ASAP7_75t_L g914 ( .A(n_864), .Y(n_914) );
OAI222xp33_ASAP7_75t_L g915 ( .A1(n_826), .A2(n_815), .B1(n_849), .B2(n_878), .C1(n_850), .C2(n_821), .Y(n_915) );
AND2x4_ASAP7_75t_L g916 ( .A(n_826), .B(n_824), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_819), .B(n_850), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_808), .B(n_866), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_822), .B(n_838), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_845), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_808), .B(n_866), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_845), .Y(n_922) );
INVx3_ASAP7_75t_L g923 ( .A(n_830), .Y(n_923) );
INVx3_ASAP7_75t_L g924 ( .A(n_830), .Y(n_924) );
INVx1_ASAP7_75t_SL g925 ( .A(n_867), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_822), .B(n_841), .Y(n_926) );
INVx1_ASAP7_75t_SL g927 ( .A(n_841), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_852), .B(n_874), .Y(n_928) );
OR2x2_ASAP7_75t_L g929 ( .A(n_857), .B(n_824), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_852), .B(n_874), .Y(n_930) );
OR2x2_ASAP7_75t_L g931 ( .A(n_806), .B(n_862), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_832), .B(n_856), .Y(n_932) );
INVxp67_ASAP7_75t_L g933 ( .A(n_859), .Y(n_933) );
OR2x2_ASAP7_75t_SL g934 ( .A(n_853), .B(n_837), .Y(n_934) );
OR2x2_ASAP7_75t_L g935 ( .A(n_871), .B(n_876), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_872), .B(n_876), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_869), .B(n_855), .Y(n_937) );
INVxp67_ASAP7_75t_L g938 ( .A(n_828), .Y(n_938) );
AO21x2_ASAP7_75t_L g939 ( .A1(n_861), .A2(n_863), .B(n_872), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_809), .B(n_823), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_827), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_842), .A2(n_851), .B1(n_836), .B2(n_829), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_809), .B(n_823), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_829), .B(n_823), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_809), .B(n_823), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_888), .B(n_809), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_891), .B(n_843), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_918), .B(n_854), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_935), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_918), .B(n_843), .Y(n_950) );
INVx1_ASAP7_75t_SL g951 ( .A(n_927), .Y(n_951) );
INVxp67_ASAP7_75t_L g952 ( .A(n_896), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_921), .B(n_854), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_921), .B(n_843), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_914), .B(n_827), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_935), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_936), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_929), .B(n_879), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_936), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_928), .B(n_848), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_939), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_929), .B(n_813), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_939), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_930), .B(n_813), .Y(n_964) );
AND2x2_ASAP7_75t_SL g965 ( .A(n_916), .B(n_886), .Y(n_965) );
INVx2_ASAP7_75t_SL g966 ( .A(n_893), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_932), .A2(n_844), .B1(n_851), .B2(n_875), .Y(n_967) );
AND2x2_ASAP7_75t_SL g968 ( .A(n_916), .B(n_886), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_905), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_901), .B(n_873), .Y(n_970) );
INVx2_ASAP7_75t_SL g971 ( .A(n_893), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_917), .A2(n_827), .B1(n_868), .B2(n_804), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_899), .B(n_877), .Y(n_973) );
INVx2_ASAP7_75t_L g974 ( .A(n_892), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_897), .A2(n_807), .B1(n_831), .B2(n_881), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_913), .A2(n_880), .B1(n_831), .B2(n_881), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_905), .Y(n_977) );
AND2x4_ASAP7_75t_L g978 ( .A(n_923), .B(n_858), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_898), .B(n_890), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_903), .B(n_807), .Y(n_980) );
AOI31xp33_ASAP7_75t_L g981 ( .A1(n_894), .A2(n_870), .A3(n_839), .B(n_846), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_910), .Y(n_982) );
NAND2xp5_ASAP7_75t_SL g983 ( .A(n_902), .B(n_807), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_940), .B(n_945), .Y(n_984) );
INVxp67_ASAP7_75t_L g985 ( .A(n_951), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_984), .B(n_944), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_969), .Y(n_987) );
INVxp67_ASAP7_75t_SL g988 ( .A(n_952), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_969), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_977), .Y(n_990) );
BUFx3_ASAP7_75t_L g991 ( .A(n_951), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_984), .B(n_940), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_948), .B(n_945), .Y(n_993) );
AOI21xp33_ASAP7_75t_L g994 ( .A1(n_967), .A2(n_896), .B(n_937), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_949), .B(n_895), .Y(n_995) );
INVx1_ASAP7_75t_SL g996 ( .A(n_970), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_982), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_948), .B(n_943), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_982), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_949), .B(n_907), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_953), .B(n_943), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_956), .B(n_906), .Y(n_1002) );
OR2x2_ASAP7_75t_L g1003 ( .A(n_962), .B(n_944), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_956), .B(n_922), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_953), .B(n_912), .Y(n_1005) );
NOR2xp33_ASAP7_75t_L g1006 ( .A(n_955), .B(n_938), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_957), .B(n_920), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_974), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_962), .B(n_931), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_946), .B(n_910), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_974), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_957), .B(n_909), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_958), .B(n_931), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_959), .B(n_889), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_958), .B(n_889), .Y(n_1015) );
OR2x6_ASAP7_75t_L g1016 ( .A(n_966), .B(n_924), .Y(n_1016) );
INVxp33_ASAP7_75t_L g1017 ( .A(n_980), .Y(n_1017) );
OAI21xp33_ASAP7_75t_L g1018 ( .A1(n_967), .A2(n_903), .B(n_933), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_1017), .B(n_925), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1015), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_986), .Y(n_1021) );
O2A1O1Ixp33_ASAP7_75t_SL g1022 ( .A1(n_994), .A2(n_983), .B(n_966), .C(n_971), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_992), .B(n_964), .Y(n_1023) );
AO21x1_ASAP7_75t_L g1024 ( .A1(n_988), .A2(n_981), .B(n_915), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1015), .Y(n_1025) );
NAND2x1_ASAP7_75t_L g1026 ( .A(n_1016), .B(n_966), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_995), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_987), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1005), .B(n_954), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_992), .B(n_964), .Y(n_1030) );
NAND3xp33_ASAP7_75t_SL g1031 ( .A(n_1018), .B(n_975), .C(n_972), .Y(n_1031) );
INVxp67_ASAP7_75t_L g1032 ( .A(n_991), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1005), .B(n_954), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1008), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1008), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_987), .Y(n_1036) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_986), .B(n_950), .Y(n_1037) );
AOI21xp33_ASAP7_75t_L g1038 ( .A1(n_1018), .A2(n_972), .B(n_911), .Y(n_1038) );
AO21x1_ASAP7_75t_L g1039 ( .A1(n_1006), .A2(n_981), .B(n_975), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_989), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_993), .B(n_960), .Y(n_1041) );
AND2x2_ASAP7_75t_SL g1042 ( .A(n_1003), .B(n_965), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_993), .B(n_959), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_998), .B(n_973), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1011), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_998), .B(n_1001), .Y(n_1046) );
NOR2xp33_ASAP7_75t_L g1047 ( .A(n_985), .B(n_979), .Y(n_1047) );
NAND2x1_ASAP7_75t_L g1048 ( .A(n_1016), .B(n_971), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1021), .Y(n_1049) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_1042), .A2(n_897), .B1(n_900), .B2(n_991), .Y(n_1050) );
INVxp67_ASAP7_75t_L g1051 ( .A(n_1019), .Y(n_1051) );
O2A1O1Ixp33_ASAP7_75t_L g1052 ( .A1(n_1039), .A2(n_1007), .B(n_904), .C(n_1014), .Y(n_1052) );
INVxp67_ASAP7_75t_L g1053 ( .A(n_1028), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1020), .Y(n_1054) );
INVx1_ASAP7_75t_SL g1055 ( .A(n_1027), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1025), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_1046), .B(n_1041), .Y(n_1057) );
O2A1O1Ixp33_ASAP7_75t_L g1058 ( .A1(n_1039), .A2(n_952), .B(n_1004), .C(n_971), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g1059 ( .A1(n_1022), .A2(n_1016), .B(n_965), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1034), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_1038), .A2(n_996), .B1(n_1002), .B2(n_1000), .C(n_1001), .Y(n_1061) );
XOR2xp5_ASAP7_75t_L g1062 ( .A(n_1031), .B(n_887), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1046), .B(n_1010), .Y(n_1063) );
OAI222xp33_ASAP7_75t_L g1064 ( .A1(n_1026), .A2(n_996), .B1(n_1016), .B2(n_1003), .C1(n_1009), .C2(n_1013), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1037), .B(n_1009), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g1066 ( .A(n_1032), .B(n_1047), .Y(n_1066) );
NOR2xp33_ASAP7_75t_L g1067 ( .A(n_1043), .B(n_1012), .Y(n_1067) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_1055), .Y(n_1068) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_1062), .A2(n_1024), .B1(n_1042), .B2(n_1022), .Y(n_1069) );
AOI21xp33_ASAP7_75t_L g1070 ( .A1(n_1058), .A2(n_1024), .B(n_1048), .Y(n_1070) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_1052), .A2(n_1048), .B1(n_1037), .B2(n_976), .C(n_1016), .Y(n_1071) );
AOI21xp5_ASAP7_75t_L g1072 ( .A1(n_1059), .A2(n_965), .B(n_968), .Y(n_1072) );
AOI211xp5_ASAP7_75t_L g1073 ( .A1(n_1064), .A2(n_1013), .B(n_978), .C(n_973), .Y(n_1073) );
INVx1_ASAP7_75t_SL g1074 ( .A(n_1049), .Y(n_1074) );
OAI21xp5_ASAP7_75t_L g1075 ( .A1(n_1050), .A2(n_1023), .B(n_1030), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1065), .Y(n_1076) );
O2A1O1Ixp33_ASAP7_75t_L g1077 ( .A1(n_1051), .A2(n_1044), .B(n_1029), .C(n_1033), .Y(n_1077) );
AOI21xp5_ASAP7_75t_L g1078 ( .A1(n_1050), .A2(n_1061), .B(n_1053), .Y(n_1078) );
INVxp67_ASAP7_75t_L g1079 ( .A(n_1066), .Y(n_1079) );
OAI321xp33_ASAP7_75t_L g1080 ( .A1(n_1069), .A2(n_1051), .A3(n_1053), .B1(n_1057), .B2(n_1056), .C(n_1054), .Y(n_1080) );
O2A1O1Ixp33_ASAP7_75t_L g1081 ( .A1(n_1070), .A2(n_1063), .B(n_1067), .C(n_1060), .Y(n_1081) );
A2O1A1O1Ixp25_ASAP7_75t_L g1082 ( .A1(n_1078), .A2(n_1040), .B(n_1036), .C(n_897), .D(n_900), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1083 ( .A1(n_1071), .A2(n_942), .B1(n_979), .B2(n_950), .C(n_947), .Y(n_1083) );
INVxp67_ASAP7_75t_L g1084 ( .A(n_1068), .Y(n_1084) );
OAI211xp5_ASAP7_75t_SL g1085 ( .A1(n_1079), .A2(n_926), .B(n_919), .C(n_941), .Y(n_1085) );
NAND3xp33_ASAP7_75t_L g1086 ( .A(n_1073), .B(n_963), .C(n_961), .Y(n_1086) );
NAND2xp5_ASAP7_75t_SL g1087 ( .A(n_1072), .B(n_1030), .Y(n_1087) );
NOR3xp33_ASAP7_75t_SL g1088 ( .A(n_1080), .B(n_1087), .C(n_1083), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1084), .Y(n_1089) );
OAI211xp5_ASAP7_75t_L g1090 ( .A1(n_1082), .A2(n_1075), .B(n_1074), .C(n_1077), .Y(n_1090) );
AOI21xp33_ASAP7_75t_L g1091 ( .A1(n_1081), .A2(n_1076), .B(n_908), .Y(n_1091) );
INVxp33_ASAP7_75t_L g1092 ( .A(n_1086), .Y(n_1092) );
NAND4xp75_ASAP7_75t_L g1093 ( .A(n_1088), .B(n_968), .C(n_908), .D(n_960), .Y(n_1093) );
OAI21xp5_ASAP7_75t_L g1094 ( .A1(n_1090), .A2(n_1089), .B(n_1092), .Y(n_1094) );
AOI211xp5_ASAP7_75t_L g1095 ( .A1(n_1092), .A2(n_1085), .B(n_880), .C(n_831), .Y(n_1095) );
OR2x6_ASAP7_75t_L g1096 ( .A(n_1094), .B(n_881), .Y(n_1096) );
OR3x1_ASAP7_75t_L g1097 ( .A(n_1093), .B(n_1091), .C(n_900), .Y(n_1097) );
AOI21xp5_ASAP7_75t_L g1098 ( .A1(n_1095), .A2(n_968), .B(n_963), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1096), .Y(n_1099) );
INVx4_ASAP7_75t_L g1100 ( .A(n_1097), .Y(n_1100) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_1100), .Y(n_1101) );
OAI22xp5_ASAP7_75t_SL g1102 ( .A1(n_1100), .A2(n_1098), .B1(n_934), .B2(n_886), .Y(n_1102) );
XOR2xp5_ASAP7_75t_L g1103 ( .A(n_1101), .B(n_1099), .Y(n_1103) );
AOI222xp33_ASAP7_75t_L g1104 ( .A1(n_1103), .A2(n_1102), .B1(n_900), .B2(n_897), .C1(n_839), .C2(n_999), .Y(n_1104) );
AOI22x1_ASAP7_75t_L g1105 ( .A1(n_1104), .A2(n_1045), .B1(n_1035), .B2(n_1034), .Y(n_1105) );
AOI222xp33_ASAP7_75t_L g1106 ( .A1(n_1105), .A2(n_989), .B1(n_999), .B2(n_997), .C1(n_990), .C2(n_961), .Y(n_1106) );
endmodule