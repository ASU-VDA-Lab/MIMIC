module real_jpeg_6057_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_1),
.A2(n_27),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_1),
.A2(n_46),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_46),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_1),
.A2(n_46),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_2),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_3),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_3),
.A2(n_160),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_3),
.A2(n_160),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_3),
.A2(n_29),
.B1(n_160),
.B2(n_415),
.Y(n_414)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_5),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_5),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_5),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_11),
.A2(n_26),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_11),
.B(n_34),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_11),
.A2(n_26),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_11),
.A2(n_26),
.B1(n_40),
.B2(n_220),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_11),
.A2(n_303),
.B(n_306),
.C(n_310),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_11),
.B(n_123),
.C(n_165),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_11),
.B(n_112),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_11),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_11),
.B(n_128),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_13),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_72),
.B1(n_108),
.B2(n_111),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_13),
.A2(n_72),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_13),
.A2(n_72),
.B1(n_132),
.B2(n_336),
.Y(n_335)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_438),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_56),
.B1(n_60),
.B2(n_433),
.C(n_436),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_22),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_22),
.B(n_56),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_23),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_24),
.B(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_49),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_30),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_31),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_26),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_30),
.Y(n_153)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_34),
.B(n_45),
.Y(n_213)
);

AO22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_42),
.Y(n_34)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_35),
.Y(n_150)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_37),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_38),
.Y(n_221)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_39),
.Y(n_149)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_40),
.Y(n_310)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_41),
.Y(n_157)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_44),
.B(n_69),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_44),
.A2(n_58),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_49),
.B(n_70),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_52),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_54),
.B(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_56),
.A2(n_258),
.B1(n_263),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_56),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_56),
.A2(n_263),
.B(n_269),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B(n_59),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_57),
.A2(n_213),
.B(n_414),
.Y(n_429)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_393),
.B(n_423),
.C(n_426),
.D(n_432),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_385),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_246),
.C(n_292),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_222),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_195),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_65),
.B(n_195),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_144),
.C(n_180),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_66),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_74),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_67),
.B(n_75),
.C(n_114),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_68),
.B(n_213),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_113),
.B1(n_114),
.B2(n_143),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_106),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_77),
.A2(n_112),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_77),
.B(n_217),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_101),
.Y(n_77)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_88),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_81),
.Y(n_305)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_91),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_100),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_96),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_96),
.Y(n_319)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_99),
.Y(n_206)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_99),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_99),
.Y(n_318)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_102),
.B(n_112),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_103),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_106),
.B(n_256),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_107),
.B(n_184),
.Y(n_183)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_112),
.A2(n_184),
.B(n_219),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_113),
.A2(n_114),
.B1(n_418),
.B2(n_419),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_113),
.B(n_400),
.C(n_403),
.Y(n_421)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_114),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_114),
.B(n_419),
.C(n_420),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_135),
.B(n_136),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_115),
.A2(n_203),
.B(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_116),
.B(n_137),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_116),
.B(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_116),
.B(n_315),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_128),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_119),
.Y(n_309)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_128),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_128),
.B(n_315),
.Y(n_330)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_128)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_132),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_135),
.A2(n_232),
.B(n_237),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_135),
.B(n_136),
.Y(n_285)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_144),
.A2(n_145),
.B1(n_180),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_158),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_146),
.B(n_158),
.Y(n_210)
);

AOI32xp33_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.A3(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_149),
.Y(n_280)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_166),
.B(n_170),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_192),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_171),
.A2(n_189),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_171),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_172),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_173),
.Y(n_339)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_187),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_181),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_182),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_182),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_184),
.B(n_219),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_184),
.A2(n_277),
.B(n_404),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_187),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_188),
.B(n_351),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_192),
.B(n_334),
.Y(n_363)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_209),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_198),
.C(n_209),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_201),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_202),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_203),
.B(n_314),
.Y(n_341)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_206),
.Y(n_327)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_212),
.C(n_215),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_222),
.A2(n_388),
.B(n_389),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_245),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_223),
.B(n_245),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_226),
.C(n_238),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_238),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_228),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_230),
.B(n_350),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_237),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_237),
.B(n_330),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_241),
.B(n_429),
.C(n_430),
.Y(n_435)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_243),
.B(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_289),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_247),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_265),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_248),
.B(n_265),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_257),
.C(n_264),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_249),
.B(n_257),
.CI(n_264),
.CON(n_290),
.SN(n_290)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_254),
.C(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_258),
.A2(n_263),
.B1(n_302),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_288),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_274),
.B2(n_275),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_268),
.B(n_274),
.C(n_288),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_284),
.B(n_287),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_276),
.B(n_284),
.Y(n_287)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_287),
.A2(n_397),
.B1(n_398),
.B2(n_405),
.Y(n_396)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_287),
.Y(n_405)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_289),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_290),
.B(n_291),
.Y(n_390)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_290),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_320),
.B(n_384),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_294),
.B(n_297),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.C(n_311),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_298),
.B(n_380),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_301),
.A2(n_311),
.B1(n_312),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_302),
.Y(n_376)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx11_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_378),
.B(n_383),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_368),
.B(n_377),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_345),
.B(n_367),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_331),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_331),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_326),
.B1(n_329),
.B2(n_348),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_340),
.Y(n_331)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_352),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_342),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_343),
.C(n_370),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_354),
.B(n_366),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_349),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_362),
.B(n_365),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_364),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_371),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_374),
.C(n_375),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_382),
.Y(n_383)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_387),
.B(n_390),
.C(n_391),
.D(n_392),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_408),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_407),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_407),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_406),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_405),
.C(n_406),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_399),
.A2(n_400),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_411),
.C(n_421),
.Y(n_431)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_422),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_409),
.B(n_422),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_421),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_416),
.B1(n_417),
.B2(n_420),
.Y(n_412)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_413),
.Y(n_420)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_431),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_431),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_435),
.Y(n_437)
);


endmodule