module fake_jpeg_13809_n_169 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_2),
.B(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_34),
.B(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_1),
.C(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_1),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_53),
.Y(n_61)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_20),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_62),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_67),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_72),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_38),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_23),
.B1(n_53),
.B2(n_3),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_28),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_37),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_93),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_51),
.B1(n_47),
.B2(n_46),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_61),
.B1(n_85),
.B2(n_68),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_105),
.Y(n_112)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_97),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_6),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_11),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_98),
.Y(n_125)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_76),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_75),
.B1(n_83),
.B2(n_77),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_77),
.B1(n_61),
.B2(n_73),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_73),
.C(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_71),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_71),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_107),
.C(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_58),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_105),
.C(n_101),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_90),
.B(n_103),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_100),
.C(n_108),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_80),
.B(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_92),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_136),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_117),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_144),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_137),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_130),
.B(n_133),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_132),
.Y(n_148)
);

AOI21x1_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_139),
.B(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_123),
.C(n_120),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_156),
.Y(n_159)
);

AOI321xp33_ASAP7_75t_L g156 ( 
.A1(n_153),
.A2(n_141),
.A3(n_126),
.B1(n_134),
.B2(n_146),
.C(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_109),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_149),
.B(n_111),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_160),
.A2(n_162),
.B1(n_111),
.B2(n_116),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_124),
.B1(n_58),
.B2(n_84),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_124),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_163),
.B(n_164),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_159),
.A3(n_124),
.B1(n_84),
.B2(n_68),
.C1(n_85),
.C2(n_80),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_80),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_167),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_166),
.Y(n_169)
);


endmodule