module fake_jpeg_14826_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_19),
.A2(n_13),
.B1(n_14),
.B2(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_12),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_12),
.B(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_26),
.Y(n_28)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_18),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_26),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_25),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.C(n_11),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_7),
.B(n_6),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_32),
.B(n_1),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_6),
.B(n_9),
.Y(n_36)
);

NAND4xp25_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_37),
.C(n_0),
.D(n_2),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_5),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_40),
.Y(n_41)
);


endmodule