module fake_jpeg_12414_n_96 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_1),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NAND2x1_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_0),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_29),
.B1(n_42),
.B2(n_38),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_23),
.B1(n_25),
.B2(n_17),
.Y(n_45)
);

OAI31xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_53),
.A3(n_37),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_13),
.B1(n_22),
.B2(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_24),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_35),
.Y(n_51)
);

OA21x2_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_19),
.B(n_25),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_19),
.C(n_21),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_16),
.C(n_13),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_54),
.C(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

CKINVDCx10_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_45),
.B(n_53),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_64),
.B(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_20),
.B1(n_16),
.B2(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_58),
.B1(n_60),
.B2(n_55),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_66),
.B(n_53),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_80),
.B1(n_34),
.B2(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_58),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_8),
.C(n_7),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_56),
.B1(n_57),
.B2(n_63),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_82),
.B(n_85),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_66),
.B(n_68),
.C(n_52),
.D(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_84),
.Y(n_88)
);

OAI322xp33_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_76),
.A3(n_74),
.B1(n_6),
.B2(n_7),
.C1(n_3),
.C2(n_4),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_3),
.B(n_15),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_6),
.B(n_3),
.C(n_15),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_90),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_92),
.C(n_32),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_29),
.Y(n_96)
);


endmodule