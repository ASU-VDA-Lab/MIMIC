module fake_jpeg_2758_n_543 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_45),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_48),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_49),
.Y(n_139)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_52),
.Y(n_160)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_56),
.Y(n_154)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_88),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_34),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_41),
.B(n_13),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_96),
.Y(n_102)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_41),
.B(n_17),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_98),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_112),
.B(n_123),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_69),
.A2(n_29),
.B1(n_15),
.B2(n_30),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_118),
.A2(n_33),
.B1(n_43),
.B2(n_37),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_17),
.B(n_39),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_119),
.A2(n_33),
.B(n_30),
.C(n_15),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_39),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_48),
.B(n_40),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_54),
.B(n_40),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_58),
.B(n_82),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_15),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_40),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_38),
.C(n_43),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_20),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_28),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_65),
.B(n_28),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_74),
.B(n_28),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_164),
.Y(n_233)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_174),
.Y(n_216)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

CKINVDCx12_ASAP7_75t_R g172 ( 
.A(n_100),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_172),
.Y(n_217)
);

BUFx4f_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

OR2x2_ASAP7_75t_SL g177 ( 
.A(n_115),
.B(n_91),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_182),
.Y(n_212)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_109),
.B(n_77),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_119),
.A2(n_78),
.B1(n_79),
.B2(n_47),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_199),
.B1(n_203),
.B2(n_143),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_49),
.B1(n_56),
.B2(n_83),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_189),
.A2(n_210),
.B1(n_143),
.B2(n_100),
.Y(n_239)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_191),
.Y(n_234)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_193),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_102),
.B(n_77),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_101),
.B(n_92),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_200),
.Y(n_220)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_198),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_63),
.B1(n_30),
.B2(n_33),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_25),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_207),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g203 ( 
.A1(n_118),
.A2(n_158),
.B1(n_120),
.B2(n_116),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_206),
.B(n_27),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_27),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_208),
.Y(n_235)
);

BUFx16f_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_133),
.B(n_20),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_209),
.B(n_124),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_124),
.A2(n_29),
.B1(n_143),
.B2(n_161),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_103),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_224),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_117),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_228),
.B1(n_107),
.B2(n_135),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_201),
.B1(n_203),
.B2(n_181),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_177),
.A2(n_147),
.B(n_152),
.C(n_113),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_204),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_238),
.B(n_242),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_243),
.B1(n_196),
.B2(n_207),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_188),
.B(n_141),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_166),
.A2(n_156),
.B1(n_120),
.B2(n_160),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_205),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_246),
.B(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_179),
.C(n_104),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_261),
.C(n_267),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_169),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_248),
.B(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_107),
.B1(n_189),
.B2(n_142),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_250),
.A2(n_263),
.B1(n_271),
.B2(n_221),
.Y(n_292)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_180),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_270),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_155),
.C(n_136),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_219),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_262),
.B(n_268),
.Y(n_298)
);

AO22x1_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_135),
.B1(n_151),
.B2(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_272),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_207),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_220),
.B(n_171),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_194),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_269),
.B(n_213),
.Y(n_304)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_228),
.A2(n_151),
.B1(n_202),
.B2(n_198),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_216),
.B(n_235),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_167),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_222),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_216),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_218),
.B1(n_224),
.B2(n_222),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_276),
.A2(n_265),
.B(n_261),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_227),
.B(n_226),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_296),
.B(n_273),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_282),
.B(n_267),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_235),
.B1(n_214),
.B2(n_234),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_284),
.A2(n_293),
.B1(n_254),
.B2(n_257),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_224),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_288),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_224),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_300),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_224),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_291),
.A2(n_225),
.B(n_130),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_270),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_263),
.A2(n_271),
.B1(n_250),
.B2(n_275),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_232),
.B(n_210),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_238),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_263),
.A2(n_271),
.B1(n_252),
.B2(n_256),
.Y(n_301)
);

AO22x1_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_265),
.B1(n_247),
.B2(n_261),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_213),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_251),
.C(n_253),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_306),
.A2(n_308),
.B(n_319),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_309),
.B(n_327),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_280),
.A2(n_246),
.B1(n_265),
.B2(n_266),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_310),
.A2(n_314),
.B1(n_324),
.B2(n_282),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_248),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_311),
.B(n_312),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_269),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_328),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_280),
.A2(n_246),
.B1(n_214),
.B2(n_247),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_249),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_320),
.Y(n_343)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_317),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_323),
.C(n_326),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_294),
.A2(n_217),
.B(n_229),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_258),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_276),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_231),
.C(n_260),
.Y(n_323)
);

OR2x2_ASAP7_75t_SL g325 ( 
.A(n_294),
.B(n_258),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_332),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_231),
.C(n_255),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_279),
.A2(n_234),
.B(n_117),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_278),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_336),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_225),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_287),
.C(n_276),
.Y(n_352)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_223),
.Y(n_334)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_334),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_245),
.C(n_136),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_319),
.Y(n_360)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_279),
.Y(n_338)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_330),
.B(n_303),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_342),
.B(n_301),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_284),
.Y(n_347)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_347),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_298),
.Y(n_350)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_290),
.Y(n_351)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_357),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_316),
.B(n_290),
.Y(n_353)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_281),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_355),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_281),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_285),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_312),
.B1(n_307),
.B2(n_332),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_313),
.B(n_245),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_364),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_315),
.B(n_236),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_288),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_309),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_366),
.A2(n_306),
.B1(n_307),
.B2(n_327),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_299),
.Y(n_367)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_368),
.A2(n_376),
.B1(n_358),
.B2(n_338),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_318),
.C(n_305),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_372),
.C(n_382),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_314),
.C(n_308),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_366),
.A2(n_315),
.B1(n_327),
.B2(n_309),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_378),
.A2(n_349),
.B1(n_367),
.B2(n_361),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_337),
.A2(n_325),
.B(n_328),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_379),
.A2(n_384),
.B(n_346),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_309),
.C(n_325),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_397),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_345),
.A2(n_322),
.B(n_277),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_333),
.Y(n_388)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_324),
.Y(n_390)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_297),
.Y(n_391)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_299),
.C(n_317),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_394),
.C(n_340),
.Y(n_402)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_393),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_317),
.C(n_296),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_342),
.B(n_322),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_383),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_337),
.A2(n_296),
.B(n_301),
.Y(n_396)
);

XOR2x1_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_341),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_399),
.A2(n_240),
.B1(n_178),
.B2(n_197),
.Y(n_449)
);

XNOR2x1_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_413),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_385),
.C(n_372),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_406),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_340),
.C(n_358),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_SL g436 ( 
.A(n_408),
.B(n_420),
.C(n_421),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_356),
.Y(n_410)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_410),
.Y(n_429)
);

OA22x2_ASAP7_75t_L g412 ( 
.A1(n_373),
.A2(n_346),
.B1(n_345),
.B2(n_362),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_368),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_414),
.A2(n_379),
.B(n_384),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_390),
.A2(n_359),
.B1(n_347),
.B2(n_362),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_415),
.A2(n_422),
.B1(n_424),
.B2(n_244),
.Y(n_447)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_356),
.Y(n_417)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_417),
.Y(n_441)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_369),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_419),
.Y(n_444)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_374),
.A2(n_338),
.B1(n_358),
.B2(n_344),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_374),
.A2(n_344),
.B1(n_350),
.B2(n_355),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_375),
.A2(n_345),
.B1(n_349),
.B2(n_337),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_423),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_375),
.A2(n_293),
.B1(n_292),
.B2(n_361),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_377),
.B(n_336),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_425),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_382),
.C(n_392),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_426),
.B(n_428),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_427),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_380),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_394),
.C(n_387),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_430),
.B(n_433),
.Y(n_467)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_404),
.B(n_376),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_397),
.C(n_395),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_439),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_373),
.C(n_396),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_295),
.C(n_297),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_442),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_295),
.C(n_244),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_399),
.C(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_446),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_423),
.Y(n_445)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_445),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_230),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_415),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_230),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_448),
.B(n_240),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_424),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_403),
.B(n_130),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_221),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_452),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_453),
.A2(n_472),
.B1(n_449),
.B2(n_429),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_412),
.C(n_407),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_457),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_405),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_417),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_460),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_412),
.C(n_408),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_421),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_462),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_414),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_420),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_471),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_410),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_464),
.B(n_465),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_425),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_442),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_470),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_486),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_477),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_467),
.A2(n_434),
.B1(n_445),
.B2(n_435),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_466),
.B(n_468),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_480),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_435),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_456),
.A2(n_438),
.B(n_427),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_483),
.A2(n_185),
.B(n_236),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_456),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_485),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_452),
.C(n_459),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_437),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_436),
.C(n_431),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_144),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_436),
.B1(n_431),
.B2(n_450),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_491),
.B(n_501),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_240),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_494),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_481),
.A2(n_142),
.B(n_191),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_493),
.A2(n_22),
.B(n_13),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_187),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g495 ( 
.A(n_474),
.Y(n_495)
);

AOI322xp5_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_475),
.A3(n_499),
.B1(n_496),
.B2(n_500),
.C1(n_490),
.C2(n_485),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_183),
.C(n_175),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_498),
.B(n_504),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_488),
.A2(n_144),
.B(n_150),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_503),
.A2(n_25),
.B1(n_22),
.B2(n_13),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_153),
.Y(n_504)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_505),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_L g506 ( 
.A1(n_502),
.A2(n_489),
.B(n_484),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_506),
.B(n_510),
.Y(n_525)
);

NOR4xp25_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_12),
.C(n_11),
.D(n_10),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_482),
.A3(n_106),
.B1(n_51),
.B2(n_126),
.C1(n_173),
.C2(n_150),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_511),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_491),
.A2(n_482),
.B1(n_160),
.B2(n_126),
.Y(n_510)
);

AOI322xp5_ASAP7_75t_L g511 ( 
.A1(n_497),
.A2(n_106),
.A3(n_51),
.B1(n_173),
.B2(n_43),
.C1(n_37),
.C2(n_27),
.Y(n_511)
);

AOI322xp5_ASAP7_75t_L g512 ( 
.A1(n_497),
.A2(n_106),
.A3(n_37),
.B1(n_25),
.B2(n_20),
.C1(n_22),
.C2(n_10),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_9),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_515),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_22),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_13),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_518),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_523),
.B(n_527),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_526),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_514),
.A2(n_12),
.B(n_11),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_524),
.A2(n_1),
.B(n_2),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_12),
.C(n_10),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_516),
.Y(n_527)
);

AOI322xp5_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_508),
.C(n_515),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_529),
.A2(n_531),
.B(n_534),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_9),
.C(n_1),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_520),
.C(n_521),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_535),
.A2(n_536),
.B(n_538),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_530),
.A2(n_2),
.B(n_4),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_532),
.A2(n_4),
.B(n_5),
.Y(n_538)
);

AOI322xp5_ASAP7_75t_L g540 ( 
.A1(n_537),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_506),
.C2(n_519),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_539),
.B(n_5),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_541),
.B(n_4),
.Y(n_542)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_542),
.Y(n_543)
);


endmodule