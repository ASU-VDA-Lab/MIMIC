module fake_ariane_1837_n_1013 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1013);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1013;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_586;
wire n_443;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_424;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_764;
wire n_979;
wire n_552;
wire n_348;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_553;
wire n_446;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_557;
wire n_405;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_331;
wire n_559;
wire n_320;
wire n_401;
wire n_485;
wire n_495;
wire n_267;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_839;
wire n_821;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_240;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_671;
wire n_303;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_429;
wire n_654;
wire n_455;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_612;
wire n_333;
wire n_449;
wire n_388;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_543;
wire n_260;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_527;
wire n_290;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_609;
wire n_444;
wire n_355;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_437;
wire n_697;
wire n_274;
wire n_622;
wire n_337;
wire n_967;
wire n_998;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_580;
wire n_358;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_548;
wire n_289;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_144),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_151),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_126),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_124),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_136),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_54),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_127),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_52),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_200),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_140),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_192),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_150),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_43),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_80),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_164),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_167),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_108),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_49),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_4),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_101),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_169),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_196),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_180),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_90),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_219),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_78),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_50),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_25),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_222),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_8),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_162),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_142),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_98),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_165),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_70),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_88),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_135),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_116),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_170),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_48),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_195),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_119),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_107),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_184),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_46),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_208),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_138),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_95),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_139),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_68),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_213),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_25),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_0),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_30),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_223),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_173),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_204),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_134),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_171),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_154),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_121),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_161),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_118),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_218),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_114),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_191),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_156),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_23),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_111),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_112),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_12),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_125),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_174),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_217),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_132),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_207),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_176),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_103),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_104),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_185),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_214),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_105),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_181),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_69),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_34),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_1),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_7),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_172),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_15),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_205),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_190),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_133),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_237),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_120),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_143),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_189),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_33),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_137),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_11),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_84),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_147),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_5),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_210),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_123),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_203),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_221),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_233),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_206),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_38),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_79),
.B(n_21),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_22),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_115),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_55),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_43),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_6),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_183),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_42),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_86),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_145),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_228),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_159),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_177),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_100),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_6),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_62),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_163),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_198),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_41),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_212),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_56),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_226),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_229),
.B(n_122),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_129),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_5),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_141),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_220),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_75),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_26),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_2),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_94),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_40),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_178),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_211),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_10),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_148),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_16),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_47),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_186),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_187),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_197),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_128),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_20),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_35),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_175),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_157),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_182),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_202),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_168),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_21),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_152),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_166),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_285),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g420 ( 
.A1(n_244),
.A2(n_3),
.B(n_4),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_241),
.B(n_7),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_352),
.B(n_296),
.Y(n_422)
);

CKINVDCx6p67_ASAP7_75t_R g423 ( 
.A(n_268),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_254),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_305),
.B(n_9),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_281),
.B(n_10),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_256),
.Y(n_427)
);

BUFx12f_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_399),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_377),
.B(n_13),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

BUFx8_ASAP7_75t_SL g437 ( 
.A(n_408),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_279),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_246),
.B(n_14),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_354),
.B(n_17),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_261),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_261),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_254),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_394),
.B(n_17),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_285),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_254),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_271),
.A2(n_53),
.B(n_51),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_285),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_261),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_285),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_318),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_269),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_251),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_332),
.Y(n_462)
);

OAI22x1_ASAP7_75t_SL g463 ( 
.A1(n_302),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_306),
.B(n_23),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_307),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_308),
.B(n_322),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_326),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_24),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_340),
.B(n_24),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_252),
.Y(n_470)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_274),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_263),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_344),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_266),
.B(n_26),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_357),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_364),
.Y(n_476)
);

BUFx8_ASAP7_75t_SL g477 ( 
.A(n_310),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_369),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_383),
.B(n_27),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_314),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_389),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_270),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_275),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_335),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_291),
.Y(n_486)
);

BUFx8_ASAP7_75t_SL g487 ( 
.A(n_338),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_294),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_297),
.Y(n_489)
);

BUFx8_ASAP7_75t_SL g490 ( 
.A(n_368),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_286),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_298),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_273),
.A2(n_58),
.B(n_57),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_319),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_311),
.A2(n_60),
.B(n_59),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_315),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_324),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_315),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_240),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_315),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_304),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_345),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_397),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_345),
.B(n_61),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_345),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_309),
.A2(n_28),
.B(n_29),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_313),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_330),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_350),
.Y(n_511)
);

BUFx8_ASAP7_75t_SL g512 ( 
.A(n_242),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_360),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_300),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_317),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_323),
.A2(n_30),
.B(n_32),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_334),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_325),
.A2(n_36),
.B(n_37),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_243),
.Y(n_519)
);

BUFx8_ASAP7_75t_L g520 ( 
.A(n_382),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_331),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_398),
.B(n_36),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_333),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_403),
.A2(n_149),
.B(n_239),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_336),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_343),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_245),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_349),
.B(n_37),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_353),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_356),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_365),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_247),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_359),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_477),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_R g536 ( 
.A(n_528),
.B(n_413),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_487),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_490),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_509),
.B(n_334),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_484),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_512),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_437),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_500),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_504),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_467),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_423),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_R g549 ( 
.A(n_427),
.B(n_248),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_519),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_473),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_499),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_R g553 ( 
.A(n_465),
.B(n_249),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_434),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_466),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_428),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_519),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_533),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_R g559 ( 
.A(n_465),
.B(n_412),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_418),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_439),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_417),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_478),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_476),
.B(n_363),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_520),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_520),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_514),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_R g571 ( 
.A(n_422),
.B(n_250),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_R g572 ( 
.A(n_485),
.B(n_411),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_421),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_475),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_481),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_472),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_454),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

INVx8_ASAP7_75t_L g580 ( 
.A(n_422),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_485),
.B(n_280),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_445),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_486),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_495),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_495),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_462),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_447),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_424),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_506),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_417),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_419),
.A2(n_351),
.B1(n_299),
.B2(n_371),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_426),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_450),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_448),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_425),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_491),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_491),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_464),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_R g600 ( 
.A(n_420),
.B(n_507),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_450),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_529),
.B(n_253),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_513),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_R g604 ( 
.A(n_531),
.B(n_255),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_536),
.B(n_431),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_576),
.B(n_529),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_539),
.A2(n_479),
.B1(n_469),
.B2(n_523),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_585),
.B(n_461),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_581),
.Y(n_609)
);

BUFx8_ASAP7_75t_L g610 ( 
.A(n_555),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_586),
.B(n_482),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_579),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_584),
.B(n_449),
.Y(n_613)
);

NOR3xp33_ASAP7_75t_L g614 ( 
.A(n_570),
.B(n_517),
.C(n_468),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_580),
.B(n_449),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_549),
.B(n_474),
.C(n_440),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_574),
.B(n_482),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_557),
.B(n_522),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_579),
.Y(n_619)
);

INVx8_ASAP7_75t_L g620 ( 
.A(n_580),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_560),
.B(n_563),
.C(n_571),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_SL g623 ( 
.A(n_546),
.B(n_420),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_550),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_593),
.A2(n_480),
.B1(n_463),
.B2(n_532),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_588),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_543),
.B(n_483),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_580),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_548),
.B(n_554),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_588),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_604),
.B(n_526),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_566),
.B(n_483),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_560),
.B(n_488),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_563),
.B(n_441),
.C(n_488),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_575),
.B(n_524),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_553),
.B(n_505),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_583),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_602),
.B(n_530),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_577),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

AOI221xp5_ASAP7_75t_L g641 ( 
.A1(n_592),
.A2(n_460),
.B1(n_530),
.B2(n_534),
.C(n_459),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_541),
.B(n_448),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_594),
.B(n_448),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_597),
.B(n_534),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_601),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_582),
.Y(n_646)
);

BUFx5_ASAP7_75t_L g647 ( 
.A(n_595),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_598),
.B(n_470),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_559),
.B(n_526),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_587),
.B(n_489),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_573),
.B(n_492),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_573),
.B(n_502),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_565),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_572),
.B(n_508),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_569),
.B(n_515),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_578),
.B(n_603),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_545),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_540),
.B(n_498),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_590),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_558),
.B(n_521),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_544),
.B(n_527),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_599),
.B(n_430),
.C(n_429),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_562),
.B(n_452),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_591),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_591),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_551),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_567),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_596),
.B(n_510),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_SL g669 ( 
.A(n_651),
.B(n_542),
.C(n_537),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_SL g670 ( 
.A(n_607),
.B(n_564),
.C(n_561),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_637),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_608),
.B(n_511),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_616),
.A2(n_611),
.B1(n_644),
.B2(n_635),
.Y(n_673)
);

BUFx8_ASAP7_75t_L g674 ( 
.A(n_657),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_667),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_628),
.B(n_547),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_645),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_617),
.B(n_511),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_SL g679 ( 
.A(n_652),
.B(n_538),
.C(n_535),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_621),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_609),
.B(n_432),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_620),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_620),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_632),
.B(n_257),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_648),
.B(n_258),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_653),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

INVx5_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_622),
.B(n_556),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_640),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_641),
.A2(n_507),
.B1(n_518),
.B2(n_516),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_639),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_666),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_668),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_646),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_658),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_654),
.B(n_259),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_638),
.B(n_260),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_614),
.A2(n_600),
.B1(n_378),
.B2(n_380),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_615),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_624),
.B(n_446),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_655),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_650),
.B(n_262),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_610),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_627),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_640),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_633),
.B(n_264),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_605),
.A2(n_381),
.B1(n_384),
.B2(n_373),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_612),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_656),
.B(n_265),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_619),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_626),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_630),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_659),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_665),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_660),
.B(n_267),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_634),
.B(n_272),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_642),
.B(n_568),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_664),
.Y(n_719)
);

NOR2x2_ASAP7_75t_L g720 ( 
.A(n_625),
.B(n_456),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_662),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_640),
.Y(n_722)
);

INVx6_ASAP7_75t_L g723 ( 
.A(n_647),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_623),
.A2(n_636),
.B(n_606),
.C(n_613),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_631),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_649),
.B(n_276),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_618),
.B(n_516),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_647),
.B(n_277),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_663),
.Y(n_729)
);

CKINVDCx6p67_ASAP7_75t_R g730 ( 
.A(n_661),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_643),
.A2(n_518),
.B1(n_505),
.B2(n_390),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_647),
.B(n_278),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_647),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_617),
.B(n_400),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_682),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_680),
.Y(n_736)
);

OAI21xp33_ASAP7_75t_SL g737 ( 
.A1(n_734),
.A2(n_493),
.B(n_453),
.Y(n_737)
);

AO32x1_ASAP7_75t_L g738 ( 
.A1(n_727),
.A2(n_443),
.A3(n_435),
.B1(n_436),
.B2(n_444),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_728),
.A2(n_525),
.B(n_496),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_673),
.A2(n_405),
.B(n_410),
.C(n_404),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_682),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_699),
.A2(n_687),
.B(n_705),
.C(n_724),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_702),
.B(n_282),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_696),
.B(n_693),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_703),
.B(n_283),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_670),
.B(n_284),
.Y(n_746)
);

O2A1O1Ixp5_ASAP7_75t_SL g747 ( 
.A1(n_697),
.A2(n_444),
.B(n_443),
.C(n_505),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_682),
.B(n_287),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_698),
.B(n_289),
.C(n_288),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_688),
.B(n_505),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_732),
.A2(n_292),
.B(n_290),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_692),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_672),
.B(n_293),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_709),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_683),
.B(n_295),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_683),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_685),
.B(n_301),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_694),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_671),
.A2(n_367),
.B1(n_312),
.B2(n_316),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_678),
.A2(n_391),
.B1(n_320),
.B2(n_321),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_SL g761 ( 
.A(n_704),
.B(n_303),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_695),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_721),
.B(n_327),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_SL g764 ( 
.A1(n_688),
.A2(n_700),
.B1(n_676),
.B2(n_720),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_686),
.B(n_328),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_714),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_677),
.A2(n_395),
.B(n_337),
.C(n_339),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_708),
.A2(n_402),
.B(n_346),
.C(n_347),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_684),
.A2(n_406),
.B(n_348),
.C(n_355),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_707),
.A2(n_385),
.B1(n_358),
.B2(n_409),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_674),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_711),
.Y(n_772)
);

OAI21xp33_ASAP7_75t_SL g773 ( 
.A1(n_710),
.A2(n_44),
.B(n_45),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_716),
.B(n_712),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_713),
.A2(n_44),
.B(n_45),
.C(n_329),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_681),
.B(n_361),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_690),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_733),
.A2(n_63),
.B(n_65),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_718),
.B(n_452),
.Y(n_779)
);

AOI21xp33_ASAP7_75t_L g780 ( 
.A1(n_717),
.A2(n_375),
.B(n_374),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_690),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_689),
.B(n_471),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_706),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_715),
.A2(n_376),
.B(n_386),
.C(n_388),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_725),
.B(n_392),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_SL g786 ( 
.A(n_726),
.B(n_66),
.C(n_67),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_674),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_723),
.A2(n_591),
.B1(n_503),
.B2(n_501),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_730),
.A2(n_503),
.B1(n_501),
.B2(n_497),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_739),
.A2(n_691),
.B(n_731),
.Y(n_790)
);

OA21x2_ASAP7_75t_L g791 ( 
.A1(n_742),
.A2(n_679),
.B(n_669),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_778),
.A2(n_719),
.B(n_701),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_744),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_766),
.Y(n_794)
);

OAI21xp5_ASAP7_75t_L g795 ( 
.A1(n_774),
.A2(n_722),
.B(n_723),
.Y(n_795)
);

INVx6_ASAP7_75t_L g796 ( 
.A(n_735),
.Y(n_796)
);

BUFx2_ASAP7_75t_R g797 ( 
.A(n_771),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_772),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_758),
.B(n_729),
.Y(n_799)
);

AO21x2_ASAP7_75t_L g800 ( 
.A1(n_740),
.A2(n_729),
.B(n_455),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_735),
.Y(n_801)
);

BUFx2_ASAP7_75t_SL g802 ( 
.A(n_735),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_777),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_777),
.Y(n_804)
);

AO21x2_ASAP7_75t_L g805 ( 
.A1(n_745),
.A2(n_455),
.B(n_451),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_747),
.A2(n_71),
.B(n_72),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_777),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_751),
.A2(n_73),
.B(n_74),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_781),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_787),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_736),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_752),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_775),
.B(n_675),
.C(n_503),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_783),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_762),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_788),
.A2(n_76),
.B(n_77),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_743),
.B(n_675),
.Y(n_817)
);

AO21x2_ASAP7_75t_L g818 ( 
.A1(n_757),
.A2(n_451),
.B(n_457),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_756),
.Y(n_819)
);

AO21x2_ASAP7_75t_L g820 ( 
.A1(n_780),
.A2(n_457),
.B(n_458),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_756),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_754),
.A2(n_81),
.B(n_82),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_763),
.B(n_501),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_750),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_741),
.Y(n_825)
);

OA21x2_ASAP7_75t_L g826 ( 
.A1(n_776),
.A2(n_457),
.B(n_494),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_750),
.B(n_83),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_782),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_737),
.A2(n_85),
.B(n_87),
.Y(n_829)
);

INVx6_ASAP7_75t_SL g830 ( 
.A(n_764),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_755),
.B(n_748),
.Y(n_831)
);

INVx5_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_779),
.A2(n_89),
.B(n_91),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_765),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_784),
.A2(n_749),
.B(n_753),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_794),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_813),
.A2(n_769),
.B1(n_746),
.B2(n_768),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_827),
.B(n_785),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_798),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_829),
.A2(n_738),
.B(n_789),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_793),
.B(n_761),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_829),
.A2(n_770),
.B(n_759),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_834),
.A2(n_760),
.B1(n_767),
.B2(n_786),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_794),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_790),
.A2(n_92),
.B(n_93),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_811),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_797),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_814),
.A2(n_817),
.B1(n_832),
.B2(n_791),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_796),
.Y(n_849)
);

AO21x1_ASAP7_75t_L g850 ( 
.A1(n_795),
.A2(n_822),
.B(n_823),
.Y(n_850)
);

AO21x2_ASAP7_75t_L g851 ( 
.A1(n_820),
.A2(n_818),
.B(n_805),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_812),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_800),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_800),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_815),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_835),
.A2(n_96),
.B(n_97),
.Y(n_856)
);

BUFx4f_ASAP7_75t_SL g857 ( 
.A(n_830),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_810),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_806),
.A2(n_99),
.B(n_102),
.Y(n_859)
);

HB1xp67_ASAP7_75t_SL g860 ( 
.A(n_797),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_799),
.Y(n_861)
);

OAI22xp33_ASAP7_75t_L g862 ( 
.A1(n_791),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_804),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_804),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_803),
.Y(n_865)
);

BUFx2_ASAP7_75t_R g866 ( 
.A(n_802),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_824),
.B(n_113),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_857),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_861),
.B(n_791),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_841),
.B(n_827),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_836),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_844),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_858),
.B(n_831),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_863),
.B(n_864),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_839),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_847),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_846),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_848),
.B(n_828),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_863),
.B(n_807),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_860),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_862),
.A2(n_828),
.B1(n_821),
.B2(n_819),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_SL g882 ( 
.A1(n_837),
.A2(n_822),
.B1(n_820),
.B2(n_816),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_838),
.B(n_833),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_852),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_838),
.B(n_792),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_849),
.B(n_809),
.Y(n_886)
);

AND2x4_ASAP7_75t_SL g887 ( 
.A(n_838),
.B(n_801),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_865),
.B(n_825),
.Y(n_888)
);

OR2x6_ASAP7_75t_L g889 ( 
.A(n_867),
.B(n_816),
.Y(n_889)
);

INVx8_ASAP7_75t_L g890 ( 
.A(n_866),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_843),
.B(n_821),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_855),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_853),
.B(n_826),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_853),
.Y(n_894)
);

NAND2xp33_ASAP7_75t_R g895 ( 
.A(n_856),
.B(n_808),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_875),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_884),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_869),
.B(n_854),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_878),
.B(n_856),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_892),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_878),
.B(n_840),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_885),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_894),
.B(n_850),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_870),
.B(n_845),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_871),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_891),
.B(n_842),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_873),
.B(n_851),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_889),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_872),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_888),
.B(n_851),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_889),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_877),
.Y(n_912)
);

INVxp67_ASAP7_75t_SL g913 ( 
.A(n_893),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_889),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_883),
.B(n_874),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_883),
.B(n_859),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_883),
.B(n_806),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_879),
.B(n_887),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_881),
.B(n_130),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_890),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_890),
.B(n_131),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_886),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_886),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_895),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_896),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_924),
.B(n_882),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_905),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_903),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_915),
.B(n_868),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_905),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_900),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_923),
.B(n_880),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_900),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_923),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_899),
.B(n_876),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_909),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_909),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_897),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_912),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_920),
.B(n_921),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_912),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_903),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_901),
.B(n_146),
.Y(n_943)
);

AND2x2_ASAP7_75t_SL g944 ( 
.A(n_902),
.B(n_153),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_898),
.B(n_913),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_906),
.B(n_155),
.Y(n_946)
);

AND2x4_ASAP7_75t_SL g947 ( 
.A(n_922),
.B(n_158),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_931),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_928),
.B(n_908),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_944),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_945),
.B(n_907),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_928),
.B(n_911),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_942),
.B(n_911),
.Y(n_953)
);

NAND2x1_ASAP7_75t_L g954 ( 
.A(n_934),
.B(n_911),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_942),
.B(n_914),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_926),
.B(n_914),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_933),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_926),
.B(n_914),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_925),
.B(n_906),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_934),
.B(n_917),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_927),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_927),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_935),
.B(n_917),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_938),
.B(n_910),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_932),
.B(n_904),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_943),
.B(n_902),
.Y(n_966)
);

AND2x4_ASAP7_75t_SL g967 ( 
.A(n_929),
.B(n_922),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_930),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_948),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_959),
.B(n_943),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_961),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_957),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_951),
.B(n_929),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_954),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_964),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_950),
.B(n_929),
.Y(n_976)
);

NAND4xp75_ASAP7_75t_SL g977 ( 
.A(n_963),
.B(n_946),
.C(n_919),
.D(n_940),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_968),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_SL g979 ( 
.A1(n_974),
.A2(n_966),
.B1(n_956),
.B2(n_958),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_973),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_975),
.A2(n_952),
.B(n_953),
.Y(n_981)
);

OAI21xp33_ASAP7_75t_L g982 ( 
.A1(n_970),
.A2(n_949),
.B(n_955),
.Y(n_982)
);

OA21x2_ASAP7_75t_L g983 ( 
.A1(n_971),
.A2(n_969),
.B(n_978),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_977),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_972),
.A2(n_960),
.B(n_965),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_976),
.B(n_967),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_983),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_983),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_980),
.Y(n_989)
);

OA21x2_ASAP7_75t_L g990 ( 
.A1(n_981),
.A2(n_962),
.B(n_936),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_922),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_985),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_986),
.B(n_916),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_982),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_979),
.B(n_916),
.Y(n_995)
);

AOI221x1_ASAP7_75t_L g996 ( 
.A1(n_994),
.A2(n_987),
.B1(n_988),
.B2(n_991),
.C(n_992),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_989),
.Y(n_997)
);

OA22x2_ASAP7_75t_L g998 ( 
.A1(n_996),
.A2(n_995),
.B1(n_993),
.B2(n_990),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_997),
.B(n_990),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_998),
.A2(n_947),
.B(n_918),
.Y(n_1000)
);

AOI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_999),
.A2(n_941),
.B1(n_939),
.B2(n_937),
.C(n_936),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_1000),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_1001),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_1002),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_1004),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_1005),
.B(n_1003),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1006),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1007),
.B(n_179),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1008),
.Y(n_1009)
);

XNOR2xp5_ASAP7_75t_L g1010 ( 
.A(n_1009),
.B(n_193),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_SL g1011 ( 
.A1(n_1010),
.A2(n_194),
.B1(n_199),
.B2(n_201),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_1011),
.B(n_209),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_1012),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_1013)
);


endmodule