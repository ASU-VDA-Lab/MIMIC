module fake_jpeg_10839_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_11),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_24),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_26),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_2),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_87),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_103),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_77),
.B1(n_64),
.B2(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_99),
.B1(n_104),
.B2(n_54),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_77),
.B1(n_64),
.B2(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_54),
.B1(n_62),
.B2(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_74),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_54),
.B1(n_63),
.B2(n_61),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_112),
.B1(n_118),
.B2(n_122),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_113),
.B(n_119),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_63),
.B1(n_73),
.B2(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_123),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_60),
.B1(n_62),
.B2(n_70),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_55),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_127),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_2),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_121),
.Y(n_131)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_66),
.B1(n_65),
.B2(n_59),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_78),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_33),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_69),
.B1(n_58),
.B2(n_3),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_69),
.B1(n_58),
.B2(n_31),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_1),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_39),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_1),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_20),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_3),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_142),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_58),
.B1(n_69),
.B2(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_144),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_141),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_119),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_36),
.C(n_38),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_137),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_34),
.B(n_35),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_10),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_12),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_13),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_152),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_156),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_28),
.B(n_32),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_162),
.B1(n_143),
.B2(n_133),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_146),
.C(n_131),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_146),
.B1(n_134),
.B2(n_139),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_172),
.B(n_175),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_133),
.B1(n_42),
.B2(n_44),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_155),
.B(n_156),
.C(n_160),
.D(n_167),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_159),
.B(n_161),
.C(n_164),
.D(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_168),
.B(n_179),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_180),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_171),
.B(n_165),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_169),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_163),
.Y(n_188)
);


endmodule