module fake_jpeg_20167_n_183 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_23),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_21),
.C(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_14),
.B1(n_13),
.B2(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_37),
.B1(n_27),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_14),
.B1(n_13),
.B2(n_16),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_16),
.B1(n_28),
.B2(n_17),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_16),
.B1(n_27),
.B2(n_19),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_22),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_16),
.B1(n_27),
.B2(n_17),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_51),
.Y(n_54)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_39),
.B1(n_52),
.B2(n_32),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_37),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_39),
.C(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_52),
.B1(n_51),
.B2(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_63),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_60),
.C(n_59),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_11),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_88),
.C(n_70),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_60),
.C(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_63),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_94),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_71),
.B(n_61),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_100),
.B(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_92),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_87),
.B(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_105),
.B1(n_91),
.B2(n_87),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_80),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_76),
.B(n_65),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_88),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_70),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_108),
.B1(n_98),
.B2(n_100),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_56),
.B1(n_82),
.B2(n_78),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_74),
.B1(n_82),
.B2(n_77),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_56),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_124),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_66),
.B1(n_41),
.B2(n_64),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_107),
.C(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_129),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_104),
.C(n_106),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_96),
.C(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_134),
.Y(n_145)
);

AOI321xp33_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_64),
.A3(n_102),
.B1(n_19),
.B2(n_12),
.C(n_31),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_20),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_18),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_64),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_24),
.C(n_25),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_37),
.A3(n_36),
.B1(n_53),
.B2(n_33),
.C1(n_49),
.C2(n_52),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_121),
.B1(n_110),
.B2(n_49),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_119),
.C(n_116),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_143),
.C(n_29),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_122),
.C(n_114),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_146),
.B1(n_139),
.B2(n_143),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_126),
.B1(n_136),
.B2(n_133),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_53),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_20),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_151),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_145),
.B(n_147),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_10),
.B(n_9),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_33),
.B1(n_27),
.B2(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_11),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_157),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_11),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_10),
.Y(n_162)
);

XOR2x2_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_15),
.Y(n_163)
);

AO221x1_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_20),
.B1(n_15),
.B2(n_24),
.C(n_29),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_9),
.B(n_8),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_8),
.B(n_1),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_151),
.B1(n_154),
.B2(n_18),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_168),
.B1(n_165),
.B2(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_18),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_170),
.A3(n_171),
.B1(n_1),
.B2(n_2),
.C1(n_3),
.C2(n_4),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_21),
.B1(n_35),
.B2(n_9),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_172),
.A2(n_176),
.B1(n_3),
.B2(n_4),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.C(n_29),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_29),
.A3(n_25),
.B1(n_24),
.B2(n_20),
.C1(n_4),
.C2(n_0),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_20),
.A3(n_24),
.B1(n_25),
.B2(n_5),
.C1(n_2),
.C2(n_3),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_29),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_24),
.C(n_25),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_179),
.B(n_4),
.Y(n_180)
);

OAI321xp33_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_181),
.A3(n_174),
.B1(n_20),
.B2(n_5),
.C(n_25),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_5),
.Y(n_183)
);


endmodule