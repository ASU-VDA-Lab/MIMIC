module real_jpeg_3765_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_1),
.Y(n_139)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_2),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_2),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_134),
.B1(n_161),
.B2(n_221),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_2),
.A2(n_161),
.B1(n_214),
.B2(n_286),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_2),
.A2(n_65),
.B1(n_161),
.B2(n_274),
.Y(n_341)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_3),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_3),
.A2(n_204),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_3),
.B(n_281),
.C(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_3),
.B(n_112),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_3),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_3),
.B(n_60),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_3),
.B(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_5),
.A2(n_63),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_5),
.A2(n_63),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_6),
.Y(n_100)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_7),
.Y(n_241)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_7),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_7),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_7),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_8),
.Y(n_153)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_10),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_75),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_11),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_11),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_11),
.A2(n_123),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_11),
.A2(n_123),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_11),
.A2(n_123),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_58),
.B1(n_129),
.B2(n_134),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_12),
.A2(n_58),
.B1(n_355),
.B2(n_357),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_13),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_13),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_13),
.A2(n_64),
.B1(n_140),
.B2(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_13),
.A2(n_140),
.B1(n_291),
.B2(n_318),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_13),
.A2(n_140),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_14),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_15),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_15),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_15),
.A2(n_89),
.B1(n_230),
.B2(n_234),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_16),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_256),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_255),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_224),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_21),
.B(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_167),
.C(n_184),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_22),
.A2(n_23),
.B1(n_167),
.B2(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_94),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_24),
.B(n_95),
.C(n_166),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_68),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_25),
.B(n_68),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_53),
.B1(n_59),
.B2(n_61),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_26),
.A2(n_265),
.B(n_271),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_26),
.A2(n_59),
.B1(n_297),
.B2(n_341),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_26),
.A2(n_271),
.B(n_341),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_27),
.A2(n_60),
.B1(n_62),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_27),
.A2(n_60),
.B1(n_169),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_27),
.B(n_272),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_40),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_30),
.Y(n_170)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_31),
.Y(n_233)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_31),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_31),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_39),
.Y(n_363)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_40),
.A2(n_297),
.B(n_301),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_46),
.Y(n_212)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_46),
.Y(n_358)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_48),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_48),
.Y(n_320)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_53),
.A2(n_59),
.B(n_301),
.Y(n_404)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_56),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_56),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_56),
.Y(n_300)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_60),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_78),
.B1(n_83),
.B2(n_92),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_73),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_77),
.Y(n_292)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_78),
.B(n_290),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_78),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_78),
.A2(n_92),
.B1(n_211),
.B2(n_354),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_79),
.Y(n_322)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_80),
.Y(n_177)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_81),
.Y(n_293)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_84),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_88),
.Y(n_311)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_88),
.Y(n_356)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_90),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_136),
.B1(n_165),
.B2(n_166),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_95),
.Y(n_165)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_112),
.B1(n_120),
.B2(n_127),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_96),
.A2(n_219),
.B(n_222),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_96),
.A2(n_222),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_96),
.B(n_120),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_97),
.A2(n_128),
.B1(n_223),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_97),
.A2(n_220),
.B1(n_223),
.B2(n_378),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_112),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B1(n_106),
.B2(n_109),
.Y(n_98)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_99),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_104),
.Y(n_196)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_104),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_105),
.Y(n_350)
);

AO22x2_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_112)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_108),
.Y(n_365)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_110),
.Y(n_252)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_121),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_124),
.Y(n_379)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_125),
.Y(n_380)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_133),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g360 ( 
.A1(n_134),
.A2(n_347),
.A3(n_361),
.B1(n_364),
.B2(n_366),
.Y(n_360)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_143),
.B1(n_159),
.B2(n_163),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_163),
.B(n_187),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_196),
.A3(n_197),
.B1(n_199),
.B2(n_203),
.Y(n_195)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_143),
.A2(n_159),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_144),
.A2(n_399),
.B(n_401),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_147),
.Y(n_400)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_163),
.B(n_204),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_164),
.B(n_188),
.Y(n_254)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_167),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_168),
.B(n_174),
.Y(n_244)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_172),
.B(n_367),
.Y(n_366)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_173),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_210),
.B1(n_216),
.B2(n_217),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_175),
.A2(n_178),
.B(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_175),
.A2(n_285),
.B(n_288),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_175),
.A2(n_204),
.B(n_288),
.Y(n_314)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_176),
.Y(n_330)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_184),
.B(n_419),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_194),
.C(n_218),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_185),
.A2(n_186),
.B1(n_218),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_194),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_208),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_195),
.A2(n_208),
.B1(n_209),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_195),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g399 ( 
.A1(n_203),
.A2(n_204),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g344 ( 
.A1(n_204),
.A2(n_345),
.B(n_346),
.Y(n_344)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_218),
.Y(n_414)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_223),
.A2(n_378),
.B(n_381),
.Y(n_377)
);

BUFx24_ASAP7_75t_SL g430 ( 
.A(n_224),
.Y(n_430)
);

FAx1_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.CI(n_243),
.CON(n_224),
.SN(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_238),
.B2(n_242),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_254),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_407),
.B(n_426),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_387),
.B(n_406),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_369),
.B(n_386),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_335),
.B(n_368),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_304),
.B(n_334),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_283),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_263),
.B(n_283),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_275),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_264),
.A2(n_275),
.B1(n_276),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_294),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_284),
.B(n_295),
.C(n_303),
.Y(n_336)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_302),
.B2(n_303),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_326),
.B(n_333),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_315),
.B(n_325),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_314),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_312),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_324),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_324),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_321),
.B(n_323),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_323),
.A2(n_353),
.B(n_359),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_331),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_337),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_351),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_342),
.C(n_351),
.Y(n_370)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx6_ASAP7_75t_SL g349 ( 
.A(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_360),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_360),
.Y(n_375)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx5_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_370),
.B(n_371),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_376),
.B2(n_385),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_375),
.C(n_385),
.Y(n_388)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_382),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_383),
.C(n_384),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_388),
.B(n_389),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_396),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.Y(n_390)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_391),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_393),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_394),
.C(n_396),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_402),
.B2(n_405),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_403),
.C(n_404),
.Y(n_417)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_402),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_421),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_410),
.A2(n_427),
.B(n_428),
.Y(n_426)
);

NOR2x1_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_418),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_418),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.C(n_417),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_416),
.B1(n_417),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_417),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_423),
.Y(n_427)
);


endmodule