module fake_jpeg_32160_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_19),
.B1(n_17),
.B2(n_11),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_37),
.B1(n_27),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_15),
.B1(n_17),
.B2(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_13),
.B1(n_20),
.B2(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_14),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_50),
.B1(n_32),
.B2(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_57),
.B1(n_26),
.B2(n_23),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_48),
.Y(n_53)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_31),
.B1(n_34),
.B2(n_33),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_56),
.B(n_40),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_43),
.A3(n_47),
.B1(n_42),
.B2(n_50),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_49),
.B1(n_40),
.B2(n_34),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_24),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_0),
.B(n_1),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

AO21x2_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_40),
.B(n_26),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_57),
.B1(n_51),
.B2(n_23),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_24),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_70),
.B1(n_2),
.B2(n_3),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_0),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_59),
.C(n_58),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_78),
.B1(n_80),
.B2(n_4),
.Y(n_87)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_76),
.B(n_3),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_2),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_6),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_86),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_66),
.C(n_65),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_85),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

INVxp33_ASAP7_75t_SL g92 ( 
.A(n_84),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_65),
.C(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_79),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_82),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_96),
.Y(n_99)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_84),
.B(n_83),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_64),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_86),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_90),
.C(n_74),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_6),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_64),
.B(n_95),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_101),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_99),
.C(n_97),
.Y(n_105)
);


endmodule