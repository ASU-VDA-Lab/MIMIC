module real_aes_6655_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_575;
wire n_210;
wire n_212;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g261 ( .A1(n_0), .A2(n_262), .B(n_263), .C(n_266), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_1), .B(n_250), .Y(n_267) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_3), .B(n_178), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_4), .A2(n_139), .B(n_142), .C(n_555), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_5), .A2(n_134), .B(n_579), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_6), .A2(n_134), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_7), .B(n_250), .Y(n_585) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_8), .A2(n_169), .B(n_206), .Y(n_205) );
AND2x6_ASAP7_75t_L g139 ( .A(n_9), .B(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_10), .A2(n_139), .B(n_142), .C(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g523 ( .A(n_11), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_41), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_12), .B(n_41), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_13), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_13), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_14), .B(n_226), .Y(n_557) );
INVx1_ASAP7_75t_L g160 ( .A(n_15), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_16), .B(n_178), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_17), .A2(n_179), .B(n_541), .C(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_18), .B(n_250), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_19), .B(n_154), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_20), .A2(n_142), .B(n_145), .C(n_153), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_21), .A2(n_214), .B(n_265), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_22), .B(n_226), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_23), .A2(n_105), .B1(n_118), .B2(n_768), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_24), .A2(n_57), .B1(n_453), .B2(n_454), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_24), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_25), .B(n_226), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g570 ( .A(n_26), .Y(n_570) );
INVx1_ASAP7_75t_L g495 ( .A(n_27), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_28), .A2(n_142), .B(n_153), .C(n_209), .Y(n_208) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_29), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_30), .Y(n_553) );
INVx1_ASAP7_75t_L g511 ( .A(n_31), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_32), .A2(n_134), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g137 ( .A(n_33), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_34), .A2(n_182), .B(n_191), .C(n_193), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_35), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_36), .A2(n_265), .B(n_582), .C(n_584), .Y(n_581) );
INVxp67_ASAP7_75t_L g512 ( .A(n_37), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_38), .B(n_211), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_39), .A2(n_142), .B(n_153), .C(n_494), .Y(n_493) );
CKINVDCx14_ASAP7_75t_R g580 ( .A(n_40), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_42), .A2(n_266), .B(n_521), .C(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_43), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_44), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_45), .B(n_178), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_46), .B(n_134), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_47), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_48), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_49), .A2(n_182), .B(n_191), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_50), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g264 ( .A(n_51), .Y(n_264) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_52), .A2(n_451), .B1(n_452), .B2(n_455), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_52), .Y(n_455) );
AOI222xp33_ASAP7_75t_L g468 ( .A1(n_53), .A2(n_469), .B1(n_470), .B2(n_479), .C1(n_758), .C2(n_762), .Y(n_468) );
INVx1_ASAP7_75t_L g236 ( .A(n_54), .Y(n_236) );
INVx1_ASAP7_75t_L g529 ( .A(n_55), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_56), .B(n_134), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_57), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_58), .Y(n_162) );
CKINVDCx14_ASAP7_75t_R g519 ( .A(n_59), .Y(n_519) );
INVx1_ASAP7_75t_L g140 ( .A(n_60), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_61), .B(n_134), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_62), .B(n_250), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_63), .A2(n_152), .B(n_175), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g159 ( .A(n_64), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_65), .A2(n_103), .B1(n_475), .B2(n_476), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_65), .Y(n_476) );
INVx1_ASAP7_75t_SL g583 ( .A(n_66), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_68), .B(n_178), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_69), .B(n_250), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_70), .B(n_179), .Y(n_224) );
INVx1_ASAP7_75t_L g573 ( .A(n_71), .Y(n_573) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_72), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_73), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_74), .A2(n_142), .B(n_173), .C(n_182), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_75), .Y(n_245) );
INVx1_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_77), .A2(n_134), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_78), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_79), .A2(n_134), .B(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_80), .A2(n_133), .B(n_507), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_81), .Y(n_492) );
INVx1_ASAP7_75t_L g539 ( .A(n_82), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_83), .B(n_150), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_84), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_85), .A2(n_134), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g542 ( .A(n_86), .Y(n_542) );
INVx2_ASAP7_75t_L g157 ( .A(n_87), .Y(n_157) );
INVx1_ASAP7_75t_L g556 ( .A(n_88), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_89), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_90), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g114 ( .A(n_91), .Y(n_114) );
OR2x2_ASAP7_75t_L g460 ( .A(n_91), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g482 ( .A(n_91), .B(n_462), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g473 ( .A1(n_92), .A2(n_474), .B1(n_477), .B2(n_478), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_92), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_93), .A2(n_142), .B(n_182), .C(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_94), .B(n_134), .Y(n_189) );
INVx1_ASAP7_75t_L g194 ( .A(n_95), .Y(n_194) );
INVxp67_ASAP7_75t_L g248 ( .A(n_96), .Y(n_248) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_97), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_97), .B(n_169), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_98), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g174 ( .A(n_99), .Y(n_174) );
INVx1_ASAP7_75t_L g220 ( .A(n_100), .Y(n_220) );
INVx2_ASAP7_75t_L g532 ( .A(n_101), .Y(n_532) );
AND2x2_ASAP7_75t_L g238 ( .A(n_102), .B(n_156), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_103), .Y(n_475) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g769 ( .A(n_108), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g462 ( .A(n_113), .B(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g483 ( .A(n_114), .B(n_462), .Y(n_483) );
NOR2x2_ASAP7_75t_L g764 ( .A(n_114), .B(n_461), .Y(n_764) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_121), .B(n_467), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g767 ( .A(n_120), .Y(n_767) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_457), .B(n_464), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_449), .B1(n_450), .B2(n_456), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_124), .A2(n_485), .B1(n_759), .B2(n_760), .Y(n_758) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g456 ( .A(n_125), .Y(n_456) );
AND3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_353), .C(n_410), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_298), .C(n_334), .Y(n_126) );
OAI211xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_200), .B(n_252), .C(n_285), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_164), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g255 ( .A(n_130), .B(n_256), .Y(n_255) );
INVx5_ASAP7_75t_L g284 ( .A(n_130), .Y(n_284) );
AND2x2_ASAP7_75t_L g357 ( .A(n_130), .B(n_273), .Y(n_357) );
AND2x2_ASAP7_75t_L g395 ( .A(n_130), .B(n_301), .Y(n_395) );
AND2x2_ASAP7_75t_L g415 ( .A(n_130), .B(n_257), .Y(n_415) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_161), .Y(n_130) );
AOI21xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_141), .B(n_154), .Y(n_131) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_135), .B(n_139), .Y(n_221) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
INVx1_ASAP7_75t_L g215 ( .A(n_137), .Y(n_215) );
INVx1_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_138), .Y(n_148) );
INVx3_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
INVx1_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_138), .Y(n_226) );
BUFx3_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
INVx4_ASAP7_75t_SL g183 ( .A(n_139), .Y(n_183) );
INVx5_ASAP7_75t_L g192 ( .A(n_142), .Y(n_192) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
BUFx3_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B(n_151), .Y(n_145) );
INVx2_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_150), .A2(n_194), .B(n_195), .C(n_196), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_150), .A2(n_196), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp5_ASAP7_75t_L g555 ( .A1(n_150), .A2(n_556), .B(n_557), .C(n_558), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g572 ( .A1(n_150), .A2(n_558), .B(n_573), .C(n_574), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_151), .A2(n_178), .B(n_495), .C(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_152), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_155), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_156), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_156), .A2(n_233), .B(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_156), .A2(n_221), .B(n_492), .C(n_493), .Y(n_491) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_156), .A2(n_517), .B(n_524), .Y(n_516) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x2_ASAP7_75t_L g170 ( .A(n_157), .B(n_158), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_163), .A2(n_552), .B(n_559), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_164), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_187), .Y(n_164) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_165), .Y(n_296) );
AND2x2_ASAP7_75t_L g310 ( .A(n_165), .B(n_256), .Y(n_310) );
INVx1_ASAP7_75t_L g333 ( .A(n_165), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_165), .B(n_284), .Y(n_372) );
OR2x2_ASAP7_75t_L g409 ( .A(n_165), .B(n_254), .Y(n_409) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_166), .Y(n_345) );
AND2x2_ASAP7_75t_L g352 ( .A(n_166), .B(n_257), .Y(n_352) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g273 ( .A(n_167), .B(n_257), .Y(n_273) );
BUFx2_ASAP7_75t_L g301 ( .A(n_167), .Y(n_301) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_185), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_168), .B(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_168), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_168), .A2(n_219), .B(n_227), .Y(n_218) );
INVx3_ASAP7_75t_L g250 ( .A(n_168), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_168), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_168), .B(n_560), .Y(n_559) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_168), .A2(n_569), .B(n_575), .Y(n_568) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_169), .A2(n_207), .B(n_208), .Y(n_206) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_184), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_177), .C(n_180), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_176), .A2(n_178), .B1(n_511), .B2(n_512), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_176), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_176), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_178), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g262 ( .A(n_178), .Y(n_262) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_179), .B(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx3_ASAP7_75t_L g584 ( .A(n_181), .Y(n_584) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_183), .A2(n_192), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_183), .A2(n_192), .B(n_260), .C(n_261), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_183), .A2(n_192), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_183), .A2(n_192), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_183), .A2(n_192), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g538 ( .A1(n_183), .A2(n_192), .B(n_539), .C(n_540), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_183), .A2(n_192), .B(n_580), .C(n_581), .Y(n_579) );
INVx5_ASAP7_75t_L g254 ( .A(n_187), .Y(n_254) );
BUFx2_ASAP7_75t_L g277 ( .A(n_187), .Y(n_277) );
AND2x2_ASAP7_75t_L g434 ( .A(n_187), .B(n_288), .Y(n_434) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_198), .Y(n_187) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g266 ( .A(n_197), .Y(n_266) );
INVx1_ASAP7_75t_L g543 ( .A(n_197), .Y(n_543) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_239), .Y(n_201) );
OAI221xp5_ASAP7_75t_L g334 ( .A1(n_202), .A2(n_335), .B1(n_342), .B2(n_343), .C(n_346), .Y(n_334) );
OR2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_216), .Y(n_202) );
AND2x2_ASAP7_75t_L g240 ( .A(n_203), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_203), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g269 ( .A(n_204), .B(n_217), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_204), .B(n_218), .Y(n_279) );
OR2x2_ASAP7_75t_L g290 ( .A(n_204), .B(n_241), .Y(n_290) );
AND2x2_ASAP7_75t_L g293 ( .A(n_204), .B(n_281), .Y(n_293) );
AND2x2_ASAP7_75t_L g309 ( .A(n_204), .B(n_230), .Y(n_309) );
OR2x2_ASAP7_75t_L g325 ( .A(n_204), .B(n_218), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_204), .B(n_241), .Y(n_387) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_205), .B(n_230), .Y(n_379) );
AND2x2_ASAP7_75t_L g382 ( .A(n_205), .B(n_218), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_212), .B(n_213), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_213), .A2(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g303 ( .A(n_216), .B(n_290), .Y(n_303) );
INVx2_ASAP7_75t_L g329 ( .A(n_216), .Y(n_329) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_230), .Y(n_216) );
AND2x2_ASAP7_75t_L g251 ( .A(n_217), .B(n_231), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_217), .B(n_241), .Y(n_308) );
OR2x2_ASAP7_75t_L g319 ( .A(n_217), .B(n_231), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_217), .B(n_281), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_217), .A2(n_412), .B1(n_414), .B2(n_416), .C(n_419), .Y(n_411) );
INVx5_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_218), .B(n_241), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_221), .A2(n_553), .B(n_554), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_221), .A2(n_570), .B(n_571), .Y(n_569) );
INVx4_ASAP7_75t_L g265 ( .A(n_226), .Y(n_265) );
INVx2_ASAP7_75t_L g521 ( .A(n_226), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g504 ( .A(n_229), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_230), .B(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_230), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g297 ( .A(n_230), .B(n_269), .Y(n_297) );
OR2x2_ASAP7_75t_L g341 ( .A(n_230), .B(n_241), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_230), .B(n_293), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_230), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g406 ( .A(n_230), .B(n_407), .Y(n_406) );
INVx5_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_231), .B(n_240), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_SL g274 ( .A1(n_231), .A2(n_275), .B(n_278), .C(n_282), .Y(n_274) );
OR2x2_ASAP7_75t_L g312 ( .A(n_231), .B(n_308), .Y(n_312) );
OR2x2_ASAP7_75t_L g348 ( .A(n_231), .B(n_290), .Y(n_348) );
OAI311xp33_ASAP7_75t_L g354 ( .A1(n_231), .A2(n_293), .A3(n_355), .B1(n_358), .C1(n_365), .Y(n_354) );
AND2x2_ASAP7_75t_L g405 ( .A(n_231), .B(n_241), .Y(n_405) );
AND2x2_ASAP7_75t_L g413 ( .A(n_231), .B(n_268), .Y(n_413) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_231), .Y(n_431) );
AND2x2_ASAP7_75t_L g448 ( .A(n_231), .B(n_269), .Y(n_448) );
OR2x6_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_251), .Y(n_239) );
AND2x2_ASAP7_75t_L g276 ( .A(n_240), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g432 ( .A(n_240), .Y(n_432) );
AND2x2_ASAP7_75t_L g268 ( .A(n_241), .B(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g281 ( .A(n_241), .Y(n_281) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_241), .Y(n_324) );
INVxp67_ASAP7_75t_L g363 ( .A(n_241), .Y(n_363) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_249), .Y(n_241) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_242), .A2(n_527), .B(n_533), .Y(n_526) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_242), .A2(n_537), .B(n_544), .Y(n_536) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_242), .A2(n_578), .B(n_585), .Y(n_577) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_250), .A2(n_258), .B(n_267), .Y(n_257) );
AND2x2_ASAP7_75t_L g441 ( .A(n_251), .B(n_289), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_268), .B1(n_270), .B2(n_271), .C(n_274), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_254), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g294 ( .A(n_254), .B(n_284), .Y(n_294) );
AND2x2_ASAP7_75t_L g302 ( .A(n_254), .B(n_256), .Y(n_302) );
OR2x2_ASAP7_75t_L g314 ( .A(n_254), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g332 ( .A(n_254), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g356 ( .A(n_254), .B(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_254), .Y(n_376) );
AND2x2_ASAP7_75t_L g428 ( .A(n_254), .B(n_352), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g436 ( .A1(n_254), .A2(n_305), .A3(n_404), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_255), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g400 ( .A(n_255), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_255), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g288 ( .A(n_256), .B(n_284), .Y(n_288) );
INVx1_ASAP7_75t_L g375 ( .A(n_256), .Y(n_375) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g425 ( .A(n_257), .B(n_284), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_265), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g558 ( .A(n_266), .Y(n_558) );
INVx1_ASAP7_75t_SL g435 ( .A(n_268), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_269), .B(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_270), .A2(n_382), .B1(n_420), .B2(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g283 ( .A(n_273), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g342 ( .A(n_273), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_273), .B(n_294), .Y(n_447) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g417 ( .A(n_276), .B(n_418), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_277), .A2(n_336), .B(n_338), .Y(n_335) );
OR2x2_ASAP7_75t_L g343 ( .A(n_277), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g364 ( .A(n_277), .B(n_352), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_277), .B(n_375), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_277), .B(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_SL g391 ( .A1(n_278), .A2(n_392), .B1(n_397), .B2(n_400), .C(n_401), .Y(n_391) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OR2x2_ASAP7_75t_L g368 ( .A(n_279), .B(n_341), .Y(n_368) );
INVx1_ASAP7_75t_L g407 ( .A(n_279), .Y(n_407) );
INVx2_ASAP7_75t_L g383 ( .A(n_280), .Y(n_383) );
INVx1_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_284), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g351 ( .A(n_284), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g439 ( .A(n_284), .B(n_409), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .B1(n_291), .B2(n_294), .C1(n_295), .C2(n_297), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g295 ( .A(n_288), .B(n_296), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_288), .A2(n_338), .B1(n_366), .B2(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_288), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OAI21xp33_ASAP7_75t_SL g326 ( .A1(n_297), .A2(n_327), .B(n_330), .Y(n_326) );
OAI211xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_303), .B(n_304), .C(n_326), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_302), .A2(n_305), .B1(n_310), .B2(n_311), .C(n_313), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_302), .B(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_L g396 ( .A(n_302), .Y(n_396) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
AND2x2_ASAP7_75t_L g398 ( .A(n_307), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g315 ( .A(n_310), .Y(n_315) );
AND2x2_ASAP7_75t_L g321 ( .A(n_310), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_320), .B2(n_323), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_317), .B(n_329), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_318), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g418 ( .A(n_322), .Y(n_418) );
AND2x2_ASAP7_75t_L g437 ( .A(n_322), .B(n_352), .Y(n_437) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_329), .B(n_386), .Y(n_445) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_332), .B(n_400), .Y(n_443) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g366 ( .A(n_344), .Y(n_366) );
BUFx2_ASAP7_75t_L g390 ( .A(n_345), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_349), .B(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR3xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_369), .C(n_391), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_364), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_373), .B(n_377), .C(n_380), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_370), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NOR2xp67_ASAP7_75t_SL g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_SL g399 ( .A(n_379), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B(n_388), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g404 ( .A(n_382), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B1(n_406), .B2(n_408), .Y(n_401) );
INVx2_ASAP7_75t_SL g422 ( .A(n_409), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_426), .C(n_438), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_422), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_433), .B2(n_435), .C(n_436), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_427), .A2(n_439), .B(n_440), .C(n_442), .Y(n_438) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_446), .B2(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_456), .A2(n_480), .B1(n_483), .B2(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_460), .Y(n_466) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_464), .B(n_468), .C(n_765), .Y(n_467) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g477 ( .A(n_474), .Y(n_477) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g759 ( .A(n_481), .Y(n_759) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g761 ( .A(n_483), .Y(n_761) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
OR5x1_ASAP7_75t_L g485 ( .A(n_486), .B(n_652), .C(n_716), .D(n_732), .E(n_747), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_487), .B(n_586), .C(n_613), .D(n_636), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_534), .B(n_545), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_499), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_SL g565 ( .A(n_490), .Y(n_565) );
AND2x4_ASAP7_75t_L g599 ( .A(n_490), .B(n_588), .Y(n_599) );
OR2x2_ASAP7_75t_L g609 ( .A(n_490), .B(n_567), .Y(n_609) );
OR2x2_ASAP7_75t_L g655 ( .A(n_490), .B(n_502), .Y(n_655) );
AND2x2_ASAP7_75t_L g669 ( .A(n_490), .B(n_566), .Y(n_669) );
AND2x2_ASAP7_75t_L g712 ( .A(n_490), .B(n_602), .Y(n_712) );
AND2x2_ASAP7_75t_L g719 ( .A(n_490), .B(n_577), .Y(n_719) );
AND2x2_ASAP7_75t_L g738 ( .A(n_490), .B(n_628), .Y(n_738) );
AND2x2_ASAP7_75t_L g756 ( .A(n_490), .B(n_598), .Y(n_756) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_497), .Y(n_490) );
INVx1_ASAP7_75t_L g721 ( .A(n_499), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_515), .Y(n_499) );
AND2x2_ASAP7_75t_L g631 ( .A(n_500), .B(n_566), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_500), .B(n_651), .Y(n_650) );
AOI32xp33_ASAP7_75t_L g664 ( .A1(n_500), .A2(n_665), .A3(n_668), .B1(n_670), .B2(n_674), .Y(n_664) );
AND2x2_ASAP7_75t_L g734 ( .A(n_500), .B(n_628), .Y(n_734) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g598 ( .A(n_502), .B(n_567), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_502), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g640 ( .A(n_502), .B(n_587), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_502), .B(n_719), .Y(n_718) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_505), .B(n_513), .Y(n_502) );
INVx1_ASAP7_75t_L g603 ( .A(n_503), .Y(n_603) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OA21x2_ASAP7_75t_L g602 ( .A1(n_506), .A2(n_514), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g605 ( .A(n_515), .B(n_549), .Y(n_605) );
AND2x2_ASAP7_75t_L g681 ( .A(n_515), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g753 ( .A(n_515), .Y(n_753) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
OR2x2_ASAP7_75t_L g548 ( .A(n_516), .B(n_526), .Y(n_548) );
AND2x2_ASAP7_75t_L g562 ( .A(n_516), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_516), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g612 ( .A(n_516), .Y(n_612) );
AND2x2_ASAP7_75t_L g639 ( .A(n_516), .B(n_526), .Y(n_639) );
BUFx3_ASAP7_75t_L g642 ( .A(n_516), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_516), .B(n_617), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_516), .B(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g593 ( .A(n_525), .Y(n_593) );
AND2x2_ASAP7_75t_L g611 ( .A(n_525), .B(n_591), .Y(n_611) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g622 ( .A(n_526), .B(n_536), .Y(n_622) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_526), .Y(n_635) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_535), .B(n_642), .Y(n_692) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_SL g563 ( .A(n_536), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_536), .B(n_611), .C(n_612), .Y(n_610) );
OR2x2_ASAP7_75t_L g618 ( .A(n_536), .B(n_591), .Y(n_618) );
AND2x2_ASAP7_75t_L g638 ( .A(n_536), .B(n_591), .Y(n_638) );
AND2x2_ASAP7_75t_L g682 ( .A(n_536), .B(n_551), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_561), .B(n_564), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_L g757 ( .A(n_547), .B(n_682), .Y(n_757) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_548), .A2(n_655), .B1(n_697), .B2(n_699), .Y(n_696) );
OR2x2_ASAP7_75t_L g703 ( .A(n_548), .B(n_618), .Y(n_703) );
OR2x2_ASAP7_75t_L g727 ( .A(n_548), .B(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_548), .B(n_647), .Y(n_740) );
AND2x2_ASAP7_75t_L g633 ( .A(n_549), .B(n_634), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_549), .A2(n_706), .B(n_721), .Y(n_720) );
AOI32xp33_ASAP7_75t_L g741 ( .A1(n_549), .A2(n_631), .A3(n_742), .B1(n_744), .B2(n_745), .Y(n_741) );
OR2x2_ASAP7_75t_L g752 ( .A(n_549), .B(n_753), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g620 ( .A(n_550), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_550), .B(n_634), .Y(n_699) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g591 ( .A(n_551), .Y(n_591) );
AND2x2_ASAP7_75t_L g657 ( .A(n_551), .B(n_622), .Y(n_657) );
AND3x2_ASAP7_75t_L g666 ( .A(n_551), .B(n_562), .C(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g592 ( .A(n_563), .B(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_563), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_563), .B(n_591), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g587 ( .A(n_565), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g627 ( .A(n_565), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g645 ( .A(n_565), .B(n_577), .Y(n_645) );
AND2x2_ASAP7_75t_L g663 ( .A(n_565), .B(n_567), .Y(n_663) );
OR2x2_ASAP7_75t_L g677 ( .A(n_565), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g723 ( .A(n_565), .B(n_651), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_566), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_577), .Y(n_566) );
AND2x2_ASAP7_75t_L g624 ( .A(n_567), .B(n_602), .Y(n_624) );
OR2x2_ASAP7_75t_L g678 ( .A(n_567), .B(n_602), .Y(n_678) );
AND2x2_ASAP7_75t_L g731 ( .A(n_567), .B(n_588), .Y(n_731) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g629 ( .A(n_568), .Y(n_629) );
AND2x2_ASAP7_75t_L g651 ( .A(n_568), .B(n_577), .Y(n_651) );
INVx2_ASAP7_75t_L g588 ( .A(n_577), .Y(n_588) );
INVx1_ASAP7_75t_L g608 ( .A(n_577), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_594), .C(n_606), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_587), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g750 ( .A(n_587), .Y(n_750) );
AND2x2_ASAP7_75t_L g628 ( .A(n_588), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_591), .B(n_592), .Y(n_600) );
INVx1_ASAP7_75t_L g685 ( .A(n_591), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_591), .B(n_612), .Y(n_709) );
AND2x2_ASAP7_75t_L g725 ( .A(n_591), .B(n_639), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_592), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g616 ( .A(n_593), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_600), .B1(n_601), .B2(n_604), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_597), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_598), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g623 ( .A(n_599), .B(n_624), .Y(n_623) );
AOI221xp5_ASAP7_75t_SL g688 ( .A1(n_599), .A2(n_641), .B1(n_689), .B2(n_694), .C(n_696), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_599), .B(n_662), .Y(n_695) );
INVx1_ASAP7_75t_L g755 ( .A(n_601), .Y(n_755) );
BUFx3_ASAP7_75t_L g662 ( .A(n_602), .Y(n_662) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI21xp33_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_609), .B(n_610), .Y(n_606) );
INVx1_ASAP7_75t_L g671 ( .A(n_608), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_608), .B(n_662), .Y(n_715) );
INVx1_ASAP7_75t_L g672 ( .A(n_609), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_609), .B(n_662), .Y(n_673) );
INVxp67_ASAP7_75t_L g693 ( .A(n_611), .Y(n_693) );
AND2x2_ASAP7_75t_L g634 ( .A(n_612), .B(n_635), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_619), .B(n_623), .C(n_625), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_SL g648 ( .A(n_616), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_617), .B(n_648), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_617), .B(n_639), .Y(n_690) );
INVx2_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_620), .A2(n_626), .B1(n_630), .B2(n_632), .Y(n_625) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g641 ( .A(n_622), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g686 ( .A(n_622), .B(n_687), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_624), .A2(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_628), .A2(n_637), .B1(n_640), .B2(n_641), .C(n_643), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_628), .B(n_662), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_628), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g744 ( .A(n_634), .Y(n_744) );
INVxp67_ASAP7_75t_L g667 ( .A(n_635), .Y(n_667) );
INVx1_ASAP7_75t_L g674 ( .A(n_637), .Y(n_674) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g713 ( .A(n_638), .B(n_642), .Y(n_713) );
INVx1_ASAP7_75t_L g687 ( .A(n_642), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_642), .B(n_657), .Y(n_717) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .A3(n_648), .B1(n_649), .B2(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_SL g656 ( .A(n_651), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_651), .B(n_683), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_651), .B(n_712), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g751 ( .A(n_651), .B(n_662), .Y(n_751) );
NAND5xp2_ASAP7_75t_L g652 ( .A(n_653), .B(n_675), .C(n_688), .D(n_700), .E(n_701), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_657), .B1(n_658), .B2(n_660), .C(n_664), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_659), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_662), .B(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_663), .A2(n_676), .B1(n_679), .B2(n_683), .Y(n_675) );
INVx2_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_666), .A2(n_671), .B(n_672), .C(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g698 ( .A(n_678), .Y(n_698) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_687), .B(n_736), .Y(n_746) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_706), .B2(n_710), .C1(n_713), .C2(n_714), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_722), .C(n_724), .Y(n_716) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
OAI21xp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_729), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g736 ( .A(n_728), .Y(n_736) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B1(n_737), .B2(n_739), .C(n_741), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_751), .B(n_752), .C(n_754), .Y(n_747) );
INVxp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI21xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B(n_757), .Y(n_754) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
endmodule