module fake_netlist_1_6705_n_881 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_881);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_881;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_836;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g101 ( .A(n_55), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_87), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_84), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_85), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_9), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_68), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_75), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_13), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_29), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_50), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_24), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_86), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_49), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_37), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_40), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_36), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_43), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_42), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_67), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_66), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_58), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_73), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_21), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_47), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_18), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_99), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_18), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_45), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_26), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_76), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_0), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_74), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_62), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_20), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_53), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_70), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_24), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_41), .Y(n_144) );
BUFx12f_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_144), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_119), .B(n_0), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_144), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_144), .B(n_38), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_119), .B(n_1), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_114), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_127), .B(n_1), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_112), .B(n_2), .Y(n_154) );
BUFx8_ASAP7_75t_SL g155 ( .A(n_129), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_101), .B(n_2), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_127), .B(n_3), .Y(n_157) );
BUFx12f_ASAP7_75t_L g158 ( .A(n_103), .Y(n_158) );
BUFx12f_ASAP7_75t_L g159 ( .A(n_108), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_101), .B(n_3), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_114), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_104), .B(n_4), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_104), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_107), .B(n_4), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_107), .B(n_5), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_113), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_167), .B(n_106), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_164), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_165), .A2(n_143), .B1(n_109), .B2(n_110), .Y(n_171) );
OAI22xp33_ASAP7_75t_SL g172 ( .A1(n_148), .A2(n_117), .B1(n_135), .B2(n_140), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_153), .A2(n_157), .B1(n_165), .B2(n_151), .Y(n_174) );
OAI22xp33_ASAP7_75t_SL g175 ( .A1(n_148), .A2(n_137), .B1(n_115), .B2(n_118), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_153), .A2(n_129), .B1(n_115), .B2(n_118), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_167), .B(n_112), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_151), .A2(n_154), .B1(n_145), .B2(n_158), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_153), .A2(n_132), .B1(n_126), .B2(n_125), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_145), .B(n_113), .Y(n_183) );
BUFx10_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_167), .B(n_132), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_164), .B(n_102), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_164), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_157), .A2(n_142), .B1(n_116), .B2(n_121), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_165), .A2(n_142), .B1(n_116), .B2(n_121), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_164), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_164), .B(n_102), .Y(n_192) );
AO22x2_ASAP7_75t_L g193 ( .A1(n_165), .A2(n_126), .B1(n_122), .B2(n_123), .Y(n_193) );
BUFx6f_ASAP7_75t_SL g194 ( .A(n_165), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_157), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_158), .B(n_122), .Y(n_198) );
BUFx10_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
OAI22xp33_ASAP7_75t_L g200 ( .A1(n_154), .A2(n_130), .B1(n_123), .B2(n_125), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_146), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_158), .B(n_105), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_156), .A2(n_128), .B1(n_130), .B2(n_133), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_158), .B(n_105), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
OA22x2_ASAP7_75t_L g207 ( .A1(n_147), .A2(n_133), .B1(n_128), .B2(n_134), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g209 ( .A1(n_160), .A2(n_134), .B1(n_139), .B2(n_138), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_156), .A2(n_141), .B1(n_136), .B2(n_131), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_161), .B(n_111), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_159), .B(n_120), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_161), .B(n_147), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_199), .Y(n_215) );
OR2x6_ASAP7_75t_L g216 ( .A(n_197), .B(n_160), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_199), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_170), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_214), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_214), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_177), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
INVxp67_ASAP7_75t_SL g223 ( .A(n_206), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_174), .B(n_146), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_199), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_176), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_171), .B(n_159), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_169), .Y(n_229) );
OR2x6_ASAP7_75t_L g230 ( .A(n_197), .B(n_159), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_186), .B(n_159), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_177), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_185), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_185), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_186), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_178), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_192), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_192), .B(n_161), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_176), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_182), .B(n_162), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_181), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_187), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_181), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_188), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_188), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_195), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_195), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_182), .B(n_162), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_196), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_168), .B(n_166), .Y(n_250) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_196), .B(n_161), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_174), .B(n_166), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_211), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_180), .B(n_124), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_211), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_202), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_183), .B(n_155), .Y(n_260) );
XOR2x2_ASAP7_75t_L g261 ( .A(n_172), .B(n_155), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_198), .B(n_146), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_189), .B(n_150), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_206), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_193), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_187), .A2(n_150), .B(n_149), .Y(n_267) );
INVxp67_ASAP7_75t_SL g268 ( .A(n_193), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_193), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_212), .B(n_146), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_189), .B(n_150), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_212), .B(n_146), .Y(n_272) );
XOR2xp5_ASAP7_75t_L g273 ( .A(n_175), .B(n_5), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_190), .B(n_150), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_202), .B(n_205), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_207), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_256), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_225), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_253), .B(n_184), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_251), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_253), .B(n_200), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_275), .B(n_184), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_275), .B(n_184), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_263), .B(n_205), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_251), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_268), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_240), .B(n_191), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_225), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_224), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_225), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_263), .B(n_204), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_251), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_265), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_263), .B(n_204), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_224), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_230), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
INVx3_ASAP7_75t_SL g299 ( .A(n_224), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_229), .A2(n_207), .B(n_191), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_240), .B(n_207), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_240), .B(n_209), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_248), .B(n_213), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_248), .B(n_150), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_235), .B(n_194), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_229), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_252), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_266), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_252), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_248), .B(n_150), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_215), .Y(n_312) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_269), .Y(n_313) );
BUFx5_ASAP7_75t_L g314 ( .A(n_219), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_241), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_238), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_243), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_238), .B(n_150), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_244), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_271), .B(n_150), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_271), .A2(n_210), .B(n_208), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_221), .B(n_150), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_245), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_224), .B(n_150), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_218), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_246), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_280), .Y(n_329) );
BUFx4f_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_280), .B(n_285), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_286), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_293), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_298), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_293), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_280), .B(n_215), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_279), .B(n_237), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_279), .B(n_247), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_293), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_279), .B(n_249), .Y(n_342) );
BUFx8_ASAP7_75t_L g343 ( .A(n_321), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_279), .B(n_232), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_321), .B(n_274), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_292), .B(n_233), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_280), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_293), .Y(n_348) );
AND2x2_ASAP7_75t_SL g349 ( .A(n_321), .B(n_274), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_298), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_285), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_292), .B(n_234), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_314), .B(n_255), .Y(n_353) );
BUFx4f_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_285), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_292), .B(n_259), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_314), .B(n_224), .Y(n_357) );
AO21x2_ASAP7_75t_L g358 ( .A1(n_322), .A2(n_267), .B(n_276), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_292), .B(n_274), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_351), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_355), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_329), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_346), .B(n_352), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_351), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_355), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_337), .B(n_307), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_343), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_334), .B(n_290), .Y(n_369) );
BUFx12f_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_337), .B(n_307), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_355), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_334), .Y(n_375) );
BUFx4f_ASAP7_75t_L g376 ( .A(n_351), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_331), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_351), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_343), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_359), .A2(n_292), .B1(n_295), .B2(n_226), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_331), .B(n_285), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_350), .B(n_290), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
BUFx10_ASAP7_75t_L g386 ( .A(n_331), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_351), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_381), .A2(n_226), .B1(n_239), .B2(n_347), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_370), .Y(n_390) );
OAI22xp5_ASAP7_75t_SL g391 ( .A1(n_368), .A2(n_239), .B1(n_254), .B2(n_258), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_370), .A2(n_349), .B1(n_258), .B2(n_254), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_370), .A2(n_349), .B1(n_345), .B2(n_356), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_362), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_382), .Y(n_396) );
OAI21xp5_ASAP7_75t_SL g397 ( .A1(n_381), .A2(n_321), .B(n_273), .Y(n_397) );
BUFx12f_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_376), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_380), .A2(n_349), .B1(n_345), .B2(n_356), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_365), .Y(n_401) );
CKINVDCx11_ASAP7_75t_R g402 ( .A(n_368), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_365), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_365), .Y(n_404) );
CKINVDCx11_ASAP7_75t_R g405 ( .A(n_386), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_373), .Y(n_409) );
BUFx4_ASAP7_75t_SL g410 ( .A(n_380), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_380), .A2(n_343), .B1(n_349), .B2(n_347), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_363), .B(n_346), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_376), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_361), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_375), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_375), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_380), .A2(n_297), .B1(n_356), .B2(n_345), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_361), .Y(n_419) );
CKINVDCx11_ASAP7_75t_R g420 ( .A(n_386), .Y(n_420) );
INVx6_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
INVx6_ASAP7_75t_L g422 ( .A(n_386), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_362), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_383), .A2(n_349), .B1(n_345), .B2(n_295), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_361), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_361), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_381), .A2(n_332), .B1(n_350), .B2(n_345), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_375), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_363), .B(n_346), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_363), .A2(n_295), .B1(n_344), .B2(n_346), .Y(n_430) );
BUFx8_ASAP7_75t_SL g431 ( .A(n_383), .Y(n_431) );
HB1xp67_ASAP7_75t_SL g432 ( .A(n_383), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_389), .A2(n_383), .B1(n_363), .B2(n_343), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_407), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_396), .B(n_382), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_397), .A2(n_383), .B1(n_361), .B2(n_372), .Y(n_436) );
CKINVDCx8_ASAP7_75t_R g437 ( .A(n_390), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_397), .A2(n_259), .B1(n_273), .B2(n_297), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_427), .A2(n_366), .B1(n_372), .B2(n_374), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_412), .A2(n_366), .B1(n_372), .B2(n_374), .Y(n_440) );
INVx6_ASAP7_75t_L g441 ( .A(n_398), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_389), .A2(n_352), .B1(n_382), .B2(n_359), .Y(n_442) );
OAI222xp33_ASAP7_75t_L g443 ( .A1(n_427), .A2(n_362), .B1(n_377), .B2(n_388), .C1(n_385), .C2(n_345), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_413), .B(n_331), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_421), .A2(n_366), .B1(n_372), .B2(n_374), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_406), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_398), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_411), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_405), .B(n_382), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_413), .B(n_331), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_420), .B(n_382), .Y(n_455) );
OAI21xp5_ASAP7_75t_SL g456 ( .A1(n_392), .A2(n_311), .B(n_305), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_432), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_431), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_398), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_394), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_394), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_400), .A2(n_374), .B1(n_366), .B2(n_377), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_393), .A2(n_377), .B1(n_345), .B2(n_382), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_432), .A2(n_377), .B1(n_345), .B2(n_382), .Y(n_465) );
BUFx5_ASAP7_75t_L g466 ( .A(n_407), .Y(n_466) );
AOI22xp5_ASAP7_75t_SL g467 ( .A1(n_410), .A2(n_331), .B1(n_388), .B2(n_261), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_411), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_391), .B(n_260), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_421), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_418), .A2(n_352), .B1(n_296), .B2(n_290), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_421), .Y(n_473) );
CKINVDCx11_ASAP7_75t_R g474 ( .A(n_415), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_391), .A2(n_352), .B1(n_296), .B2(n_290), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_424), .A2(n_332), .B1(n_367), .B2(n_371), .Y(n_476) );
AOI222xp33_ASAP7_75t_L g477 ( .A1(n_429), .A2(n_295), .B1(n_303), .B2(n_304), .C1(n_302), .C2(n_261), .Y(n_477) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_416), .A2(n_228), .B(n_303), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_421), .A2(n_296), .B1(n_290), .B2(n_344), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_429), .A2(n_359), .B1(n_386), .B2(n_344), .Y(n_481) );
OAI21xp33_ASAP7_75t_L g482 ( .A1(n_417), .A2(n_303), .B(n_305), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_421), .A2(n_367), .B1(n_371), .B2(n_335), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_422), .A2(n_386), .B1(n_376), .B2(n_351), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_422), .Y(n_485) );
OAI222xp33_ASAP7_75t_L g486 ( .A1(n_415), .A2(n_385), .B1(n_371), .B2(n_367), .C1(n_378), .C2(n_335), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_428), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_422), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_419), .B(n_385), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_422), .A2(n_296), .B1(n_344), .B2(n_338), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_430), .B(n_302), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_422), .A2(n_296), .B1(n_338), .B2(n_386), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_428), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_394), .B(n_302), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_419), .A2(n_338), .B1(n_359), .B2(n_224), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_414), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_425), .A2(n_338), .B1(n_302), .B2(n_339), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_425), .A2(n_335), .B1(n_376), .B2(n_286), .Y(n_498) );
INVx6_ASAP7_75t_L g499 ( .A(n_426), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_426), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_399), .A2(n_376), .B1(n_351), .B2(n_378), .Y(n_501) );
BUFx12f_ASAP7_75t_L g502 ( .A(n_399), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_401), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_503), .B(n_401), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_467), .A2(n_399), .B1(n_414), .B2(n_395), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_433), .A2(n_414), .B1(n_311), .B2(n_305), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_447), .B(n_401), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_464), .A2(n_311), .B1(n_302), .B2(n_351), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_438), .A2(n_351), .B1(n_408), .B2(n_404), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_477), .A2(n_299), .B1(n_340), .B2(n_337), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_446), .B(n_304), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_439), .A2(n_299), .B1(n_340), .B2(n_357), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_449), .B(n_403), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_470), .A2(n_299), .B1(n_325), .B2(n_336), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_436), .A2(n_325), .B1(n_336), .B2(n_284), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g516 ( .A1(n_442), .A2(n_304), .B1(n_281), .B2(n_284), .C1(n_339), .C2(n_342), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_442), .A2(n_336), .B1(n_284), .B2(n_342), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_465), .A2(n_325), .B1(n_336), .B2(n_284), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_441), .A2(n_423), .B1(n_395), .B2(n_404), .Y(n_519) );
OAI211xp5_ASAP7_75t_SL g520 ( .A1(n_437), .A2(n_281), .B(n_287), .C(n_250), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_441), .A2(n_423), .B1(n_408), .B2(n_404), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_450), .B(n_403), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_497), .A2(n_378), .B1(n_403), .B2(n_408), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_475), .A2(n_325), .B1(n_336), .B2(n_360), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_474), .A2(n_325), .B1(n_360), .B2(n_379), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_484), .B(n_163), .C(n_152), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_497), .A2(n_325), .B1(n_360), .B2(n_379), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_441), .A2(n_378), .B1(n_360), .B2(n_230), .Y(n_528) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_486), .A2(n_378), .B(n_301), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_451), .B(n_360), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_491), .A2(n_281), .B1(n_301), .B2(n_287), .C1(n_257), .C2(n_353), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_476), .A2(n_325), .B1(n_387), .B2(n_379), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_495), .A2(n_387), .B1(n_379), .B2(n_364), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_463), .A2(n_387), .B1(n_379), .B2(n_364), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_481), .A2(n_369), .B1(n_384), .B2(n_379), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_472), .A2(n_387), .B1(n_379), .B2(n_364), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_500), .A2(n_387), .B1(n_379), .B2(n_364), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_452), .B(n_364), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_468), .B(n_364), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_478), .A2(n_387), .B1(n_379), .B2(n_364), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_469), .B(n_364), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_459), .B(n_236), .C(n_287), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_479), .B(n_364), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_440), .A2(n_387), .B1(n_348), .B2(n_341), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_482), .A2(n_387), .B1(n_348), .B2(n_341), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_459), .A2(n_230), .B1(n_369), .B2(n_384), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_445), .A2(n_369), .B1(n_384), .B2(n_328), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_484), .A2(n_369), .B1(n_384), .B2(n_236), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_435), .A2(n_328), .B1(n_333), .B2(n_341), .Y(n_549) );
NAND2xp33_ASAP7_75t_SL g550 ( .A(n_488), .B(n_328), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_487), .B(n_328), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_483), .A2(n_328), .B1(n_333), .B2(n_341), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_490), .A2(n_328), .B1(n_333), .B2(n_341), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_445), .A2(n_502), .B1(n_454), .B2(n_444), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_461), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_460), .A2(n_369), .B1(n_384), .B2(n_333), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_501), .B(n_163), .C(n_152), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_485), .A2(n_328), .B1(n_333), .B2(n_341), .Y(n_558) );
OAI222xp33_ASAP7_75t_L g559 ( .A1(n_457), .A2(n_369), .B1(n_216), .B2(n_353), .C1(n_316), .C2(n_327), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_493), .B(n_328), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_485), .A2(n_328), .B1(n_333), .B2(n_348), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_489), .B(n_333), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_462), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_489), .A2(n_473), .B1(n_492), .B2(n_458), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_456), .A2(n_319), .B1(n_315), .B2(n_317), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_448), .A2(n_319), .B1(n_315), .B2(n_317), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_496), .B(n_333), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_457), .A2(n_333), .B1(n_341), .B2(n_348), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_496), .Y(n_569) );
OAI221xp5_ASAP7_75t_SL g570 ( .A1(n_453), .A2(n_216), .B1(n_231), .B2(n_320), .C(n_316), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_455), .A2(n_341), .B1(n_348), .B2(n_319), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_499), .A2(n_348), .B1(n_317), .B2(n_315), .Y(n_572) );
OAI221xp5_ASAP7_75t_SL g573 ( .A1(n_471), .A2(n_216), .B1(n_320), .B2(n_316), .C(n_323), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_499), .A2(n_348), .B1(n_319), .B2(n_327), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_466), .A2(n_324), .B1(n_327), .B2(n_294), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g576 ( .A1(n_501), .A2(n_216), .B1(n_306), .B2(n_301), .C(n_322), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_480), .A2(n_313), .B1(n_309), .B2(n_324), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_466), .A2(n_324), .B1(n_327), .B2(n_294), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_466), .A2(n_324), .B1(n_294), .B2(n_320), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_466), .A2(n_320), .B1(n_310), .B2(n_298), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_494), .B(n_314), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_466), .A2(n_300), .B1(n_310), .B2(n_298), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_466), .A2(n_300), .B1(n_310), .B2(n_298), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_434), .B(n_314), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g585 ( .A1(n_443), .A2(n_486), .B(n_498), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_434), .B(n_314), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_434), .A2(n_310), .B1(n_300), .B2(n_308), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_443), .A2(n_310), .B1(n_300), .B2(n_308), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_467), .A2(n_354), .B1(n_330), .B2(n_314), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_503), .B(n_152), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_433), .A2(n_300), .B1(n_308), .B2(n_314), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_447), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_433), .A2(n_323), .B(n_306), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_433), .A2(n_308), .B1(n_314), .B2(n_150), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_433), .A2(n_314), .B1(n_313), .B2(n_309), .Y(n_595) );
AOI221xp5_ASAP7_75t_SL g596 ( .A1(n_433), .A2(n_152), .B1(n_163), .B2(n_149), .C(n_322), .Y(n_596) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_460), .B(n_330), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_499), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_505), .A2(n_152), .B1(n_163), .B2(n_306), .C(n_149), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_542), .A2(n_314), .B1(n_309), .B2(n_323), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_593), .B(n_6), .Y(n_601) );
NAND4xp25_ASAP7_75t_SL g602 ( .A(n_589), .B(n_6), .C(n_7), .D(n_8), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_511), .B(n_152), .C(n_163), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_504), .B(n_152), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_504), .B(n_7), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_592), .B(n_8), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_538), .B(n_163), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_510), .A2(n_314), .B1(n_163), .B2(n_149), .Y(n_608) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_585), .A2(n_163), .B(n_149), .Y(n_609) );
OA21x2_ASAP7_75t_L g610 ( .A1(n_585), .A2(n_262), .B(n_173), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_565), .A2(n_354), .B1(n_330), .B2(n_291), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_592), .B(n_9), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_563), .B(n_10), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_538), .B(n_149), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_564), .A2(n_149), .B1(n_323), .B2(n_270), .C(n_272), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_520), .B(n_318), .C(n_288), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_555), .B(n_10), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_516), .A2(n_314), .B1(n_289), .B2(n_277), .Y(n_618) );
OAI21xp5_ASAP7_75t_SL g619 ( .A1(n_565), .A2(n_318), .B(n_282), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_516), .A2(n_314), .B1(n_289), .B2(n_277), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_521), .B(n_330), .Y(n_621) );
OA21x2_ASAP7_75t_L g622 ( .A1(n_596), .A2(n_173), .B(n_201), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_563), .B(n_11), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_590), .B(n_11), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_569), .B(n_179), .C(n_201), .Y(n_625) );
OA211x2_ASAP7_75t_L g626 ( .A1(n_588), .A2(n_12), .B(n_13), .C(n_14), .Y(n_626) );
OAI221xp5_ASAP7_75t_SL g627 ( .A1(n_593), .A2(n_318), .B1(n_277), .B2(n_289), .C(n_283), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_598), .B(n_12), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_598), .B(n_14), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_590), .B(n_15), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_567), .B(n_15), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_560), .B(n_16), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_560), .B(n_16), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_554), .B(n_17), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_507), .B(n_17), .Y(n_635) );
OAI221xp5_ASAP7_75t_SL g636 ( .A1(n_517), .A2(n_318), .B1(n_277), .B2(n_289), .C(n_283), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_569), .B(n_179), .C(n_208), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_513), .B(n_19), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_522), .B(n_20), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_555), .B(n_21), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_530), .B(n_22), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_523), .B(n_22), .Y(n_642) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_597), .B(n_330), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_526), .B(n_179), .C(n_210), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_509), .A2(n_179), .B1(n_220), .B2(n_282), .C(n_283), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_519), .B(n_354), .Y(n_646) );
NAND2xp33_ASAP7_75t_SL g647 ( .A(n_547), .B(n_194), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_523), .B(n_23), .Y(n_648) );
OA21x2_ASAP7_75t_L g649 ( .A1(n_557), .A2(n_277), .B(n_289), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_531), .B(n_23), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_508), .A2(n_314), .B1(n_358), .B2(n_354), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_531), .B(n_25), .Y(n_652) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_547), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_537), .B(n_354), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g655 ( .A1(n_548), .A2(n_25), .B(n_26), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_566), .A2(n_291), .B1(n_288), .B2(n_278), .C(n_312), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_556), .B(n_314), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_539), .B(n_27), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_526), .B(n_326), .C(n_291), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_528), .A2(n_314), .B1(n_291), .B2(n_358), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_570), .B(n_283), .C(n_282), .D(n_30), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_541), .B(n_28), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_567), .B(n_28), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_562), .B(n_29), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_597), .B(n_30), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_597), .B(n_31), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_573), .B(n_278), .C(n_288), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_549), .B(n_31), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_566), .A2(n_291), .B1(n_278), .B2(n_288), .C(n_312), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_543), .B(n_32), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_559), .B(n_576), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_546), .B(n_278), .C(n_288), .Y(n_672) );
NOR2xp33_ASAP7_75t_SL g673 ( .A(n_535), .B(n_314), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_515), .A2(n_312), .B1(n_278), .B2(n_288), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_551), .B(n_33), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_532), .B(n_34), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_594), .A2(n_326), .B(n_36), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_552), .B(n_35), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g679 ( .A1(n_517), .A2(n_282), .B1(n_37), .B2(n_35), .C(n_326), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_529), .B(n_39), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_529), .B(n_314), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g682 ( .A1(n_529), .A2(n_586), .B(n_584), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_529), .B(n_358), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_534), .B(n_44), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_535), .B(n_46), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_544), .B(n_48), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_512), .B(n_326), .C(n_288), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_518), .A2(n_312), .B1(n_278), .B2(n_326), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_525), .A2(n_312), .B1(n_278), .B2(n_194), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_581), .B(n_358), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_540), .B(n_51), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_571), .B(n_52), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_591), .A2(n_312), .B1(n_217), .B2(n_223), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_568), .B(n_54), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_572), .B(n_56), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_506), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_696) );
OAI21xp5_ASAP7_75t_SL g697 ( .A1(n_595), .A2(n_63), .B(n_64), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_650), .B(n_577), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_604), .B(n_533), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_610), .B(n_550), .C(n_536), .Y(n_700) );
NAND4xp75_ASAP7_75t_L g701 ( .A(n_610), .B(n_527), .C(n_524), .D(n_574), .Y(n_701) );
NAND4xp75_ASAP7_75t_L g702 ( .A(n_610), .B(n_514), .C(n_553), .D(n_580), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_690), .B(n_558), .Y(n_703) );
BUFx3_ASAP7_75t_L g704 ( .A(n_607), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_653), .B(n_561), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_607), .B(n_583), .Y(n_706) );
NOR2x1_ASAP7_75t_R g707 ( .A(n_665), .B(n_577), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_614), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_671), .B(n_545), .C(n_582), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_671), .A2(n_579), .B1(n_578), .B2(n_575), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_652), .B(n_587), .C(n_242), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_634), .B(n_242), .C(n_222), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_614), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_617), .Y(n_714) );
NOR3xp33_ASAP7_75t_SL g715 ( .A(n_661), .B(n_65), .C(n_69), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_647), .B(n_222), .C(n_218), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_628), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_602), .B(n_71), .C(n_72), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_605), .B(n_77), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_617), .Y(n_720) );
AO21x2_ASAP7_75t_L g721 ( .A1(n_680), .A2(n_78), .B(n_79), .Y(n_721) );
AO21x2_ASAP7_75t_L g722 ( .A1(n_680), .A2(n_81), .B(n_82), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_640), .Y(n_723) );
BUFx2_ASAP7_75t_L g724 ( .A(n_647), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_603), .B(n_88), .C(n_89), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_681), .B(n_90), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_601), .B(n_91), .C(n_92), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_632), .B(n_94), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_601), .B(n_95), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_618), .A2(n_96), .B1(n_97), .B2(n_98), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_643), .B(n_100), .Y(n_731) );
NAND4xp75_ASAP7_75t_L g732 ( .A(n_666), .B(n_643), .C(n_646), .D(n_626), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_657), .B(n_682), .C(n_673), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_618), .A2(n_620), .B1(n_672), .B2(n_616), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_633), .B(n_631), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_663), .B(n_664), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_642), .B(n_648), .C(n_635), .Y(n_737) );
AO21x2_ASAP7_75t_L g738 ( .A1(n_606), .A2(n_612), .B(n_623), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_685), .B(n_654), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_683), .B(n_658), .Y(n_740) );
AO21x2_ASAP7_75t_L g741 ( .A1(n_613), .A2(n_662), .B(n_670), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_629), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_685), .B(n_654), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_638), .B(n_639), .C(n_621), .Y(n_744) );
OAI221xp5_ASAP7_75t_SL g745 ( .A1(n_619), .A2(n_620), .B1(n_697), .B2(n_677), .C(n_651), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_649), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_655), .B(n_679), .C(n_641), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_624), .B(n_630), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_621), .B(n_675), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_660), .B(n_668), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_691), .B(n_684), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_676), .A2(n_615), .B1(n_678), .B2(n_651), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_691), .B(n_684), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_622), .Y(n_754) );
INVx2_ASAP7_75t_SL g755 ( .A(n_694), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_686), .B(n_692), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_599), .B(n_659), .C(n_645), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_627), .B(n_696), .C(n_636), .Y(n_758) );
NAND4xp75_ASAP7_75t_L g759 ( .A(n_622), .B(n_686), .C(n_695), .D(n_600), .Y(n_759) );
NAND4xp75_ASAP7_75t_L g760 ( .A(n_622), .B(n_611), .C(n_687), .D(n_689), .Y(n_760) );
NAND4xp25_ASAP7_75t_L g761 ( .A(n_608), .B(n_667), .C(n_656), .D(n_669), .Y(n_761) );
OR2x6_ASAP7_75t_L g762 ( .A(n_644), .B(n_625), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_608), .B(n_637), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_688), .B(n_674), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_693), .B(n_609), .C(n_610), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_650), .B(n_652), .Y(n_766) );
INVx2_ASAP7_75t_SL g767 ( .A(n_604), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_609), .B(n_610), .C(n_671), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_604), .B(n_607), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_604), .B(n_607), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_704), .Y(n_771) );
INVx5_ASAP7_75t_L g772 ( .A(n_762), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_705), .B(n_740), .Y(n_773) );
NOR4xp25_ASAP7_75t_L g774 ( .A(n_768), .B(n_745), .C(n_766), .D(n_723), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_717), .B(n_707), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_704), .Y(n_776) );
OAI22xp5_ASAP7_75t_SL g777 ( .A1(n_717), .A2(n_724), .B1(n_716), .B2(n_765), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_708), .B(n_713), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_767), .Y(n_779) );
NAND4xp25_ASAP7_75t_L g780 ( .A(n_745), .B(n_744), .C(n_698), .D(n_747), .Y(n_780) );
NAND4xp75_ASAP7_75t_SL g781 ( .A(n_729), .B(n_731), .C(n_698), .D(n_743), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_720), .B(n_703), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_714), .B(n_770), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_769), .Y(n_784) );
NOR3xp33_ASAP7_75t_SL g785 ( .A(n_701), .B(n_702), .C(n_732), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_739), .B(n_749), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_699), .B(n_742), .Y(n_787) );
XNOR2xp5_ASAP7_75t_L g788 ( .A(n_736), .B(n_735), .Y(n_788) );
OAI31xp33_ASAP7_75t_L g789 ( .A1(n_709), .A2(n_757), .A3(n_733), .B(n_737), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_750), .B(n_738), .Y(n_790) );
XNOR2xp5_ASAP7_75t_L g791 ( .A(n_748), .B(n_710), .Y(n_791) );
XNOR2x2_ASAP7_75t_L g792 ( .A(n_760), .B(n_759), .Y(n_792) );
NAND4xp25_ASAP7_75t_SL g793 ( .A(n_758), .B(n_734), .C(n_718), .D(n_753), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_738), .Y(n_794) );
NAND4xp75_ASAP7_75t_L g795 ( .A(n_715), .B(n_729), .C(n_764), .D(n_755), .Y(n_795) );
XOR2x2_ASAP7_75t_L g796 ( .A(n_758), .B(n_718), .Y(n_796) );
XNOR2xp5_ASAP7_75t_L g797 ( .A(n_751), .B(n_756), .Y(n_797) );
XOR2x2_ASAP7_75t_L g798 ( .A(n_747), .B(n_727), .Y(n_798) );
INVx1_ASAP7_75t_SL g799 ( .A(n_706), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_719), .Y(n_800) );
AND2x4_ASAP7_75t_L g801 ( .A(n_700), .B(n_746), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_741), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_741), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_761), .B(n_752), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_752), .B(n_763), .Y(n_805) );
NAND2xp33_ASAP7_75t_L g806 ( .A(n_712), .B(n_711), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_746), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_754), .B(n_762), .Y(n_808) );
XOR2x2_ASAP7_75t_L g809 ( .A(n_734), .B(n_711), .Y(n_809) );
INVx2_ASAP7_75t_SL g810 ( .A(n_762), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_712), .B(n_726), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_721), .B(n_722), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_783), .Y(n_813) );
INVxp67_ASAP7_75t_L g814 ( .A(n_775), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_775), .A2(n_730), .B1(n_725), .B2(n_728), .Y(n_815) );
XOR2x2_ASAP7_75t_L g816 ( .A(n_796), .B(n_791), .Y(n_816) );
XNOR2xp5_ASAP7_75t_L g817 ( .A(n_785), .B(n_730), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_783), .Y(n_818) );
INVx2_ASAP7_75t_SL g819 ( .A(n_771), .Y(n_819) );
OA22x2_ASAP7_75t_L g820 ( .A1(n_777), .A2(n_805), .B1(n_810), .B2(n_801), .Y(n_820) );
OA22x2_ASAP7_75t_L g821 ( .A1(n_810), .A2(n_801), .B1(n_788), .B2(n_774), .Y(n_821) );
INVxp67_ASAP7_75t_L g822 ( .A(n_804), .Y(n_822) );
INVx1_ASAP7_75t_SL g823 ( .A(n_808), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_790), .B(n_802), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_782), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_808), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_778), .Y(n_827) );
INVxp67_ASAP7_75t_L g828 ( .A(n_804), .Y(n_828) );
INVxp67_ASAP7_75t_L g829 ( .A(n_780), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_803), .B(n_794), .Y(n_830) );
INVxp67_ASAP7_75t_L g831 ( .A(n_793), .Y(n_831) );
XOR2x2_ASAP7_75t_L g832 ( .A(n_809), .B(n_781), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_784), .Y(n_833) );
XOR2x2_ASAP7_75t_L g834 ( .A(n_809), .B(n_792), .Y(n_834) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_829), .Y(n_835) );
AOI22x1_ASAP7_75t_L g836 ( .A1(n_831), .A2(n_801), .B1(n_792), .B2(n_776), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_827), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_813), .Y(n_838) );
OA22x2_ASAP7_75t_L g839 ( .A1(n_822), .A2(n_799), .B1(n_797), .B2(n_789), .Y(n_839) );
OA22x2_ASAP7_75t_L g840 ( .A1(n_822), .A2(n_797), .B1(n_776), .B2(n_786), .Y(n_840) );
AOI22x1_ASAP7_75t_L g841 ( .A1(n_817), .A2(n_798), .B1(n_800), .B2(n_779), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_818), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_833), .Y(n_843) );
INVx1_ASAP7_75t_SL g844 ( .A(n_823), .Y(n_844) );
BUFx2_ASAP7_75t_L g845 ( .A(n_819), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_820), .A2(n_772), .B1(n_773), .B2(n_795), .Y(n_846) );
AO22x1_ASAP7_75t_L g847 ( .A1(n_814), .A2(n_772), .B1(n_812), .B2(n_811), .Y(n_847) );
OAI22x1_ASAP7_75t_SL g848 ( .A1(n_834), .A2(n_772), .B1(n_798), .B2(n_807), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_821), .A2(n_806), .B1(n_772), .B2(n_786), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_844), .Y(n_850) );
XOR2x2_ASAP7_75t_L g851 ( .A(n_839), .B(n_816), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_837), .Y(n_852) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_844), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_843), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_838), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_842), .Y(n_856) );
AOI322xp5_ASAP7_75t_L g857 ( .A1(n_835), .A2(n_828), .A3(n_821), .B1(n_823), .B2(n_826), .C1(n_825), .C2(n_787), .Y(n_857) );
INVx2_ASAP7_75t_SL g858 ( .A(n_850), .Y(n_858) );
INVx2_ASAP7_75t_SL g859 ( .A(n_850), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_853), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_852), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_852), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_858), .Y(n_863) );
INVx2_ASAP7_75t_SL g864 ( .A(n_858), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_860), .A2(n_849), .B1(n_839), .B2(n_841), .Y(n_865) );
AO22x2_ASAP7_75t_L g866 ( .A1(n_865), .A2(n_863), .B1(n_864), .B2(n_859), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_865), .A2(n_851), .B1(n_832), .B2(n_820), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_866), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_867), .A2(n_851), .B1(n_848), .B2(n_846), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_869), .A2(n_859), .B1(n_836), .B2(n_840), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_868), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_871), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_870), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_873), .A2(n_862), .B1(n_861), .B2(n_840), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_874), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_875), .A2(n_873), .B1(n_872), .B2(n_845), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_876), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_877), .A2(n_856), .B1(n_855), .B2(n_854), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_878), .Y(n_879) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_879), .A2(n_847), .B1(n_826), .B2(n_824), .C(n_857), .Y(n_880) );
AOI211xp5_ASAP7_75t_L g881 ( .A1(n_880), .A2(n_815), .B(n_824), .C(n_830), .Y(n_881) );
endmodule