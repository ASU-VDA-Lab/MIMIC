module real_jpeg_6805_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_1),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_1),
.A2(n_205),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_1),
.A2(n_174),
.B1(n_193),
.B2(n_205),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_1),
.A2(n_198),
.B1(n_205),
.B2(n_415),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_2),
.A2(n_244),
.B1(n_246),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_259),
.C(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_2),
.B(n_145),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_2),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_2),
.B(n_89),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_2),
.B(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_4),
.A2(n_155),
.B1(n_158),
.B2(n_161),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_4),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_161),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_4),
.A2(n_99),
.B1(n_161),
.B2(n_216),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_4),
.A2(n_161),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_6),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_6),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_6),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_9),
.A2(n_49),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_9),
.A2(n_38),
.B1(n_49),
.B2(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g387 ( 
.A(n_10),
.Y(n_387)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_10),
.Y(n_439)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_11),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_11),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_95),
.B1(n_166),
.B2(n_198),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_11),
.A2(n_95),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_11),
.A2(n_95),
.B1(n_191),
.B2(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_12),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_12),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_12),
.A2(n_115),
.B1(n_174),
.B2(n_252),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_12),
.A2(n_115),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_12),
.A2(n_115),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_13),
.A2(n_192),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_13),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_13),
.A2(n_271),
.B1(n_279),
.B2(n_300),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_13),
.A2(n_227),
.B1(n_279),
.B2(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_13),
.A2(n_279),
.B1(n_386),
.B2(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_14),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_15),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_15),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_15),
.A2(n_80),
.B1(n_181),
.B2(n_185),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_15),
.A2(n_80),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_43),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_16),
.A2(n_36),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_234),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_232),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_208),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_20),
.B(n_208),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_128),
.C(n_177),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_21),
.A2(n_22),
.B1(n_128),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_90),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_23),
.A2(n_24),
.B(n_92),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_47),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_91),
.B1(n_92),
.B2(n_127),
.Y(n_90)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_24),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_24),
.A2(n_47),
.B1(n_127),
.B2(n_428),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_25),
.A2(n_35),
.B1(n_180),
.B2(n_187),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_25),
.A2(n_263),
.B(n_268),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_25),
.A2(n_249),
.B(n_268),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_25),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_397)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_26),
.B(n_270),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_26),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_26),
.A2(n_340),
.B1(n_371),
.B2(n_374),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_26),
.A2(n_374),
.B1(n_401),
.B2(n_434),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_27),
.Y(n_304)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_28),
.Y(n_188)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_28),
.Y(n_375)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_29),
.Y(n_274)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_31),
.Y(n_344)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_31),
.Y(n_372)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_40),
.Y(n_186)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_41),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_42),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_42),
.Y(n_273)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_45),
.Y(n_267)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_46),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_47),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_57),
.B1(n_79),
.B2(n_89),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_48),
.A2(n_57),
.B1(n_89),
.B2(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_52),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_52),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_52),
.Y(n_174)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_53),
.Y(n_175)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g352 ( 
.A(n_54),
.B(n_353),
.Y(n_352)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_56),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_56),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_56),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_56),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_57),
.A2(n_79),
.B1(n_89),
.B2(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_57),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_57),
.B(n_251),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_68),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_59),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_67),
.Y(n_349)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_68),
.A2(n_278),
.B(n_283),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_89),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_89),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_113),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_94),
.Y(n_213)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_101),
.B(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_101),
.Y(n_214)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_105),
.Y(n_391)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_108),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_108),
.Y(n_332)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_113),
.A2(n_214),
.B(n_437),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_120),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_121),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_121),
.A2(n_409),
.B(n_411),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_123),
.Y(n_389)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx8_ASAP7_75t_L g410 ( 
.A(n_124),
.Y(n_410)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_128),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_170),
.B(n_176),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_171),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_145),
.B1(n_153),
.B2(n_162),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_131),
.A2(n_326),
.B(n_333),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_131),
.B(n_367),
.Y(n_366)
);

AOI22x1_ASAP7_75t_L g440 ( 
.A1(n_131),
.A2(n_145),
.B1(n_367),
.B2(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_131),
.A2(n_333),
.B(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_132),
.A2(n_154),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_132),
.A2(n_200),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_132),
.A2(n_200),
.B1(n_364),
.B2(n_414),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_145),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_136),
.B1(n_140),
.B2(n_143),
.Y(n_133)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_134),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_136),
.Y(n_335)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_139),
.Y(n_327)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_139),
.Y(n_385)
);

AO22x2_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_146),
.B1(n_149),
.B2(n_151),
.Y(n_145)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_142),
.Y(n_351)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_169),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_173),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_209),
.CI(n_210),
.CON(n_208),
.SN(n_208)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_177),
.B(n_443),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_196),
.C(n_201),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_178),
.B(n_426),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_179),
.B(n_189),
.Y(n_451)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_180),
.Y(n_434)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_184),
.Y(n_293)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_184),
.Y(n_342)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_185),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_187),
.Y(n_312)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_190),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_196),
.B(n_201),
.Y(n_426)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_197),
.Y(n_441)
);

AOI32xp33_ASAP7_75t_L g346 ( 
.A1(n_198),
.A2(n_329),
.A3(n_347),
.B1(n_350),
.B2(n_352),
.Y(n_346)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_200),
.B(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_200),
.A2(n_364),
.B(n_366),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B(n_207),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_202),
.A2(n_203),
.B1(n_214),
.B2(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_207),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g484 ( 
.A(n_208),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_217),
.B2(n_231),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_214),
.B(n_249),
.Y(n_369)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_230),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_243),
.B(n_250),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_219),
.A2(n_220),
.B1(n_278),
.B2(n_323),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_219),
.A2(n_250),
.B(n_323),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_219),
.A2(n_220),
.B1(n_417),
.B2(n_432),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_220),
.A2(n_283),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_225),
.B(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_228),
.Y(n_336)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI311xp33_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_422),
.A3(n_459),
.B1(n_477),
.C1(n_478),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_378),
.B(n_421),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_355),
.B(n_377),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_317),
.B(n_354),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_286),
.B(n_316),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_261),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_241),
.B(n_261),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_253),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_242),
.A2(n_253),
.B1(n_254),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_249),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_249),
.B(n_393),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_SL g409 ( 
.A1(n_249),
.A2(n_392),
.B(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_275),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_276),
.C(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_266),
.Y(n_373)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_273),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_284),
.B2(n_285),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_308),
.B(n_315),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_297),
.B(n_307),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_294),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_306),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_306),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_303),
.B(n_305),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_339),
.B(n_345),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_313),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_319),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_337),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_324),
.C(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx6_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_334),
.Y(n_367)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_346),
.Y(n_361)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx5_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_356),
.B(n_357),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_362),
.B2(n_376),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_361),
.C(n_376),
.Y(n_379)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_368),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_369),
.C(n_370),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_379),
.B(n_380),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_406),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_381)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_396),
.B2(n_397),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_384),
.B(n_396),
.Y(n_455)
);

OAI32xp33_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.A3(n_388),
.B1(n_390),
.B2(n_392),
.Y(n_384)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_403),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_403),
.B(n_404),
.C(n_406),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_412),
.B2(n_420),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_407),
.B(n_413),
.C(n_416),
.Y(n_468)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_412),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_414),
.Y(n_457)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_445),
.Y(n_422)
);

A2O1A1Ixp33_ASAP7_75t_SL g478 ( 
.A1(n_423),
.A2(n_445),
.B(n_479),
.C(n_482),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_442),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_442),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_427),
.C(n_429),
.Y(n_424)
);

FAx1_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_427),
.CI(n_429),
.CON(n_458),
.SN(n_458)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_435),
.C(n_440),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_433),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_435),
.A2(n_436),
.B1(n_440),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_440),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_458),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_458),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.C(n_452),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_448),
.B1(n_451),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.C(n_456),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_453),
.A2(n_454),
.B1(n_456),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_472),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_480),
.B(n_481),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_469),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_469),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.C(n_468),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_475),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_467),
.B1(n_468),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_474),
.Y(n_480)
);


endmodule