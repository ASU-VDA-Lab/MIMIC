module fake_jpeg_27430_n_169 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_1),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_21),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_15),
.B1(n_26),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_77)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_38),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_32),
.B1(n_48),
.B2(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_67),
.B1(n_56),
.B2(n_49),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_14),
.B(n_28),
.C(n_27),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_3),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_41),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_65),
.Y(n_101)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_76),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_23),
.B1(n_18),
.B2(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_84),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_40),
.B1(n_21),
.B2(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_16),
.B1(n_22),
.B2(n_5),
.Y(n_87)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_52),
.B(n_43),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_105),
.B(n_80),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_43),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_104),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_58),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_3),
.B(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_64),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_81),
.B1(n_83),
.B2(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_115),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_112),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_119),
.B(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_69),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_120),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_122),
.B(n_123),
.Y(n_134)
);

HAxp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_63),
.CON(n_119),
.SN(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_131),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_98),
.C(n_104),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_117),
.C(n_112),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_96),
.B(n_107),
.C(n_106),
.D(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_113),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_131),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_142),
.C(n_134),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_122),
.B1(n_110),
.B2(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_141),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_88),
.B1(n_118),
.B2(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_114),
.C(n_97),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_111),
.C(n_69),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_78),
.C(n_76),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_151),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

OAI322xp33_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_129),
.A3(n_128),
.B1(n_111),
.B2(n_92),
.C1(n_8),
.C2(n_9),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_78),
.C(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_136),
.B1(n_140),
.B2(n_144),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_146),
.B(n_8),
.Y(n_159)
);

NAND4xp25_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_148),
.C(n_9),
.D(n_11),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_159),
.A2(n_161),
.B1(n_12),
.B2(n_4),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_72),
.B1(n_7),
.B2(n_11),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_155),
.B(n_161),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_157),
.B(n_6),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_163),
.B(n_3),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_166),
.B(n_164),
.C(n_157),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_6),
.Y(n_169)
);


endmodule