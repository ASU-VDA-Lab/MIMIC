module fake_ariane_1296_n_198 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_198);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_198;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_194;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_10),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_R g55 ( 
.A(n_49),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_R g61 ( 
.A(n_34),
.B(n_19),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_R g65 ( 
.A(n_33),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_R g67 ( 
.A(n_38),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_0),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_39),
.B(n_0),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_R g73 ( 
.A(n_43),
.B(n_2),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_52),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_52),
.B(n_50),
.C(n_40),
.Y(n_78)
);

NAND2x1p5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_47),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_42),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_72),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_71),
.B1(n_75),
.B2(n_68),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_60),
.B(n_69),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_44),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_37),
.B(n_40),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_85),
.B(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_41),
.Y(n_100)
);

OR2x6_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_73),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_73),
.B1(n_55),
.B2(n_65),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_55),
.B1(n_65),
.B2(n_67),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_79),
.B(n_91),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_79),
.B(n_91),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_79),
.B(n_89),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_89),
.B(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_96),
.B1(n_99),
.B2(n_93),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_84),
.B(n_86),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

OR2x6_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_104),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_103),
.B1(n_101),
.B2(n_90),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_R g118 ( 
.A(n_109),
.B(n_83),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_117),
.A2(n_90),
.B(n_5),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AND2x4_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_107),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_108),
.B1(n_77),
.B2(n_112),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

NAND2x1p5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_114),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_107),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_115),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_114),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_105),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_127),
.Y(n_145)
);

NOR4xp25_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_118),
.C(n_128),
.D(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_127),
.B1(n_77),
.B2(n_129),
.C(n_128),
.Y(n_148)
);

OAI31xp33_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_129),
.A3(n_76),
.B(n_134),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_133),
.B(n_61),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_142),
.B(n_141),
.Y(n_151)
);

NAND2x1p5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_141),
.B(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_142),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_142),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_76),
.CON(n_158),
.SN(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_148),
.C(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_157),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_140),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_154),
.B1(n_153),
.B2(n_157),
.C(n_158),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_R g166 ( 
.A(n_160),
.B(n_140),
.Y(n_166)
);

NAND5xp2_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_152),
.C(n_141),
.D(n_108),
.E(n_112),
.Y(n_167)
);

OAI222xp33_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_130),
.B1(n_135),
.B2(n_152),
.C1(n_142),
.C2(n_125),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_140),
.Y(n_169)
);

NAND4xp75_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_142),
.C(n_141),
.D(n_152),
.Y(n_170)
);

AOI222xp33_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_159),
.B1(n_138),
.B2(n_140),
.C1(n_139),
.C2(n_8),
.Y(n_171)
);

OAI211xp5_ASAP7_75t_SL g172 ( 
.A1(n_169),
.A2(n_159),
.B(n_140),
.C(n_139),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_159),
.B(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_140),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_140),
.B1(n_139),
.B2(n_135),
.Y(n_176)
);

AOI222xp33_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_162),
.B1(n_138),
.B2(n_170),
.C1(n_140),
.C2(n_139),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_139),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_139),
.C(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

AND3x1_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_173),
.C(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_177),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

AOI211x1_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_180),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_180),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_105),
.C(n_138),
.Y(n_188)
);

NAND4xp25_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_4),
.C(n_6),
.D(n_7),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

OAI221xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_130),
.B1(n_9),
.B2(n_12),
.C(n_13),
.Y(n_192)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_138),
.B1(n_9),
.B2(n_13),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_7),
.Y(n_194)
);

AOI211xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_190),
.B(n_192),
.C(n_188),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_187),
.B1(n_186),
.B2(n_138),
.Y(n_197)
);

NAND4xp25_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_195),
.C(n_14),
.D(n_16),
.Y(n_198)
);


endmodule