module fake_jpeg_4244_n_11 (n_3, n_2, n_1, n_0, n_4, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

OA22x2_ASAP7_75t_L g5 ( 
.A1(n_1),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_5)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_2),
.B(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_5),
.C(n_7),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_9),
.A2(n_5),
.B1(n_6),
.B2(n_3),
.Y(n_10)
);

XNOR2x2_ASAP7_75t_SL g11 ( 
.A(n_10),
.B(n_3),
.Y(n_11)
);


endmodule