module fake_aes_10717_n_38 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
OA21x2_ASAP7_75t_L g15 ( .A1(n_0), .A2(n_3), .B(n_6), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_10), .Y(n_17) );
O2A1O1Ixp33_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_0), .B(n_1), .C(n_2), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_14), .B(n_3), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g20 ( .A(n_17), .B(n_7), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_14), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_16), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_16), .Y(n_23) );
NOR2xp67_ASAP7_75t_L g24 ( .A(n_22), .B(n_19), .Y(n_24) );
OAI22xp33_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_13), .B1(n_12), .B2(n_15), .Y(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_23), .B1(n_18), .B2(n_20), .C(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_26), .B(n_15), .Y(n_28) );
NOR3xp33_ASAP7_75t_SL g29 ( .A(n_27), .B(n_15), .C(n_5), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_4), .Y(n_30) );
NAND3xp33_ASAP7_75t_SL g31 ( .A(n_29), .B(n_15), .C(n_5), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_28), .B(n_4), .Y(n_32) );
AND2x4_ASAP7_75t_SL g33 ( .A(n_31), .B(n_11), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_35), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_33), .B1(n_36), .B2(n_31), .Y(n_38) );
endmodule