module fake_jpeg_9523_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_21),
.B1(n_26),
.B2(n_18),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_19),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_21),
.B1(n_14),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_22),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_60),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_29),
.B1(n_19),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_76),
.B1(n_65),
.B2(n_26),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_66),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_16),
.B(n_27),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_17),
.B(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_70),
.Y(n_99)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_39),
.B(n_25),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_91),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_34),
.B(n_1),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_35),
.A3(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_3),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_92),
.B(n_24),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_50),
.B(n_31),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_75),
.B1(n_60),
.B2(n_71),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_98),
.B1(n_73),
.B2(n_75),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_58),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_42),
.B1(n_38),
.B2(n_44),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_97),
.B1(n_64),
.B2(n_1),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_42),
.B1(n_38),
.B2(n_44),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_38),
.B1(n_24),
.B2(n_23),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_55),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_104),
.C(n_112),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_55),
.B1(n_75),
.B2(n_63),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_106),
.B(n_107),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_119),
.B1(n_122),
.B2(n_88),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_69),
.C(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_23),
.B1(n_20),
.B2(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_0),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_117),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_35),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_115),
.B1(n_90),
.B2(n_79),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_64),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_0),
.C(n_2),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_87),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_86),
.B1(n_83),
.B2(n_81),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_133),
.B1(n_135),
.B2(n_137),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_128),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_88),
.B1(n_84),
.B2(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_79),
.B1(n_85),
.B2(n_89),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_85),
.B1(n_95),
.B2(n_89),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_107),
.B1(n_113),
.B2(n_121),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_93),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_135),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_158),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_115),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_153),
.C(n_156),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_95),
.B(n_93),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_151),
.B(n_126),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_138),
.B1(n_134),
.B2(n_128),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_3),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_4),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_4),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_140),
.C(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_164),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_142),
.C(n_129),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_165),
.C(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_155),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_124),
.C(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_148),
.B(n_144),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_175),
.B(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_173),
.B(n_175),
.Y(n_184)
);

AOI31xp67_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_127),
.A3(n_157),
.B(n_138),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_165),
.C(n_162),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_4),
.C(n_6),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_187),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_158),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_178),
.C(n_174),
.Y(n_186)
);

OAI21x1_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_9),
.B(n_10),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_9),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_8),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_188),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_8),
.B(n_9),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_192),
.A2(n_11),
.B(n_12),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_193),
.A2(n_183),
.B(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_198),
.B(n_191),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_189),
.B(n_194),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_200),
.B(n_11),
.Y(n_203)
);


endmodule