module real_jpeg_23254_n_16 (n_5, n_4, n_8, n_0, n_12, n_345, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_345;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_66),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_47),
.C(n_50),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_132),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_4),
.B(n_30),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_104),
.B1(n_207),
.B2(n_210),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_59),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_6),
.A2(n_42),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_6),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_7),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_127),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_127),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_127),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_9),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_9),
.A2(n_26),
.B1(n_58),
.B2(n_65),
.Y(n_293)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_29),
.C(n_63),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_68),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_12),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_129),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_129),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_12),
.A2(n_58),
.B1(n_65),
.B2(n_129),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_13),
.A2(n_57),
.B1(n_75),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_136),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_136),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_136),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_15),
.Y(n_107)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_78),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_20),
.A2(n_72),
.B1(n_328),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_20),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_22),
.B(n_44),
.C(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_24),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_25),
.A2(n_30),
.B(n_38),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_25),
.A2(n_38),
.B(n_81),
.Y(n_273)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_27),
.A2(n_62),
.B(n_133),
.C(n_153),
.Y(n_152)
);

HAxp5_ASAP7_75t_SL g224 ( 
.A(n_27),
.B(n_132),
.CON(n_224),
.SN(n_224)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g225 ( 
.A(n_29),
.B(n_32),
.C(n_34),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_30),
.A2(n_38),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_30),
.A2(n_38),
.B1(n_167),
.B2(n_224),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_30),
.A2(n_38),
.B1(n_80),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_31),
.A2(n_146),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_31),
.A2(n_37),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_31)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_33),
.A2(n_36),
.B(n_223),
.C(n_225),
.Y(n_222)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_34),
.B(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_38),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_38),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_72),
.C(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_43),
.A2(n_44),
.B1(n_79),
.B2(n_331),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_45),
.A2(n_49),
.B1(n_182),
.B2(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_45),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_45),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_49),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_49),
.B(n_121),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_49),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_49),
.B(n_132),
.Y(n_205)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_51),
.B(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_53),
.A2(n_119),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_53),
.B(n_180),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_66),
.B2(n_67),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_61),
.B(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_67),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_60),
.A2(n_66),
.B1(n_131),
.B2(n_134),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_60),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_60),
.A2(n_66),
.B1(n_143),
.B2(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_61),
.A2(n_135),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_66),
.B(n_293),
.Y(n_292)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_72),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_72),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_75),
.B(n_132),
.Y(n_133)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_78),
.B(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_79),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_88),
.A2(n_141),
.B(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_325),
.A3(n_337),
.B1(n_342),
.B2(n_343),
.C(n_345),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_302),
.B(n_324),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_276),
.B(n_301),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_169),
.B(n_257),
.C(n_275),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_155),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_100),
.B(n_155),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_137),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_122),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_102),
.B(n_122),
.C(n_137),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_116),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_103),
.B(n_116),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.B(n_110),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_104),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_104),
.A2(n_113),
.B1(n_200),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_104),
.A2(n_110),
.B(n_189),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_104),
.A2(n_189),
.B(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_109),
.B1(n_112),
.B2(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_105),
.B(n_111),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_105),
.A2(n_112),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_151),
.B(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_115),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_117),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_118),
.B(n_247),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_119),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_119),
.A2(n_180),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_119),
.A2(n_180),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.C(n_130),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_125),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_124),
.Y(n_285)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_132),
.B(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_147),
.B2(n_154),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_140),
.B(n_144),
.C(n_154),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_141),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_156),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_158),
.B(n_160),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_165),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_162),
.B(n_186),
.Y(n_263)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_165),
.B(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_256),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_251),
.B(n_255),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_235),
.B(n_250),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_218),
.B(n_234),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_196),
.B(n_217),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_183),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_183),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_178),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_191),
.C(n_194),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_203),
.B(n_216),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_202),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_208),
.B(n_215),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_233),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_233),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_229),
.C(n_230),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_237),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_245),
.C(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_254),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_259),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_274),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_268),
.C(n_274),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_267),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_267),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_271),
.C(n_273),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_277),
.B(n_278),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_300),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_287),
.B1(n_298),
.B2(n_299),
.Y(n_279)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_299),
.C(n_300),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_286),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_281),
.A2(n_282),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_281),
.A2(n_312),
.B(n_316),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_283),
.Y(n_313)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_294),
.C(n_297),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_294),
.B1(n_295),
.B2(n_297),
.Y(n_289)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_293),
.Y(n_317)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_303),
.B(n_304),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_304)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_311),
.B1(n_319),
.B2(n_320),
.Y(n_305)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_309),
.B(n_310),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_307),
.B(n_309),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_310),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_327),
.B1(n_332),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_319),
.C(n_323),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_321),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_334),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_334),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_332),
.C(n_333),
.Y(n_326)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_338),
.B(n_339),
.Y(n_342)
);


endmodule