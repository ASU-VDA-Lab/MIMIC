module real_aes_16614_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g103 ( .A(n_0), .B(n_104), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_1), .A2(n_4), .B1(n_251), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_2), .A2(n_41), .B1(n_146), .B2(n_148), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_3), .A2(n_22), .B1(n_148), .B2(n_191), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_5), .A2(n_15), .B1(n_173), .B2(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_6), .A2(n_58), .B1(n_193), .B2(n_218), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_7), .A2(n_16), .B1(n_146), .B2(n_177), .Y(n_607) );
INVx1_ASAP7_75t_L g104 ( .A(n_8), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_9), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_10), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_11), .A2(n_17), .B1(n_175), .B2(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
OR2x2_ASAP7_75t_L g120 ( .A(n_12), .B(n_37), .Y(n_120) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_13), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_14), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_18), .A2(n_97), .B1(n_173), .B2(n_251), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_19), .A2(n_38), .B1(n_209), .B2(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_20), .B(n_174), .Y(n_206) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_21), .A2(n_55), .B(n_163), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_23), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_24), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_25), .B(n_152), .Y(n_515) );
INVx4_ASAP7_75t_R g570 ( .A(n_26), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_27), .A2(n_45), .B1(n_154), .B2(n_156), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_28), .A2(n_100), .B1(n_112), .B2(n_857), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_29), .A2(n_51), .B1(n_156), .B2(n_173), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_30), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_31), .B(n_209), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_32), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_33), .B(n_148), .Y(n_522) );
INVx1_ASAP7_75t_L g531 ( .A(n_34), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_SL g588 ( .A1(n_35), .A2(n_146), .B(n_158), .C(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_36), .A2(n_52), .B1(n_146), .B2(n_156), .Y(n_504) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_37), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_39), .A2(n_83), .B1(n_146), .B2(n_190), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_40), .A2(n_44), .B1(n_146), .B2(n_177), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_42), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_43), .A2(n_57), .B1(n_173), .B2(n_228), .Y(n_253) );
INVx1_ASAP7_75t_L g519 ( .A(n_46), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_47), .B(n_146), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_48), .Y(n_540) );
INVx2_ASAP7_75t_L g126 ( .A(n_49), .Y(n_126) );
BUFx3_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
INVx1_ASAP7_75t_L g118 ( .A(n_50), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_53), .A2(n_130), .B1(n_836), .B2(n_837), .Y(n_129) );
INVx1_ASAP7_75t_L g836 ( .A(n_53), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_54), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_56), .A2(n_85), .B1(n_146), .B2(n_156), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_59), .A2(n_72), .B1(n_154), .B2(n_228), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_60), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_61), .A2(n_74), .B1(n_146), .B2(n_177), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_62), .A2(n_95), .B1(n_173), .B2(n_175), .Y(n_172) );
AND2x4_ASAP7_75t_L g142 ( .A(n_63), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g163 ( .A(n_64), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_65), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_66), .A2(n_88), .B1(n_154), .B2(n_156), .Y(n_527) );
AO22x1_ASAP7_75t_L g557 ( .A1(n_67), .A2(n_73), .B1(n_239), .B2(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g143 ( .A(n_68), .Y(n_143) );
AND2x2_ASAP7_75t_L g591 ( .A(n_69), .B(n_160), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_70), .B(n_193), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_71), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_75), .B(n_148), .Y(n_541) );
INVx2_ASAP7_75t_L g152 ( .A(n_76), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_77), .B(n_160), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_78), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_79), .A2(n_96), .B1(n_156), .B2(n_193), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_80), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_81), .B(n_170), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_82), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_84), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_86), .A2(n_131), .B1(n_844), .B2(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_86), .Y(n_844) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_87), .B(n_160), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_89), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_90), .B(n_160), .Y(n_537) );
INVx1_ASAP7_75t_L g106 ( .A(n_91), .Y(n_106) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_92), .B(n_174), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_93), .A2(n_179), .B(n_193), .C(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g572 ( .A(n_94), .B(n_573), .Y(n_572) );
NAND2xp33_ASAP7_75t_L g545 ( .A(n_98), .B(n_155), .Y(n_545) );
AND2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_108), .Y(n_100) );
AND2x4_ASAP7_75t_L g858 ( .A(n_101), .B(n_108), .Y(n_858) );
NOR3x1_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .C(n_107), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
AND3x2_ASAP7_75t_L g116 ( .A(n_105), .B(n_117), .C(n_119), .Y(n_116) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g490 ( .A(n_106), .Y(n_490) );
INVx1_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
NOR2x1_ASAP7_75t_L g856 ( .A(n_107), .B(n_120), .Y(n_856) );
NOR2x1p5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_121), .Y(n_112) );
INVxp67_ASAP7_75t_SL g846 ( .A(n_113), .Y(n_846) );
NOR2x1_ASAP7_75t_R g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx3_ASAP7_75t_L g842 ( .A(n_115), .Y(n_842) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_119), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_129), .B(n_838), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
BUFx12f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_SL g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx3_ASAP7_75t_L g848 ( .A(n_125), .Y(n_848) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_126), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g837 ( .A(n_130), .Y(n_837) );
OA22x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_487), .B1(n_491), .B2(n_493), .Y(n_130) );
INVx2_ASAP7_75t_L g845 ( .A(n_131), .Y(n_845) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_383), .Y(n_131) );
NOR2x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_335), .Y(n_132) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_282), .C(n_320), .Y(n_133) );
AOI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_213), .B1(n_233), .B2(n_261), .C(n_267), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_135), .A2(n_460), .B1(n_463), .B2(n_464), .Y(n_459) );
INVx2_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_184), .Y(n_136) );
INVx1_ASAP7_75t_L g374 ( .A(n_137), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_166), .Y(n_137) );
INVx1_ASAP7_75t_L g326 ( .A(n_138), .Y(n_326) );
AND2x4_ASAP7_75t_L g369 ( .A(n_138), .B(n_290), .Y(n_369) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g297 ( .A(n_139), .B(n_200), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_139), .B(n_266), .Y(n_357) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g265 ( .A(n_140), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g281 ( .A(n_140), .B(n_186), .Y(n_281) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_140), .Y(n_288) );
INVx1_ASAP7_75t_L g344 ( .A(n_140), .Y(n_344) );
AO31x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .A3(n_159), .B(n_164), .Y(n_140) );
INVx2_ASAP7_75t_L g181 ( .A(n_141), .Y(n_181) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_141), .A2(n_168), .A3(n_215), .B(n_221), .Y(n_214) );
AO31x2_ASAP7_75t_L g236 ( .A1(n_141), .A2(n_187), .A3(n_237), .B(n_244), .Y(n_236) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_141), .A2(n_232), .A3(n_606), .B(n_609), .Y(n_605) );
BUFx10_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
BUFx10_ASAP7_75t_L g506 ( .A(n_142), .Y(n_506) );
INVx1_ASAP7_75t_L g561 ( .A(n_142), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B1(n_153), .B2(n_157), .Y(n_144) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
INVx4_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
INVx1_ASAP7_75t_L g228 ( .A(n_146), .Y(n_228) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_147), .Y(n_148) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
INVx2_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
INVx1_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
INVx1_ASAP7_75t_L g219 ( .A(n_147), .Y(n_219) );
INVx1_ASAP7_75t_L g240 ( .A(n_147), .Y(n_240) );
INVx1_ASAP7_75t_L g243 ( .A(n_147), .Y(n_243) );
INVx1_ASAP7_75t_L g252 ( .A(n_147), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_148), .B(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_149), .A2(n_157), .B1(n_227), .B2(n_229), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_149), .A2(n_157), .B1(n_238), .B2(n_241), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_149), .A2(n_157), .B1(n_250), .B2(n_253), .Y(n_249) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g505 ( .A(n_150), .Y(n_505) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g543 ( .A(n_151), .Y(n_543) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx8_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx1_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
INVx1_ASAP7_75t_L g518 ( .A(n_152), .Y(n_518) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_155), .A2(n_243), .B1(n_570), .B2(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_156), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g529 ( .A(n_156), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_157), .A2(n_172), .B1(n_176), .B2(n_178), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_157), .A2(n_189), .B1(n_192), .B2(n_194), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_157), .A2(n_208), .B(n_210), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_157), .A2(n_178), .B1(n_216), .B2(n_220), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_157), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_157), .A2(n_194), .B1(n_527), .B2(n_528), .Y(n_526) );
OAI22x1_ASAP7_75t_L g606 ( .A1(n_157), .A2(n_194), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx6_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
O2A1O1Ixp5_ASAP7_75t_L g204 ( .A1(n_158), .A2(n_177), .B(n_205), .C(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_158), .A2(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_158), .B(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_158), .A2(n_553), .B(n_557), .C(n_560), .Y(n_619) );
AO31x2_ASAP7_75t_L g501 ( .A1(n_159), .A2(n_502), .A3(n_506), .B(n_507), .Y(n_501) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_160), .B(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_161), .B(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_161), .B(n_183), .Y(n_182) );
BUFx3_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
INVx2_ASAP7_75t_SL g202 ( .A(n_161), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_161), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g523 ( .A(n_161), .B(n_506), .Y(n_523) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g170 ( .A(n_162), .Y(n_170) );
INVx3_ASAP7_75t_L g264 ( .A(n_166), .Y(n_264) );
AND2x2_ASAP7_75t_L g279 ( .A(n_166), .B(n_200), .Y(n_279) );
INVx2_ASAP7_75t_L g285 ( .A(n_166), .Y(n_285) );
AND2x4_ASAP7_75t_L g347 ( .A(n_166), .B(n_186), .Y(n_347) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_166), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_166), .B(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g296 ( .A(n_167), .B(n_186), .Y(n_296) );
AND2x2_ASAP7_75t_L g324 ( .A(n_167), .B(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g403 ( .A(n_167), .Y(n_403) );
AO31x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .A3(n_180), .B(n_182), .Y(n_167) );
AO31x2_ASAP7_75t_L g525 ( .A1(n_168), .A2(n_195), .A3(n_526), .B(n_530), .Y(n_525) );
AOI21x1_ASAP7_75t_L g580 ( .A1(n_168), .A2(n_581), .B(n_591), .Y(n_580) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_169), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_169), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g573 ( .A(n_169), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_169), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g198 ( .A(n_170), .Y(n_198) );
INVx2_ASAP7_75t_L g232 ( .A(n_170), .Y(n_232) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_170), .A2(n_555), .B(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_174), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_177), .A2(n_540), .B(n_541), .C(n_542), .Y(n_539) );
INVx1_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_180), .A2(n_224), .A3(n_249), .B(n_254), .Y(n_248) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_181), .A2(n_565), .B(n_568), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
INVx1_ASAP7_75t_L g359 ( .A(n_185), .Y(n_359) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_185), .B(n_279), .Y(n_387) );
BUFx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g289 ( .A(n_186), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g325 ( .A(n_186), .Y(n_325) );
INVx1_ASAP7_75t_L g401 ( .A(n_186), .Y(n_401) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .A3(n_195), .B(n_197), .Y(n_186) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_191), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_194), .B(n_569), .Y(n_568) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_195), .A2(n_224), .A3(n_226), .B(n_230), .Y(n_223) );
INVx2_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_SL g211 ( .A(n_196), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g221 ( .A(n_198), .B(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g225 ( .A(n_198), .Y(n_225) );
AND2x4_ASAP7_75t_L g340 ( .A(n_200), .B(n_325), .Y(n_340) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g362 ( .A(n_201), .Y(n_362) );
OAI21x1_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_212), .Y(n_201) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_202), .A2(n_203), .B(n_212), .Y(n_266) );
OAI21x1_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_207), .B(n_211), .Y(n_203) );
AND2x4_ASAP7_75t_L g234 ( .A(n_213), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_223), .Y(n_213) );
INVx4_ASAP7_75t_SL g258 ( .A(n_214), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_214), .B(n_260), .Y(n_270) );
BUFx2_ASAP7_75t_L g334 ( .A(n_214), .Y(n_334) );
AND2x2_ASAP7_75t_L g378 ( .A(n_214), .B(n_236), .Y(n_378) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_219), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
OR2x2_ASAP7_75t_L g294 ( .A(n_223), .B(n_236), .Y(n_294) );
INVx2_ASAP7_75t_L g305 ( .A(n_223), .Y(n_305) );
AND2x4_ASAP7_75t_L g308 ( .A(n_223), .B(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_223), .Y(n_349) );
INVx1_ASAP7_75t_L g390 ( .A(n_223), .Y(n_390) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_224), .A2(n_564), .B(n_572), .Y(n_563) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_232), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_246), .Y(n_233) );
INVx2_ASAP7_75t_L g483 ( .A(n_234), .Y(n_483) );
AND2x4_ASAP7_75t_L g444 ( .A(n_235), .B(n_247), .Y(n_444) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx2_ASAP7_75t_L g309 ( .A(n_236), .Y(n_309) );
INVx1_ASAP7_75t_L g365 ( .A(n_236), .Y(n_365) );
AND2x2_ASAP7_75t_L g391 ( .A(n_236), .B(n_316), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_236), .B(n_304), .Y(n_395) );
OAI21xp33_ASAP7_75t_SL g514 ( .A1(n_239), .A2(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_257), .Y(n_246) );
INVx3_ASAP7_75t_L g372 ( .A(n_247), .Y(n_372) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_256), .Y(n_247) );
INVx2_ASAP7_75t_L g276 ( .A(n_248), .Y(n_276) );
INVx2_ASAP7_75t_L g316 ( .A(n_248), .Y(n_316) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_252), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_256), .B(n_258), .Y(n_317) );
AND2x2_ASAP7_75t_L g345 ( .A(n_256), .B(n_316), .Y(n_345) );
INVx1_ASAP7_75t_L g271 ( .A(n_257), .Y(n_271) );
NAND2x1_ASAP7_75t_L g407 ( .A(n_257), .B(n_381), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_257), .B(n_345), .Y(n_456) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g274 ( .A(n_258), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_258), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g364 ( .A(n_258), .B(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_258), .Y(n_441) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_261), .A2(n_454), .B1(n_455), .B2(n_457), .Y(n_453) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_263), .B(n_297), .Y(n_332) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g355 ( .A(n_264), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g454 ( .A(n_264), .B(n_265), .Y(n_454) );
AND2x2_ASAP7_75t_L g327 ( .A(n_265), .B(n_296), .Y(n_327) );
AND2x4_ASAP7_75t_L g346 ( .A(n_265), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g397 ( .A(n_265), .B(n_324), .Y(n_397) );
INVx1_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
AOI31xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .A3(n_272), .B(n_277), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_269), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_269), .Y(n_463) );
OAI21xp33_ASAP7_75t_L g481 ( .A1(n_269), .A2(n_271), .B(n_301), .Y(n_481) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g323 ( .A(n_270), .Y(n_323) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g458 ( .A(n_273), .B(n_294), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g292 ( .A(n_274), .Y(n_292) );
INVx1_ASAP7_75t_L g313 ( .A(n_275), .Y(n_313) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_275), .Y(n_420) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g302 ( .A(n_276), .Y(n_302) );
OR2x2_ASAP7_75t_L g330 ( .A(n_276), .B(n_305), .Y(n_330) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2x1p5_ASAP7_75t_L g319 ( .A(n_281), .B(n_285), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_291), .B1(n_295), .B2(n_298), .C(n_310), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2x1_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g399 ( .A(n_288), .B(n_302), .Y(n_399) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OR2x2_ASAP7_75t_L g329 ( .A(n_292), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g416 ( .A(n_292), .B(n_308), .Y(n_416) );
AND2x4_ASAP7_75t_L g333 ( .A(n_293), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g352 ( .A(n_294), .B(n_315), .Y(n_352) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_296), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g409 ( .A(n_296), .Y(n_409) );
INVx2_ASAP7_75t_L g418 ( .A(n_296), .Y(n_418) );
AND2x2_ASAP7_75t_L g432 ( .A(n_296), .B(n_362), .Y(n_432) );
INVx1_ASAP7_75t_L g410 ( .A(n_297), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_306), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_300), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_301), .B(n_308), .Y(n_342) );
AND2x2_ASAP7_75t_L g363 ( .A(n_301), .B(n_364), .Y(n_363) );
NAND2x1_ASAP7_75t_L g471 ( .A(n_301), .B(n_333), .Y(n_471) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B(n_318), .Y(n_310) );
NAND2x1_ASAP7_75t_L g472 ( .A(n_312), .B(n_416), .Y(n_472) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_313), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx4_ASAP7_75t_L g381 ( .A(n_315), .Y(n_381) );
AND2x2_ASAP7_75t_L g451 ( .A(n_315), .B(n_356), .Y(n_451) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g348 ( .A(n_316), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g361 ( .A(n_319), .B(n_362), .Y(n_361) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_319), .B(n_432), .Y(n_431) );
AOI322xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .A3(n_326), .B1(n_327), .B2(n_328), .C1(n_331), .C2(n_333), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g414 ( .A(n_324), .B(n_362), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_324), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g438 ( .A(n_324), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g443 ( .A(n_324), .B(n_428), .Y(n_443) );
INVx1_ASAP7_75t_L g452 ( .A(n_324), .Y(n_452) );
OR2x2_ASAP7_75t_L g338 ( .A(n_326), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g465 ( .A(n_326), .Y(n_465) );
AND2x2_ASAP7_75t_L g468 ( .A(n_327), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR3xp33_ASAP7_75t_L g404 ( .A(n_330), .B(n_344), .C(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g446 ( .A(n_330), .Y(n_446) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND3xp33_ASAP7_75t_SL g335 ( .A(n_336), .B(n_350), .C(n_360), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B1(n_343), .B2(n_345), .C1(n_346), .C2(n_348), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22x1_ASAP7_75t_L g482 ( .A1(n_339), .A2(n_483), .B1(n_484), .B2(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g343 ( .A(n_340), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_340), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g436 ( .A(n_340), .B(n_402), .Y(n_436) );
AND2x4_ASAP7_75t_L g466 ( .A(n_340), .B(n_403), .Y(n_466) );
AND2x2_ASAP7_75t_L g447 ( .A(n_341), .B(n_414), .Y(n_447) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g439 ( .A(n_344), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_345), .B(n_378), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_345), .B(n_364), .Y(n_462) );
INVx1_ASAP7_75t_L g382 ( .A(n_346), .Y(n_382) );
INVx2_ASAP7_75t_L g426 ( .A(n_348), .Y(n_426) );
INVx1_ASAP7_75t_L g376 ( .A(n_349), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
AOI221xp5_ASAP7_75t_SL g442 ( .A1(n_355), .A2(n_443), .B1(n_444), .B2(n_445), .C(n_447), .Y(n_442) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g428 ( .A(n_357), .Y(n_428) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_357), .Y(n_480) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_359), .B(n_465), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B1(n_366), .B2(n_377), .C(n_379), .Y(n_360) );
OR2x2_ASAP7_75t_L g417 ( .A(n_362), .B(n_418), .Y(n_417) );
AOI32xp33_ASAP7_75t_L g398 ( .A1(n_364), .A2(n_378), .A3(n_399), .B1(n_400), .B2(n_404), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_364), .B(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B1(n_373), .B2(n_375), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_369), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g440 ( .A(n_372), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g433 ( .A(n_376), .B(n_378), .Y(n_433) );
AND2x2_ASAP7_75t_L g486 ( .A(n_376), .B(n_391), .Y(n_486) );
AND2x2_ASAP7_75t_L g445 ( .A(n_377), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_378), .B(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_448), .Y(n_383) );
NAND4xp75_ASAP7_75t_L g384 ( .A(n_385), .B(n_411), .C(n_429), .D(n_442), .Y(n_384) );
AOI211x1_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_392), .C(n_406), .Y(n_385) );
INVxp67_ASAP7_75t_L g484 ( .A(n_386), .Y(n_484) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B(n_398), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
BUFx2_ASAP7_75t_L g405 ( .A(n_401), .Y(n_405) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g477 ( .A(n_405), .Y(n_477) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .C(n_410), .Y(n_406) );
INVx2_ASAP7_75t_L g469 ( .A(n_407), .Y(n_469) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_421), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_417), .B2(n_419), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_426), .B2(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_434), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B(n_440), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_441), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g461 ( .A(n_444), .Y(n_461) );
NAND4xp75_ASAP7_75t_SL g448 ( .A(n_449), .B(n_459), .C(n_467), .D(n_475), .Y(n_448) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NOR2xp67_ASAP7_75t_SL g467 ( .A(n_468), .B(n_470), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_473), .Y(n_470) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
AOI21x1_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_481), .B(n_482), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx8_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
BUFx8_ASAP7_75t_SL g492 ( .A(n_490), .Y(n_492) );
AND2x2_ASAP7_75t_L g855 ( .A(n_490), .B(n_856), .Y(n_855) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_726), .Y(n_493) );
NOR4xp25_ASAP7_75t_L g494 ( .A(n_495), .B(n_626), .C(n_668), .D(n_700), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_532), .B(n_574), .C(n_611), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_509), .Y(n_498) );
INVx2_ASAP7_75t_L g639 ( .A(n_499), .Y(n_639) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g718 ( .A(n_500), .B(n_511), .Y(n_718) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_501), .B(n_525), .Y(n_577) );
AND2x2_ASAP7_75t_L g600 ( .A(n_501), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g625 ( .A(n_501), .Y(n_625) );
OR2x2_ASAP7_75t_L g688 ( .A(n_501), .B(n_525), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_505), .A2(n_521), .B(n_522), .Y(n_520) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_505), .A2(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g548 ( .A(n_506), .Y(n_548) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g622 ( .A(n_510), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g634 ( .A(n_510), .Y(n_634) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_510), .Y(n_812) );
OR2x2_ASAP7_75t_L g825 ( .A(n_510), .B(n_826), .Y(n_825) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_524), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_511), .B(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g598 ( .A(n_511), .Y(n_598) );
AND2x2_ASAP7_75t_L g645 ( .A(n_511), .B(n_646), .Y(n_645) );
NAND2x1p5_ASAP7_75t_SL g664 ( .A(n_511), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_511), .B(n_599), .Y(n_714) );
INVx1_ASAP7_75t_L g803 ( .A(n_511), .Y(n_803) );
AND2x2_ASAP7_75t_L g832 ( .A(n_511), .B(n_525), .Y(n_832) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_520), .B(n_523), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
BUFx4f_ASAP7_75t_L g587 ( .A(n_518), .Y(n_587) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g599 ( .A(n_525), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_525), .B(n_625), .Y(n_647) );
INVx1_ASAP7_75t_L g667 ( .A(n_525), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_525), .B(n_601), .Y(n_719) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_549), .Y(n_533) );
OR2x2_ASAP7_75t_L g616 ( .A(n_534), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g723 ( .A(n_534), .B(n_672), .Y(n_723) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g632 ( .A(n_535), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_535), .B(n_652), .Y(n_651) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_535), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g595 ( .A(n_536), .Y(n_595) );
BUFx3_ASAP7_75t_L g643 ( .A(n_536), .Y(n_643) );
AND2x2_ASAP7_75t_L g679 ( .A(n_536), .B(n_660), .Y(n_679) );
AND2x2_ASAP7_75t_L g759 ( .A(n_536), .B(n_605), .Y(n_759) );
AND2x2_ASAP7_75t_L g772 ( .A(n_536), .B(n_563), .Y(n_772) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
OAI21x1_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_544), .B(n_547), .Y(n_538) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g712 ( .A(n_549), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_549), .B(n_642), .Y(n_720) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_562), .Y(n_549) );
AND2x2_ASAP7_75t_L g631 ( .A(n_550), .B(n_563), .Y(n_631) );
INVx1_ASAP7_75t_L g739 ( .A(n_550), .Y(n_739) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g593 ( .A(n_551), .B(n_563), .Y(n_593) );
AND2x2_ASAP7_75t_L g656 ( .A(n_551), .B(n_562), .Y(n_656) );
AOI21x1_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_556), .B(n_559), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_561), .A2(n_582), .B(n_588), .Y(n_581) );
AND2x2_ASAP7_75t_L g614 ( .A(n_562), .B(n_605), .Y(n_614) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g604 ( .A(n_563), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g672 ( .A(n_563), .B(n_605), .Y(n_672) );
INVx1_ASAP7_75t_L g683 ( .A(n_563), .Y(n_683) );
AND2x2_ASAP7_75t_L g746 ( .A(n_563), .B(n_595), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_592), .B1(n_596), .B2(n_602), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_575), .A2(n_645), .B1(n_648), .B2(n_650), .Y(n_644) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
OR2x2_ASAP7_75t_L g724 ( .A(n_577), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g830 ( .A(n_577), .Y(n_830) );
INVx1_ASAP7_75t_L g689 ( .A(n_578), .Y(n_689) );
OR2x2_ASAP7_75t_L g752 ( .A(n_578), .B(n_647), .Y(n_752) );
OR2x2_ASAP7_75t_L g623 ( .A(n_579), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_579), .B(n_598), .Y(n_699) );
AND2x2_ASAP7_75t_L g716 ( .A(n_579), .B(n_643), .Y(n_716) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_579), .Y(n_733) );
INVxp67_ASAP7_75t_L g781 ( .A(n_579), .Y(n_781) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g601 ( .A(n_580), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_587), .Y(n_582) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_593), .Y(n_691) );
INVx3_ASAP7_75t_L g696 ( .A(n_593), .Y(n_696) );
AND2x2_ASAP7_75t_L g709 ( .A(n_593), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g809 ( .A(n_593), .B(n_771), .Y(n_809) );
INVx1_ASAP7_75t_L g603 ( .A(n_594), .Y(n_603) );
OR2x2_ASAP7_75t_L g786 ( .A(n_594), .B(n_761), .Y(n_786) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g710 ( .A(n_595), .B(n_620), .Y(n_710) );
AND2x2_ASAP7_75t_L g731 ( .A(n_595), .B(n_656), .Y(n_731) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_597), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g732 ( .A(n_597), .Y(n_732) );
AND2x2_ASAP7_75t_L g774 ( .A(n_597), .B(n_775), .Y(n_774) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g675 ( .A(n_598), .Y(n_675) );
AND2x2_ASAP7_75t_L g706 ( .A(n_598), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_598), .B(n_665), .Y(n_725) );
AND2x2_ASAP7_75t_L g674 ( .A(n_600), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g790 ( .A(n_600), .Y(n_790) );
AND2x2_ASAP7_75t_L g813 ( .A(n_600), .B(n_803), .Y(n_813) );
INVx1_ASAP7_75t_L g826 ( .A(n_600), .Y(n_826) );
INVx2_ASAP7_75t_L g665 ( .A(n_601), .Y(n_665) );
OR2x2_ASAP7_75t_L g761 ( .A(n_601), .B(n_625), .Y(n_761) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_604), .B(n_642), .Y(n_649) );
INVx2_ASAP7_75t_L g620 ( .A(n_605), .Y(n_620) );
INVx2_ASAP7_75t_L g660 ( .A(n_605), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_605), .B(n_618), .Y(n_682) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B(n_621), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_614), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g755 ( .A(n_617), .B(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx2_ASAP7_75t_L g661 ( .A(n_618), .Y(n_661) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g652 ( .A(n_620), .Y(n_652) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g635 ( .A(n_623), .Y(n_635) );
INVxp67_ASAP7_75t_L g806 ( .A(n_623), .Y(n_806) );
OR2x2_ASAP7_75t_L g708 ( .A(n_624), .B(n_665), .Y(n_708) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_627), .B(n_636), .C(n_644), .D(n_653), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_633), .C(n_635), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g822 ( .A1(n_629), .A2(n_823), .B(n_825), .C(n_827), .Y(n_822) );
OR2x6_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_631), .B(n_679), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_631), .B(n_735), .C(n_737), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_631), .B(n_710), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_631), .A2(n_736), .B1(n_828), .B2(n_831), .C(n_833), .Y(n_827) );
INVx1_ASAP7_75t_L g818 ( .A(n_632), .Y(n_818) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_640), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_637), .A2(n_645), .B1(n_680), .B2(n_754), .C(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_639), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g704 ( .A(n_640), .Y(n_704) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2x1p5_ASAP7_75t_L g658 ( .A(n_642), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g819 ( .A(n_642), .B(n_670), .Y(n_819) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx2_ASAP7_75t_L g655 ( .A(n_643), .Y(n_655) );
AND3x1_ASAP7_75t_L g828 ( .A(n_643), .B(n_829), .C(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g698 ( .A(n_647), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g768 ( .A(n_650), .Y(n_768) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g744 ( .A(n_652), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g771 ( .A(n_652), .Y(n_771) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_657), .B(n_662), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
NAND2x1_ASAP7_75t_L g669 ( .A(n_655), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g736 ( .A(n_656), .Y(n_736) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g692 ( .A(n_660), .Y(n_692) );
OR2x2_ASAP7_75t_L g671 ( .A(n_661), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g784 ( .A(n_661), .Y(n_784) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_663), .B(n_811), .Y(n_810) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
OR2x2_ASAP7_75t_L g740 ( .A(n_664), .B(n_688), .Y(n_740) );
INVx2_ASAP7_75t_L g829 ( .A(n_664), .Y(n_829) );
INVx1_ASAP7_75t_L g703 ( .A(n_665), .Y(n_703) );
NOR4xp25_ASAP7_75t_L g833 ( .A(n_665), .B(n_696), .C(n_834), .D(n_835), .Y(n_833) );
INVx1_ASAP7_75t_L g835 ( .A(n_666), .Y(n_835) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx3_ASAP7_75t_L g821 ( .A(n_667), .Y(n_821) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_673), .B(n_676), .C(n_684), .Y(n_668) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g808 ( .A(n_671), .Y(n_808) );
INVx2_ASAP7_75t_L g793 ( .A(n_672), .Y(n_793) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_674), .A2(n_677), .B(n_680), .Y(n_676) );
OR2x2_ASAP7_75t_L g760 ( .A(n_675), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g778 ( .A(n_675), .B(n_779), .Y(n_778) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g694 ( .A(n_679), .Y(n_694) );
AND2x4_ASAP7_75t_SL g783 ( .A(n_679), .B(n_784), .Y(n_783) );
INVx3_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_682), .Y(n_749) );
INVx1_ASAP7_75t_L g756 ( .A(n_683), .Y(n_756) );
AOI32xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_690), .A3(n_692), .B1(n_693), .B2(n_697), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_687), .B(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_687), .Y(n_748) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g765 ( .A(n_688), .B(n_703), .Y(n_765) );
INVx2_ASAP7_75t_L g779 ( .A(n_688), .Y(n_779) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_696), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_704), .B(n_705), .C(n_721), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_711), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g762 ( .A(n_710), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_710), .B(n_797), .Y(n_796) );
OAI32xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .A3(n_715), .B1(n_717), .B2(n_720), .Y(n_711) );
INVx1_ASAP7_75t_L g797 ( .A(n_712), .Y(n_797) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g789 ( .A(n_714), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_798), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g727 ( .A(n_728), .B(n_753), .C(n_766), .D(n_794), .Y(n_727) );
NOR2xp67_ASAP7_75t_L g728 ( .A(n_729), .B(n_741), .Y(n_728) );
OAI32xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .A3(n_733), .B1(n_734), .B2(n_740), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g780 ( .A(n_732), .B(n_781), .Y(n_780) );
OAI32xp33_ASAP7_75t_L g785 ( .A1(n_732), .A2(n_786), .A3(n_787), .B1(n_789), .B2(n_791), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_733), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g799 ( .A(n_735), .B(n_800), .Y(n_799) );
INVx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g792 ( .A(n_738), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g824 ( .A(n_738), .Y(n_824) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g788 ( .A(n_739), .Y(n_788) );
OAI22x1_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_747), .B1(n_749), .B2(n_750), .Y(n_741) );
INVx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_751), .B(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NOR2x1_ASAP7_75t_L g817 ( .A(n_755), .B(n_818), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B1(n_762), .B2(n_763), .Y(n_757) );
NAND2x1_ASAP7_75t_L g823 ( .A(n_759), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g834 ( .A(n_759), .Y(n_834) );
INVx2_ASAP7_75t_L g775 ( .A(n_761), .Y(n_775) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NOR3xp33_ASAP7_75t_SL g766 ( .A(n_767), .B(n_776), .C(n_785), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B(n_773), .Y(n_767) );
NAND2xp33_ASAP7_75t_L g795 ( .A(n_769), .B(n_796), .Y(n_795) );
INVx2_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x4_ASAP7_75t_L g831 ( .A(n_775), .B(n_832), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_780), .B(n_782), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x4_ASAP7_75t_L g802 ( .A(n_779), .B(n_803), .Y(n_802) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_781), .Y(n_801) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVxp67_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND3xp33_ASAP7_75t_SL g798 ( .A(n_799), .B(n_804), .C(n_816), .Y(n_798) );
AND2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g807 ( .A(n_803), .Y(n_807) );
AOI222xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_808), .B1(n_809), .B2(n_810), .C1(n_813), .C2(n_814), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
O2A1O1Ixp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_819), .B(n_820), .C(n_822), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_847), .B(n_849), .Y(n_838) );
OAI21xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_843), .B(n_846), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
INVx6_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx10_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
endmodule