module fake_jpeg_4188_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_20),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_28),
.B1(n_22),
.B2(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_51),
.Y(n_82)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_22),
.B(n_19),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_17),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_59),
.B1(n_70),
.B2(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_19),
.B1(n_20),
.B2(n_44),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_88),
.B1(n_71),
.B2(n_20),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_19),
.B1(n_21),
.B2(n_31),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_94),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_31),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_37),
.C(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_61),
.Y(n_114)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_102),
.Y(n_148)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_81),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_106),
.A2(n_108),
.B1(n_115),
.B2(n_18),
.Y(n_158)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_114),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_51),
.B1(n_75),
.B2(n_59),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_70),
.B1(n_74),
.B2(n_73),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_123),
.B1(n_128),
.B2(n_85),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_71),
.B1(n_62),
.B2(n_65),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_66),
.B1(n_53),
.B2(n_55),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_56),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_129),
.Y(n_133)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_95),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_84),
.A2(n_41),
.B1(n_50),
.B2(n_21),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_141),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_93),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_135),
.A2(n_23),
.B(n_32),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_140),
.C(n_145),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_97),
.B1(n_91),
.B2(n_92),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_144),
.B1(n_102),
.B2(n_101),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_92),
.B1(n_97),
.B2(n_91),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_153),
.B1(n_158),
.B2(n_114),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_85),
.C(n_83),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_83),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_99),
.C(n_50),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_23),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_157),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_120),
.B1(n_129),
.B2(n_110),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_25),
.B1(n_118),
.B2(n_116),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_41),
.B1(n_61),
.B2(n_33),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_33),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_25),
.A3(n_18),
.B1(n_34),
.B2(n_23),
.Y(n_157)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_161),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_150),
.A2(n_152),
.B1(n_147),
.B2(n_143),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_184),
.B(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_174),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_171),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_130),
.B1(n_155),
.B2(n_131),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

BUFx24_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_104),
.B1(n_24),
.B2(n_30),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_176),
.Y(n_201)
);

BUFx24_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_105),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_134),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_126),
.B1(n_122),
.B2(n_116),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_181),
.A2(n_152),
.B1(n_131),
.B2(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_112),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_197),
.B(n_181),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_206),
.B(n_184),
.Y(n_220)
);

NAND2xp67_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_136),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_214),
.B1(n_174),
.B2(n_182),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_133),
.B(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_133),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_157),
.B1(n_132),
.B2(n_154),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_160),
.B(n_112),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_203),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_218),
.A2(n_227),
.B(n_230),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_162),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_222),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_225),
.B(n_232),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_223),
.A2(n_226),
.B1(n_203),
.B2(n_191),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_165),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_209),
.B(n_193),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_183),
.B(n_178),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_192),
.A2(n_198),
.B1(n_201),
.B2(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_164),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_231),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_161),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_169),
.C(n_172),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_242),
.C(n_191),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_186),
.B(n_166),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_237),
.B1(n_200),
.B2(n_213),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_185),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_240),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_167),
.B1(n_173),
.B2(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_177),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_177),
.C(n_173),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_0),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_201),
.B1(n_190),
.B2(n_193),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_252),
.B1(n_224),
.B2(n_235),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_240),
.B1(n_216),
.B2(n_223),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_210),
.C(n_205),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_220),
.C(n_225),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_210),
.B1(n_208),
.B2(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_256),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_200),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_264),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_238),
.B1(n_32),
.B2(n_2),
.Y(n_271)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_0),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_189),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_189),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_3),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_253),
.B1(n_250),
.B2(n_246),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_272),
.B1(n_255),
.B2(n_251),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_270),
.C(n_273),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_234),
.C(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_79),
.C(n_32),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_277),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_0),
.C(n_2),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_16),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_282),
.B(n_283),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_3),
.C(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_283),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_261),
.B1(n_247),
.B2(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_289),
.B1(n_292),
.B2(n_295),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_266),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_253),
.C(n_257),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_6),
.C(n_8),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_269),
.A2(n_270),
.B1(n_259),
.B2(n_273),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_285),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_297),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_11),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_288),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_244),
.B1(n_7),
.B2(n_8),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.C(n_306),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_12),
.B1(n_7),
.B2(n_8),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_308),
.A2(n_312),
.B(n_313),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_13),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_13),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_286),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_294),
.Y(n_316)
);

OAI21x1_ASAP7_75t_SL g329 ( 
.A1(n_316),
.A2(n_319),
.B(n_320),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_13),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_321),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_306),
.B(n_309),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_9),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_9),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_6),
.C(n_10),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_14),
.B(n_15),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_10),
.B(n_12),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_327),
.A2(n_328),
.B(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_10),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_317),
.B(n_324),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_14),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_334),
.B(n_322),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_328),
.A2(n_323),
.B(n_316),
.Y(n_337)
);

AOI21xp33_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_338),
.B(n_333),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_320),
.B(n_15),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_335),
.C(n_336),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_343),
.Y(n_344)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_341),
.B(n_15),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_16),
.Y(n_346)
);


endmodule