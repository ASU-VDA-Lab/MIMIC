module real_jpeg_32461_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_578;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_634;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_0),
.Y(n_258)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_0),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_0),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_0),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_0),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_2),
.A2(n_64),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_2),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_2),
.A2(n_232),
.B1(n_324),
.B2(n_519),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_2),
.A2(n_324),
.B1(n_579),
.B2(n_584),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_3),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_4),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_4),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_4),
.A2(n_286),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_4),
.A2(n_286),
.B1(n_453),
.B2(n_455),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_4),
.A2(n_286),
.B1(n_544),
.B2(n_546),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_5),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_6),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_6),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22x1_ASAP7_75t_L g166 ( 
.A1(n_7),
.A2(n_52),
.B1(n_167),
.B2(n_171),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_7),
.A2(n_52),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_7),
.A2(n_52),
.B1(n_312),
.B2(n_316),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_8),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_8),
.Y(n_425)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_8),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_9),
.A2(n_62),
.B1(n_121),
.B2(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_9),
.A2(n_62),
.B1(n_145),
.B2(n_149),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_9),
.A2(n_62),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_10),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_10),
.A2(n_79),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_10),
.A2(n_79),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_10),
.A2(n_79),
.B1(n_421),
.B2(n_426),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_11),
.B(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_11),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_11),
.B(n_68),
.Y(n_506)
);

OAI32xp33_ASAP7_75t_L g526 ( 
.A1(n_11),
.A2(n_519),
.A3(n_527),
.B1(n_532),
.B2(n_536),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_11),
.A2(n_439),
.B1(n_465),
.B2(n_560),
.Y(n_559)
);

OAI21xp33_ASAP7_75t_L g644 ( 
.A1(n_11),
.A2(n_318),
.B(n_588),
.Y(n_644)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_12),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_13),
.A2(n_63),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_13),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_13),
.A2(n_145),
.B1(n_374),
.B2(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_13),
.A2(n_374),
.B1(n_565),
.B2(n_568),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g599 ( 
.A1(n_13),
.A2(n_374),
.B1(n_600),
.B2(n_603),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_20),
.B(n_679),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_14),
.B(n_680),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_15),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_15),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_15),
.A2(n_86),
.B1(n_207),
.B2(n_211),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_15),
.A2(n_86),
.B1(n_272),
.B2(n_274),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_15),
.A2(n_86),
.B1(n_356),
.B2(n_359),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_16),
.Y(n_108)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_16),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_16),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_17),
.A2(n_192),
.B1(n_193),
.B2(n_197),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_17),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_17),
.A2(n_192),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_17),
.A2(n_192),
.B1(n_365),
.B2(n_370),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_17),
.A2(n_192),
.B1(n_499),
.B2(n_503),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_18),
.Y(n_148)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_18),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_182),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_181),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_69),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_24),
.B(n_69),
.Y(n_181)
);

AOI22x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_51),
.B1(n_61),
.B2(n_67),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_25),
.A2(n_51),
.B1(n_67),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_26),
.A2(n_72),
.B1(n_80),
.B2(n_90),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_27),
.A2(n_67),
.B1(n_73),
.B2(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_28),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_28),
.B(n_323),
.Y(n_322)
);

AO22x1_ASAP7_75t_L g372 ( 
.A1(n_28),
.A2(n_68),
.B1(n_323),
.B2(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_28),
.B(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_42),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_37),
.Y(n_417)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_45),
.Y(n_153)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_46),
.Y(n_170)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_46),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_47),
.Y(n_410)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_50),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_50),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_50),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_50),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_60),
.Y(n_464)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_66),
.Y(n_200)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_68),
.B(n_191),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_68),
.B(n_282),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_68),
.B(n_373),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_177),
.C(n_179),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_70),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_91),
.C(n_128),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_71),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_80),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_85),
.Y(n_288)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_85),
.Y(n_379)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_87),
.Y(n_411)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_92),
.B(n_190),
.C(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_93),
.B(n_128),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_93),
.A2(n_204),
.B1(n_205),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_93),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_118),
.B(n_120),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_94),
.A2(n_118),
.B1(n_120),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_94),
.A2(n_118),
.B1(n_452),
.B2(n_459),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_94),
.B(n_452),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_94),
.B(n_634),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_95),
.A2(n_119),
.B1(n_231),
.B2(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_95),
.A2(n_119),
.B1(n_271),
.B2(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_95),
.A2(n_119),
.B1(n_301),
.B2(n_364),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_95),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_95),
.A2(n_119),
.B1(n_518),
.B2(n_564),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_103),
.B2(n_105),
.Y(n_96)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_97),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_98),
.Y(n_234)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_98),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_98),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_98),
.Y(n_638)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_103),
.Y(n_630)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_106),
.B(n_465),
.Y(n_631)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_107),
.Y(n_304)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22x1_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_109)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

BUFx2_ASAP7_75t_SL g602 ( 
.A(n_110),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_111),
.Y(n_361)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_111),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_118),
.B(n_452),
.Y(n_523)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_118),
.Y(n_574)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_123),
.Y(n_273)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AO22x2_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_144),
.B1(n_154),
.B2(n_166),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_129),
.A2(n_144),
.B(n_154),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_129),
.A2(n_154),
.B1(n_166),
.B2(n_206),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_129),
.A2(n_154),
.B1(n_206),
.B2(n_240),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_129),
.A2(n_468),
.B(n_469),
.Y(n_467)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22x1_ASAP7_75t_L g381 ( 
.A1(n_130),
.A2(n_382),
.B1(n_386),
.B2(n_387),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_130),
.A2(n_491),
.B(n_492),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_R g576 ( 
.A(n_130),
.B(n_465),
.Y(n_576)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_131),
.A2(n_154),
.B1(n_240),
.B2(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_131),
.B(n_383),
.Y(n_442)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_137),
.B1(n_140),
.B2(n_142),
.Y(n_132)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_133),
.Y(n_617)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_135),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_136),
.Y(n_278)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_143),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_156),
.B1(n_159),
.B2(n_163),
.Y(n_155)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_147),
.Y(n_384)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_147),
.Y(n_472)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_148),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_148),
.Y(n_562)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_152),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_154),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_154),
.B(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_154),
.B(n_383),
.Y(n_492)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_164),
.Y(n_336)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_164),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_165),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_169),
.B(n_533),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_179),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_339),
.B(n_670),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_219),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_184),
.A2(n_671),
.B(n_677),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_217),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_185),
.B(n_217),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_201),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_190),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_196),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_196),
.Y(n_327)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_210),
.Y(n_531)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_215),
.Y(n_408)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_290),
.Y(n_220)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_221),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g676 ( 
.A(n_222),
.B(n_224),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.C(n_248),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_225),
.B(n_228),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_239),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_229),
.B(n_239),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_234),
.Y(n_454)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_249),
.B(n_338),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_279),
.B(n_280),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_270),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_251),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_251),
.B(n_270),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_259),
.B(n_264),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_253),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_253),
.A2(n_355),
.B1(n_419),
.B2(n_427),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_253),
.B(n_543),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_253),
.A2(n_427),
.B1(n_598),
.B2(n_605),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_254),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_258),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_259),
.A2(n_542),
.B(n_599),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_259),
.B(n_465),
.Y(n_646)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_260),
.Y(n_362)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_310),
.B1(n_311),
.B2(n_318),
.Y(n_309)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_265),
.Y(n_545)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_266),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx4f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

XNOR2x1_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_280),
.Y(n_294)
);

NAND2x1_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_281),
.B(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_337),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_291),
.B(n_337),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.C(n_297),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_293),
.B(n_296),
.Y(n_389)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2x2_ASAP7_75t_L g388 ( 
.A(n_297),
.B(n_389),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_319),
.C(n_328),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

BUFx4f_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_309),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_309),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_318),
.B1(n_354),
.B2(n_362),
.Y(n_353)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_316),
.Y(n_546)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_317),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_317),
.Y(n_587)
);

OA22x2_ASAP7_75t_L g494 ( 
.A1(n_318),
.A2(n_420),
.B1(n_495),
.B2(n_498),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_318),
.A2(n_578),
.B(n_588),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_320),
.A2(n_329),
.B1(n_330),
.B2(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_322),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_321),
.B(n_461),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_324),
.A2(n_435),
.B(n_438),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_324),
.B(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_507),
.B(n_662),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_444),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_342),
.A2(n_663),
.B(n_665),
.Y(n_662)
);

OA21x2_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_388),
.B(n_390),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_343),
.B(n_388),
.Y(n_669)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_344),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.C(n_350),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_346),
.B(n_349),
.Y(n_392)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_371),
.C(n_380),
.Y(n_351)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_363),
.Y(n_352)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_353),
.Y(n_475)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_363),
.Y(n_476)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx4f_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_369),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_372),
.B(n_381),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_386),
.A2(n_434),
.B(n_442),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_386),
.A2(n_442),
.B(n_559),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_388),
.B(n_668),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_391),
.B(n_393),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_403),
.B(n_443),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_400),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_400),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_395),
.A2(n_396),
.B1(n_400),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_400),
.Y(n_479)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_403),
.B(n_478),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_429),
.C(n_432),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_449),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_418),
.Y(n_405)
);

XOR2x2_ASAP7_75t_L g487 ( 
.A(n_406),
.B(n_418),
.Y(n_487)
);

AOI32xp33_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_409),
.A3(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_424),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx6_ASAP7_75t_L g502 ( 
.A(n_425),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_429),
.A2(n_430),
.B1(n_432),
.B2(n_433),
.Y(n_449)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_434),
.Y(n_468)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx8_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_477),
.B(n_480),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_445),
.B(n_477),
.C(n_664),
.Y(n_663)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_450),
.C(n_473),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_483),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_474),
.Y(n_483)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_460),
.C(n_467),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_467),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_458),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_486),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_463),
.A2(n_465),
.B(n_466),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_537),
.Y(n_536)
);

OAI21xp33_ASAP7_75t_SL g634 ( 
.A1(n_465),
.A2(n_631),
.B(n_635),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_465),
.B(n_574),
.Y(n_641)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

INVx3_ASAP7_75t_SL g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_484),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_482),
.B(n_484),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_487),
.C(n_488),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_485),
.B(n_548),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_487),
.A2(n_488),
.B1(n_489),
.B2(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_487),
.Y(n_549)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.C(n_506),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_506),
.Y(n_514)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx4f_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_498),
.A2(n_539),
.B(n_542),
.Y(n_538)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OAI21x1_ASAP7_75t_SL g508 ( 
.A1(n_509),
.A2(n_550),
.B(n_660),
.Y(n_508)
);

AND2x4_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_547),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_511),
.B(n_661),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_515),
.C(n_524),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_513),
.B(n_554),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_515),
.A2(n_516),
.B1(n_525),
.B2(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

OAI21xp33_ASAP7_75t_SL g516 ( 
.A1(n_517),
.A2(n_518),
.B(n_523),
.Y(n_516)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_523),
.B(n_633),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_525),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_538),
.Y(n_525)
);

XOR2x2_ASAP7_75t_L g557 ( 
.A(n_526),
.B(n_538),
.Y(n_557)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_541),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_543),
.B(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_545),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_547),
.Y(n_661)
);

AOI21x1_ASAP7_75t_L g550 ( 
.A1(n_551),
.A2(n_594),
.B(n_659),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_569),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_553),
.B(n_556),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_553),
.B(n_556),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_558),
.C(n_563),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_571),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_563),
.Y(n_571)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_564),
.A2(n_574),
.B(n_575),
.Y(n_573)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx3_ASAP7_75t_SL g566 ( 
.A(n_567),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_570),
.B(n_572),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_570),
.B(n_572),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_576),
.C(n_577),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_573),
.B(n_576),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_577),
.B(n_655),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_578),
.Y(n_605)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

OAI211xp5_ASAP7_75t_SL g594 ( 
.A1(n_595),
.A2(n_653),
.B(n_657),
.C(n_658),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_596),
.A2(n_639),
.B(n_652),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_597),
.B(n_606),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_597),
.B(n_606),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_632),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_607),
.B(n_632),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_608),
.A2(n_614),
.B(n_623),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_615),
.B(n_618),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_624),
.A2(n_629),
.B(n_631),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_636),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_640),
.A2(n_643),
.B(n_651),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_641),
.B(n_642),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_641),
.B(n_642),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_644),
.B(n_645),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_646),
.B(n_647),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_648),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

NOR2x1_ASAP7_75t_L g653 ( 
.A(n_654),
.B(n_656),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_654),
.B(n_656),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_666),
.A2(n_667),
.B(n_669),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_672),
.A2(n_674),
.B(n_675),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_673),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_676),
.Y(n_675)
);

CKINVDCx16_ASAP7_75t_R g677 ( 
.A(n_678),
.Y(n_677)
);


endmodule