module fake_netlist_6_4064_n_1897 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1897);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1897;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_0),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_73),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

BUFx8_ASAP7_75t_SL g198 ( 
.A(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_88),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_118),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_116),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_138),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_62),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_42),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_131),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_92),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_84),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_164),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_50),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_48),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_25),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_7),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_10),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_18),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_18),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_117),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_38),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_113),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_20),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_139),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_119),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_151),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_3),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_145),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_15),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_42),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_56),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_53),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_15),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_94),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_149),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_85),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_181),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_27),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_135),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_159),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_167),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_29),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_51),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_57),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_101),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_33),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_171),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_67),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_57),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_62),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_0),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_124),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_71),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_157),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_179),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_87),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_33),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_58),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_95),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_79),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_150),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_99),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_19),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_37),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_165),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_185),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_115),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_170),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_161),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_19),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_40),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_53),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_107),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_86),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_29),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_153),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_28),
.Y(n_289)
);

BUFx2_ASAP7_75t_R g290 ( 
.A(n_100),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_121),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_187),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_154),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_1),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_8),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_7),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_175),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_24),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_65),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_105),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_60),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_44),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_41),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_24),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_32),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_69),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_166),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_186),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_74),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_59),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_40),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_52),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_9),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_190),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_162),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_97),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_136),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_160),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_180),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_17),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_89),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_36),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_93),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_127),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_44),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_177),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_146),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_14),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_22),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_39),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_132),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_148),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_55),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_76),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_48),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_98),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_111),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_46),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_46),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_188),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_3),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_147),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_23),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_77),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_60),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_6),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_4),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_112),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_109),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_43),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_39),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_126),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_27),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_81),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_61),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_63),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_22),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_26),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_45),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_9),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_59),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_47),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_1),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_134),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_52),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_25),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_43),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_172),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_72),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_183),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_96),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_80),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_30),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_28),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_251),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_210),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_268),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_251),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_198),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_263),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_193),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_191),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_251),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_208),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_307),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_226),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_251),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_196),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_200),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_215),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_201),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_251),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_202),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_223),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_258),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_287),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_258),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_203),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_191),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_209),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_211),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_287),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_287),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_287),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_287),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_214),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_218),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_227),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_229),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_274),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_204),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_328),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_226),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_351),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_225),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_237),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_208),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_237),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_216),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_204),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_235),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_205),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_329),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_331),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_331),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_243),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_244),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_352),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_350),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_207),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_207),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_246),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_249),
.Y(n_451)
);

BUFx2_ASAP7_75t_SL g452 ( 
.A(n_231),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_257),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_261),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_221),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_205),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_221),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_316),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_228),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_274),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_269),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_264),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_228),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_373),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_316),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_266),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_271),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_272),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_377),
.B(n_231),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_377),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_380),
.B(n_286),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_398),
.B(n_288),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_380),
.B(n_286),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_382),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_387),
.B(n_225),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_386),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_382),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_386),
.B(n_245),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_384),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_269),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_391),
.B(n_245),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_392),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_416),
.A2(n_375),
.B1(n_224),
.B2(n_303),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_416),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_403),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_393),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_414),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_396),
.B(n_276),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_400),
.B(n_192),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_407),
.B(n_279),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_407),
.B(n_281),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_425),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_398),
.B(n_288),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_457),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_408),
.B(n_291),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_409),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_395),
.Y(n_519)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_387),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_457),
.A2(n_410),
.B(n_409),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_410),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_420),
.B(n_292),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_457),
.A2(n_197),
.B(n_192),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_430),
.B(n_426),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_421),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_430),
.B(n_252),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_422),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_423),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_423),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_430),
.B(n_252),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_424),
.B(n_293),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_429),
.B(n_297),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_429),
.B(n_284),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_433),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_435),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_435),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_436),
.B(n_452),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_436),
.B(n_197),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_527),
.B(n_397),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_521),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_482),
.B(n_389),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_402),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_488),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_521),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_521),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_527),
.B(n_405),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_394),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_488),
.B(n_432),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_493),
.B(n_406),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_526),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_496),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_547),
.B(n_411),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_526),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_483),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_478),
.A2(n_419),
.B1(n_431),
.B2(n_427),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_412),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_483),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_526),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_526),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_483),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_541),
.B(n_466),
.C(n_459),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_493),
.B(n_413),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_518),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_518),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_545),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_478),
.A2(n_379),
.B1(n_437),
.B2(n_415),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_505),
.B(n_443),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_481),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_518),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_518),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_528),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_500),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_529),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_528),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_514),
.A2(n_321),
.B1(n_363),
.B2(n_239),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_528),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_496),
.B(n_499),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_541),
.B(n_404),
.C(n_385),
.Y(n_597)
);

INVxp33_ASAP7_75t_L g598 ( 
.A(n_499),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_537),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_500),
.B(n_444),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_528),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_474),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_477),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_519),
.B(n_450),
.Y(n_604)
);

AO21x2_ASAP7_75t_L g605 ( 
.A1(n_524),
.A2(n_511),
.B(n_505),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_476),
.B(n_194),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_474),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_519),
.B(n_451),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_495),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_475),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_495),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_514),
.B(n_482),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_511),
.B(n_453),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_544),
.B(n_454),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_L g616 ( 
.A1(n_489),
.A2(n_195),
.B1(n_417),
.B2(n_230),
.Y(n_616)
);

OAI22x1_ASAP7_75t_L g617 ( 
.A1(n_494),
.A2(n_232),
.B1(n_241),
.B2(n_240),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_545),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_501),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_512),
.B(n_463),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_501),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_512),
.B(n_467),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_516),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_482),
.B(n_194),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_476),
.A2(n_452),
.B1(n_302),
.B2(n_313),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_510),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_510),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_516),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_522),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_477),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_544),
.B(n_468),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_517),
.B(n_469),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_541),
.B(n_434),
.C(n_206),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_522),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_525),
.Y(n_636)
);

AND3x2_ASAP7_75t_L g637 ( 
.A(n_537),
.B(n_314),
.C(n_250),
.Y(n_637)
);

BUFx6f_ASAP7_75t_SL g638 ( 
.A(n_476),
.Y(n_638)
);

HB1xp67_ASAP7_75t_SL g639 ( 
.A(n_470),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_525),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_476),
.B(n_199),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_530),
.B(n_439),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_532),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_492),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_530),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_489),
.A2(n_323),
.B1(n_315),
.B2(n_236),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_532),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_533),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_530),
.B(n_439),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_533),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_489),
.B(n_381),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_542),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_477),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_475),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_477),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_534),
.B(n_440),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_543),
.Y(n_660)
);

BUFx4f_ASAP7_75t_L g661 ( 
.A(n_477),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_517),
.B(n_256),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_534),
.B(n_288),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

AOI21x1_ASAP7_75t_L g665 ( 
.A1(n_472),
.A2(n_206),
.B(n_199),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_477),
.B(n_213),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_523),
.B(n_285),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_476),
.B(n_480),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_476),
.B(n_440),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_531),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_520),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_494),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_475),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_508),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_472),
.A2(n_524),
.B(n_508),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_523),
.B(n_299),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_508),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_520),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_531),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_481),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_486),
.B(n_217),
.C(n_213),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_480),
.B(n_441),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_535),
.B(n_540),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_492),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_531),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_531),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_480),
.B(n_217),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_508),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_535),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_481),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_481),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_540),
.B(n_320),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_480),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_520),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_480),
.B(n_441),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_480),
.B(n_300),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_546),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_689),
.B(n_349),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_596),
.B(n_438),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_596),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_683),
.B(n_520),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_669),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_612),
.B(n_284),
.Y(n_703)
);

BUFx5_ASAP7_75t_L g704 ( 
.A(n_550),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_620),
.B(n_520),
.Y(n_705)
);

AND2x2_ASAP7_75t_SL g706 ( 
.A(n_606),
.B(n_212),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_643),
.B(n_448),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_689),
.B(n_520),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_570),
.B(n_378),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_598),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_599),
.B(n_383),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_662),
.B(n_486),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_574),
.B(n_220),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_667),
.B(n_692),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_646),
.B(n_238),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_567),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_SL g717 ( 
.A(n_555),
.B(n_290),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_567),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_569),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_585),
.B(n_486),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_562),
.B(n_388),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_551),
.B(n_418),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_643),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_571),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_613),
.B(n_486),
.Y(n_725)
);

BUFx6f_ASAP7_75t_SL g726 ( 
.A(n_612),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_571),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_669),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_639),
.Y(n_730)
);

AO22x2_ASAP7_75t_L g731 ( 
.A1(n_681),
.A2(n_219),
.B1(n_222),
.B2(n_233),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_622),
.B(n_486),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_579),
.B(n_253),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_633),
.B(n_447),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_556),
.B(n_486),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_573),
.B(n_465),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_556),
.B(n_491),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_684),
.B(n_456),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_573),
.B(n_306),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_682),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_693),
.B(n_308),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_682),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_L g743 ( 
.A(n_693),
.B(n_317),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_556),
.B(n_491),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_668),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_568),
.B(n_491),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_579),
.B(n_259),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_568),
.B(n_491),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_674),
.A2(n_524),
.B(n_491),
.C(n_322),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_584),
.B(n_318),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_568),
.B(n_491),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_610),
.B(n_508),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_650),
.B(n_448),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_550),
.A2(n_449),
.B(n_455),
.C(n_464),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_554),
.A2(n_338),
.B1(n_319),
.B2(n_325),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_626),
.B(n_327),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_695),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_650),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_684),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_610),
.B(n_508),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_658),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_668),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_580),
.B(n_565),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_616),
.B(n_332),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_658),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_610),
.B(n_548),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_656),
.B(n_548),
.Y(n_767)
);

OR2x6_ASAP7_75t_L g768 ( 
.A(n_612),
.B(n_302),
.Y(n_768)
);

AO221x1_ASAP7_75t_L g769 ( 
.A1(n_617),
.A2(n_372),
.B1(n_247),
.B2(n_242),
.C(n_368),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_555),
.B(n_260),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_576),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_576),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_597),
.B(n_295),
.C(n_294),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_594),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_577),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_552),
.B(n_553),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_614),
.B(n_296),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_661),
.A2(n_548),
.B(n_473),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_563),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_572),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_656),
.B(n_673),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_673),
.B(n_548),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_673),
.B(n_548),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_552),
.B(n_546),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_668),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_668),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_553),
.B(n_546),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_SL g788 ( 
.A(n_557),
.B(n_372),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_557),
.A2(n_275),
.B1(n_301),
.B2(n_289),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_549),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_559),
.B(n_546),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_575),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_647),
.B(n_335),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_577),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_632),
.B(n_337),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_575),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_674),
.A2(n_212),
.B(n_250),
.C(n_365),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_582),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_559),
.B(n_560),
.Y(n_799)
);

INVx5_ASAP7_75t_L g800 ( 
.A(n_666),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_612),
.A2(n_341),
.B1(n_343),
.B2(n_371),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_561),
.B(n_298),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_583),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_560),
.B(n_546),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_641),
.B(n_304),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_634),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_591),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_634),
.B(n_310),
.C(n_305),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_578),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_SL g810 ( 
.A(n_681),
.B(n_372),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_625),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_581),
.B(n_222),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_645),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_591),
.B(n_345),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_676),
.B(n_353),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_589),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_589),
.Y(n_817)
);

INVx8_ASAP7_75t_L g818 ( 
.A(n_612),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_625),
.A2(n_449),
.B(n_455),
.C(n_458),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_566),
.B(n_355),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_587),
.B(n_234),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_600),
.B(n_357),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_587),
.B(n_234),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_615),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_588),
.B(n_248),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_588),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_590),
.B(n_593),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_590),
.B(n_248),
.Y(n_828)
);

BUFx6f_ASAP7_75t_SL g829 ( 
.A(n_606),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_677),
.A2(n_365),
.B1(n_322),
.B2(n_273),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_593),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_582),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_604),
.B(n_456),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_595),
.B(n_601),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_608),
.B(n_370),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_652),
.B(n_311),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_606),
.B(n_458),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_606),
.B(n_460),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_617),
.A2(n_275),
.B1(n_280),
.B2(n_267),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_595),
.B(n_254),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_677),
.A2(n_688),
.B1(n_625),
.B2(n_601),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_688),
.B(n_254),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_642),
.B(n_687),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_602),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_602),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_642),
.B(n_262),
.Y(n_846)
);

BUFx8_ASAP7_75t_L g847 ( 
.A(n_638),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_SL g848 ( 
.A(n_672),
.B(n_260),
.Y(n_848)
);

OAI21xp33_ASAP7_75t_L g849 ( 
.A1(n_663),
.A2(n_358),
.B(n_313),
.Y(n_849)
);

INVxp33_ASAP7_75t_L g850 ( 
.A(n_594),
.Y(n_850)
);

AO221x1_ASAP7_75t_L g851 ( 
.A1(n_582),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.C(n_344),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_615),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_607),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_642),
.B(n_265),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_607),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_687),
.B(n_265),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_L g857 ( 
.A(n_672),
.B(n_270),
.C(n_273),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_618),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_789),
.A2(n_687),
.B1(n_242),
.B2(n_241),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_781),
.A2(n_661),
.B(n_631),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_776),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_723),
.B(n_687),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_758),
.B(n_609),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_714),
.B(n_609),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_711),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_761),
.B(n_611),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_784),
.A2(n_675),
.B(n_586),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_779),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_800),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_799),
.B(n_611),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_789),
.A2(n_232),
.B1(n_240),
.B2(n_247),
.Y(n_871)
);

INVxp67_ASAP7_75t_SL g872 ( 
.A(n_704),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_774),
.B(n_619),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_704),
.B(n_621),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_780),
.Y(n_875)
);

NOR2xp67_ASAP7_75t_L g876 ( 
.A(n_730),
.B(n_665),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_704),
.B(n_785),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_704),
.B(n_776),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_738),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_850),
.B(n_621),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_765),
.B(n_627),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_857),
.A2(n_731),
.B1(n_769),
.B2(n_727),
.Y(n_882)
);

BUFx4f_ASAP7_75t_L g883 ( 
.A(n_703),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_792),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_719),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_857),
.A2(n_255),
.B1(n_267),
.B2(n_344),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_701),
.A2(n_661),
.B(n_631),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_796),
.Y(n_888)
);

AND2x6_ASAP7_75t_L g889 ( 
.A(n_785),
.B(n_664),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_745),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_731),
.A2(n_727),
.B1(n_839),
.B2(n_776),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_818),
.B(n_666),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_704),
.B(n_627),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_700),
.B(n_628),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_809),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_700),
.B(n_628),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_SL g897 ( 
.A1(n_807),
.A2(n_462),
.B1(n_364),
.B2(n_362),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_699),
.B(n_696),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_800),
.B(n_582),
.Y(n_899)
);

AND2x2_ASAP7_75t_SL g900 ( 
.A(n_706),
.B(n_839),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_800),
.B(n_582),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_800),
.B(n_664),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_720),
.A2(n_638),
.B1(n_666),
.B2(n_660),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_702),
.B(n_660),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_725),
.B(n_670),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_732),
.B(n_670),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_710),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_826),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_831),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_759),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_729),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_716),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_740),
.B(n_637),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_742),
.B(n_666),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_718),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_R g916 ( 
.A(n_717),
.B(n_665),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_734),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_715),
.B(n_260),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_731),
.A2(n_255),
.B1(n_330),
.B2(n_366),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_724),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_776),
.B(n_630),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_715),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_745),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_728),
.Y(n_924)
);

BUFx6f_ASAP7_75t_SL g925 ( 
.A(n_790),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_762),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_713),
.B(n_635),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_706),
.B(n_679),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_847),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_757),
.B(n_707),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_L g931 ( 
.A(n_818),
.B(n_635),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_735),
.A2(n_654),
.B(n_603),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_762),
.B(n_558),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_771),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_707),
.B(n_753),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_772),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_775),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_844),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_794),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_713),
.B(n_636),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_803),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_845),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_832),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_SL g944 ( 
.A(n_722),
.B(n_326),
.C(n_312),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_730),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_709),
.A2(n_638),
.B1(n_605),
.B2(n_636),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_853),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_818),
.B(n_666),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_712),
.A2(n_605),
.B1(n_640),
.B2(n_655),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_855),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_806),
.B(n_640),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_837),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_733),
.A2(n_270),
.B(n_277),
.C(n_278),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_813),
.B(n_644),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_837),
.B(n_648),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_786),
.B(n_685),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_843),
.A2(n_726),
.B1(n_708),
.B2(n_733),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_753),
.B(n_558),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_838),
.B(n_747),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_838),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_763),
.B(n_649),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_787),
.B(n_685),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_747),
.B(n_705),
.Y(n_963)
);

AND2x2_ASAP7_75t_SL g964 ( 
.A(n_811),
.B(n_277),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_811),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_847),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_851),
.A2(n_280),
.B1(n_289),
.B2(n_301),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_736),
.B(n_336),
.C(n_334),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_703),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_737),
.B(n_649),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_744),
.B(n_686),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_816),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_698),
.B(n_651),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_827),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_703),
.B(n_558),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_746),
.B(n_651),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_748),
.B(n_653),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_721),
.B(n_653),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_726),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_768),
.B(n_657),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_805),
.B(n_260),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_777),
.B(n_848),
.C(n_802),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_777),
.B(n_655),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_751),
.B(n_791),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_817),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_SL g986 ( 
.A(n_773),
.B(n_342),
.C(n_339),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_754),
.A2(n_659),
.B(n_623),
.C(n_624),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_841),
.B(n_686),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_739),
.B(n_659),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_830),
.A2(n_367),
.B1(n_282),
.B2(n_283),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_834),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_SL g992 ( 
.A1(n_770),
.A2(n_330),
.B1(n_282),
.B2(n_283),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_824),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_832),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_768),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_852),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_768),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_858),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_842),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_832),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_798),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_752),
.A2(n_654),
.B1(n_603),
.B2(n_678),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_812),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_802),
.B(n_623),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_804),
.B(n_760),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_766),
.B(n_624),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_764),
.B(n_629),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_833),
.B(n_605),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_767),
.B(n_697),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_782),
.B(n_697),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_829),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_821),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_783),
.B(n_678),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_801),
.B(n_657),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_829),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_808),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_823),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_836),
.B(n_340),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_795),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_825),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_828),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_819),
.B(n_278),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_840),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_854),
.B(n_671),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_836),
.B(n_460),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_846),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_754),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_856),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_814),
.B(n_464),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_869),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_872),
.A2(n_963),
.B(n_1005),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_864),
.B(n_849),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_1018),
.A2(n_819),
.B(n_750),
.C(n_793),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_869),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_864),
.B(n_741),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_1018),
.A2(n_743),
.B1(n_815),
.B2(n_756),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_917),
.B(n_675),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_982),
.A2(n_835),
.B1(n_822),
.B2(n_820),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_922),
.A2(n_749),
.B(n_755),
.C(n_778),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_938),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_900),
.A2(n_797),
.B1(n_309),
.B2(n_369),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1025),
.B(n_788),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_922),
.A2(n_900),
.B1(n_959),
.B2(n_957),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_905),
.A2(n_810),
.B(n_618),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_891),
.A2(n_694),
.B1(n_671),
.B2(n_369),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_984),
.A2(n_694),
.B(n_671),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_869),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_SL g1048 ( 
.A(n_883),
.B(n_309),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_970),
.A2(n_977),
.B(n_976),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_974),
.B(n_991),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_873),
.A2(n_324),
.B(n_564),
.C(n_586),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_879),
.B(n_346),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_935),
.A2(n_586),
.B1(n_564),
.B2(n_324),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_868),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_873),
.A2(n_586),
.B(n_564),
.C(n_347),
.Y(n_1055)
);

AND2x2_ASAP7_75t_SL g1056 ( 
.A(n_883),
.B(n_442),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_869),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_910),
.Y(n_1058)
);

INVx6_ASAP7_75t_L g1059 ( 
.A(n_1015),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_942),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_947),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_907),
.B(n_442),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_950),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_859),
.A2(n_348),
.B1(n_354),
.B2(n_356),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_875),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_888),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_953),
.A2(n_446),
.B(n_445),
.C(n_509),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_909),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_859),
.A2(n_871),
.B1(n_891),
.B2(n_919),
.Y(n_1069)
);

OAI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_918),
.A2(n_981),
.B(n_886),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_885),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_871),
.A2(n_359),
.B1(n_361),
.B2(n_374),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_880),
.B(n_592),
.Y(n_1073)
);

AND2x4_ASAP7_75t_SL g1074 ( 
.A(n_1015),
.B(n_445),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_930),
.B(n_446),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_979),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_SL g1077 ( 
.A1(n_964),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_884),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_874),
.A2(n_691),
.B(n_690),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_930),
.B(n_862),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_893),
.A2(n_691),
.B(n_690),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_SL g1082 ( 
.A1(n_992),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_929),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_865),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_SL g1085 ( 
.A(n_897),
.B(n_11),
.C(n_12),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_885),
.B(n_945),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_949),
.A2(n_867),
.B(n_905),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_895),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1006),
.A2(n_691),
.B(n_690),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_894),
.B(n_11),
.C(n_13),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1004),
.A2(n_504),
.B(n_502),
.C(n_507),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_954),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_861),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_965),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_SL g1095 ( 
.A1(n_995),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_1095)
);

CKINVDCx16_ASAP7_75t_R g1096 ( 
.A(n_966),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_887),
.A2(n_870),
.B(n_878),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_892),
.B(n_529),
.Y(n_1098)
);

INVxp33_ASAP7_75t_L g1099 ( 
.A(n_1011),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_SL g1100 ( 
.A(n_861),
.B(n_680),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_898),
.B(n_16),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_952),
.B(n_64),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_890),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_983),
.B(n_1004),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_965),
.B(n_21),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_906),
.A2(n_471),
.B(n_473),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_892),
.B(n_529),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_960),
.B(n_66),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_862),
.B(n_680),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_894),
.B(n_896),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1016),
.A2(n_1019),
.B1(n_1029),
.B2(n_973),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_995),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_997),
.Y(n_1113)
);

AND2x2_ASAP7_75t_SL g1114 ( 
.A(n_964),
.B(n_21),
.Y(n_1114)
);

NOR2xp67_ASAP7_75t_L g1115 ( 
.A(n_978),
.B(n_1011),
.Y(n_1115)
);

BUFx2_ASAP7_75t_SL g1116 ( 
.A(n_925),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_946),
.A2(n_471),
.B(n_479),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_861),
.B(n_680),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_SL g1119 ( 
.A(n_968),
.B(n_479),
.C(n_484),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_951),
.B(n_23),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_SL g1121 ( 
.A1(n_988),
.A2(n_502),
.B(n_504),
.C(n_507),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_863),
.B(n_866),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_R g1123 ( 
.A(n_925),
.B(n_125),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_919),
.A2(n_479),
.B1(n_484),
.B2(n_487),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_R g1125 ( 
.A(n_931),
.B(n_130),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_863),
.B(n_26),
.Y(n_1126)
);

AOI22x1_ASAP7_75t_L g1127 ( 
.A1(n_999),
.A2(n_490),
.B1(n_479),
.B2(n_484),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_943),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_908),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_961),
.A2(n_504),
.B(n_507),
.C(n_502),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_866),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_904),
.A2(n_881),
.B1(n_1028),
.B2(n_958),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1010),
.A2(n_515),
.B(n_485),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_986),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_896),
.A2(n_484),
.B(n_487),
.C(n_490),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_SL g1136 ( 
.A(n_926),
.B(n_120),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_912),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_943),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_915),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_997),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_882),
.A2(n_509),
.B1(n_498),
.B2(n_497),
.Y(n_1141)
);

BUFx8_ASAP7_75t_L g1142 ( 
.A(n_913),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_920),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_927),
.A2(n_940),
.B1(n_1023),
.B2(n_1021),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_969),
.B(n_110),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_881),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1003),
.A2(n_1012),
.B1(n_1020),
.B2(n_1017),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_911),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_904),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1013),
.A2(n_487),
.B(n_490),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_932),
.A2(n_487),
.B(n_490),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_860),
.A2(n_485),
.B(n_503),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_975),
.B(n_108),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_961),
.B(n_30),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_973),
.B(n_507),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_989),
.A2(n_502),
.B1(n_504),
.B2(n_485),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_955),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_994),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_892),
.B(n_948),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_986),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_SL g1161 ( 
.A1(n_928),
.A2(n_877),
.B(n_1014),
.C(n_1027),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_924),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_L g1163 ( 
.A(n_913),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_890),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_1007),
.A2(n_497),
.B(n_509),
.C(n_498),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_989),
.A2(n_509),
.B(n_497),
.C(n_498),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_958),
.B(n_497),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_968),
.A2(n_498),
.B(n_32),
.C(n_34),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1058),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1031),
.A2(n_1014),
.B(n_877),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1040),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1041),
.A2(n_903),
.A3(n_1007),
.B(n_1002),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1050),
.B(n_1026),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1070),
.B(n_944),
.C(n_886),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1150),
.A2(n_988),
.B(n_987),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1152),
.A2(n_971),
.B(n_1013),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1049),
.A2(n_1008),
.B(n_971),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1151),
.A2(n_1009),
.B(n_921),
.Y(n_1178)
);

OAI22x1_ASAP7_75t_L g1179 ( 
.A1(n_1043),
.A2(n_944),
.B1(n_980),
.B2(n_975),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1039),
.A2(n_1009),
.B(n_928),
.Y(n_1180)
);

AO22x2_ASAP7_75t_L g1181 ( 
.A1(n_1069),
.A2(n_882),
.B1(n_914),
.B2(n_980),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1060),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1087),
.A2(n_1024),
.B(n_876),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_1158),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1041),
.A2(n_1055),
.A3(n_1097),
.B(n_1033),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1110),
.B(n_914),
.Y(n_1186)
);

AOI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1044),
.A2(n_901),
.B(n_899),
.Y(n_1187)
);

OA22x2_ASAP7_75t_L g1188 ( 
.A1(n_1082),
.A2(n_1022),
.B1(n_948),
.B2(n_902),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1061),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1087),
.A2(n_962),
.B(n_956),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1161),
.A2(n_916),
.B(n_901),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1077),
.A2(n_990),
.B(n_967),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1093),
.Y(n_1193)
);

AND2x6_ASAP7_75t_L g1194 ( 
.A(n_1153),
.B(n_923),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1154),
.A2(n_1026),
.B(n_996),
.C(n_998),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1059),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1092),
.B(n_1026),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_L g1198 ( 
.A(n_1069),
.B(n_1104),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1035),
.A2(n_994),
.B(n_899),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1051),
.A2(n_1001),
.A3(n_1000),
.B(n_937),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1144),
.B(n_1026),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1042),
.A2(n_902),
.B(n_933),
.Y(n_1202)
);

OR2x6_ASAP7_75t_L g1203 ( 
.A(n_1159),
.B(n_948),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1122),
.B(n_990),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1063),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1159),
.B(n_926),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1036),
.A2(n_934),
.B(n_941),
.C(n_993),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1101),
.A2(n_936),
.B(n_985),
.C(n_972),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1038),
.A2(n_1111),
.B(n_1032),
.C(n_1147),
.Y(n_1209)
);

BUFx4f_ASAP7_75t_SL g1210 ( 
.A(n_1083),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_1142),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1157),
.B(n_916),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_L g1213 ( 
.A(n_1057),
.B(n_1000),
.Y(n_1213)
);

INVxp67_ASAP7_75t_L g1214 ( 
.A(n_1086),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_R g1215 ( 
.A(n_1037),
.B(n_1022),
.Y(n_1215)
);

OR2x6_ASAP7_75t_L g1216 ( 
.A(n_1159),
.B(n_943),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1073),
.A2(n_943),
.B(n_939),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1059),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1112),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1133),
.A2(n_967),
.B(n_962),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1114),
.A2(n_962),
.B1(n_889),
.B2(n_539),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1092),
.B(n_962),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1071),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1165),
.A2(n_889),
.B(n_539),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1168),
.A2(n_889),
.B(n_539),
.C(n_538),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1047),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1046),
.A2(n_889),
.B(n_515),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1078),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1088),
.Y(n_1229)
);

NOR4xp25_ASAP7_75t_L g1230 ( 
.A(n_1064),
.B(n_31),
.C(n_34),
.D(n_35),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1121),
.A2(n_889),
.B(n_515),
.Y(n_1231)
);

OA21x2_ASAP7_75t_L g1232 ( 
.A1(n_1155),
.A2(n_1166),
.B(n_1106),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1149),
.B(n_31),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1129),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1148),
.B(n_538),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1091),
.A2(n_515),
.B(n_503),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1130),
.A2(n_515),
.B(n_503),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1056),
.B(n_539),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1079),
.A2(n_515),
.B(n_503),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1090),
.B(n_539),
.C(n_538),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1141),
.A2(n_35),
.A3(n_36),
.B(n_38),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1149),
.B(n_45),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1120),
.A2(n_539),
.B(n_538),
.C(n_536),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1081),
.A2(n_1127),
.B(n_1089),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1141),
.A2(n_47),
.A3(n_49),
.B(n_50),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1132),
.B(n_1131),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1045),
.A2(n_49),
.A3(n_54),
.B(n_55),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1146),
.B(n_54),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1115),
.A2(n_539),
.B(n_538),
.C(n_536),
.Y(n_1249)
);

AO32x2_ASAP7_75t_L g1250 ( 
.A1(n_1064),
.A2(n_1072),
.A3(n_1124),
.B1(n_1156),
.B2(n_1138),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1054),
.B(n_61),
.Y(n_1251)
);

AO32x2_ASAP7_75t_L g1252 ( 
.A1(n_1072),
.A2(n_68),
.A3(n_70),
.B1(n_75),
.B2(n_78),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_1136),
.A2(n_82),
.B(n_83),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1135),
.A2(n_513),
.B(n_506),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1047),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1047),
.Y(n_1256)
);

AO22x2_ASAP7_75t_L g1257 ( 
.A1(n_1119),
.A2(n_90),
.B1(n_91),
.B2(n_102),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1094),
.B(n_103),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1084),
.B(n_539),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1065),
.B(n_538),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1066),
.B(n_538),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1062),
.Y(n_1262)
);

AOI22x1_ASAP7_75t_SL g1263 ( 
.A1(n_1134),
.A2(n_104),
.B1(n_123),
.B2(n_141),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1068),
.B(n_538),
.Y(n_1264)
);

NOR2xp67_ASAP7_75t_L g1265 ( 
.A(n_1052),
.B(n_142),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1093),
.A2(n_513),
.B(n_506),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1126),
.B(n_536),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1117),
.A2(n_513),
.B(n_506),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1142),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1137),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1105),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1163),
.B(n_536),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1153),
.B(n_536),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1139),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1163),
.B(n_536),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1124),
.A2(n_1053),
.B(n_1067),
.Y(n_1276)
);

NOR2x1_ASAP7_75t_L g1277 ( 
.A(n_1057),
.B(n_513),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1103),
.A2(n_1164),
.B(n_1118),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1143),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1164),
.A2(n_529),
.B(n_155),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1162),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1080),
.A2(n_1167),
.B(n_1100),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1098),
.A2(n_529),
.B(n_158),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1109),
.A2(n_529),
.B(n_174),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1113),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1085),
.B(n_143),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1160),
.A2(n_176),
.B1(n_178),
.B2(n_1140),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1075),
.Y(n_1288)
);

AOI31xp33_ASAP7_75t_L g1289 ( 
.A1(n_1095),
.A2(n_1099),
.A3(n_1108),
.B(n_1102),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1108),
.A2(n_1098),
.B(n_1107),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1074),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1048),
.B(n_1145),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1048),
.B(n_1138),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1096),
.B(n_1116),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1128),
.B(n_1098),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1107),
.A2(n_1128),
.B(n_1125),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1107),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1123),
.A2(n_963),
.B(n_1031),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1050),
.B(n_922),
.Y(n_1299)
);

NOR2xp67_ASAP7_75t_L g1300 ( 
.A(n_1111),
.B(n_813),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_SL g1301 ( 
.A1(n_1147),
.A2(n_1168),
.B(n_1144),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1110),
.B(n_1104),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1110),
.A2(n_900),
.B1(n_1069),
.B2(n_1050),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1031),
.A2(n_963),
.B(n_1049),
.Y(n_1304)
);

NOR2x1_ASAP7_75t_SL g1305 ( 
.A(n_1098),
.B(n_1107),
.Y(n_1305)
);

AO21x2_ASAP7_75t_L g1306 ( 
.A1(n_1087),
.A2(n_946),
.B(n_963),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1110),
.B(n_917),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1110),
.B(n_1104),
.Y(n_1308)
);

INVx3_ASAP7_75t_SL g1309 ( 
.A(n_1076),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1150),
.A2(n_1152),
.B(n_1151),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1070),
.A2(n_1018),
.B1(n_900),
.B2(n_982),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_L g1312 ( 
.A(n_1111),
.B(n_813),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1110),
.B(n_1104),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1041),
.A2(n_1055),
.A3(n_1039),
.B(n_1097),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1171),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1188),
.A2(n_1292),
.B1(n_1174),
.B2(n_1303),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1226),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1228),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1229),
.Y(n_1319)
);

AND2x6_ASAP7_75t_L g1320 ( 
.A(n_1221),
.B(n_1311),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1203),
.B(n_1206),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1204),
.B(n_1233),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1169),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1304),
.A2(n_1244),
.B(n_1310),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1206),
.B(n_1193),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1262),
.B(n_1307),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1182),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1209),
.A2(n_1313),
.B(n_1302),
.C(n_1308),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1239),
.A2(n_1176),
.B(n_1175),
.Y(n_1329)
);

AO221x2_ASAP7_75t_L g1330 ( 
.A1(n_1303),
.A2(n_1179),
.B1(n_1174),
.B2(n_1192),
.C(n_1298),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1226),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1262),
.B(n_1186),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1300),
.A2(n_1312),
.B1(n_1311),
.B2(n_1215),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1189),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1192),
.A2(n_1289),
.B(n_1195),
.C(n_1301),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1198),
.A2(n_1299),
.B1(n_1286),
.B2(n_1181),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1205),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1178),
.A2(n_1227),
.B(n_1280),
.Y(n_1338)
);

AOI22x1_ASAP7_75t_L g1339 ( 
.A1(n_1298),
.A2(n_1304),
.B1(n_1257),
.B2(n_1287),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1170),
.A2(n_1201),
.B(n_1212),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1196),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1203),
.B(n_1216),
.Y(n_1342)
);

INVx8_ASAP7_75t_L g1343 ( 
.A(n_1216),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1183),
.A2(n_1190),
.B(n_1268),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1234),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1220),
.A2(n_1187),
.B(n_1190),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1284),
.A2(n_1177),
.B(n_1180),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1225),
.A2(n_1243),
.A3(n_1249),
.B(n_1199),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1285),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1177),
.A2(n_1180),
.B(n_1183),
.Y(n_1350)
);

OR2x6_ASAP7_75t_L g1351 ( 
.A(n_1290),
.B(n_1203),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1270),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1218),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1173),
.B(n_1214),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1197),
.B(n_1194),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1274),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1208),
.A2(n_1202),
.B(n_1207),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1221),
.A2(n_1290),
.B1(n_1184),
.B2(n_1289),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1181),
.A2(n_1242),
.B1(n_1253),
.B2(n_1306),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1217),
.A2(n_1231),
.B(n_1237),
.Y(n_1360)
);

BUFx8_ASAP7_75t_SL g1361 ( 
.A(n_1211),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1281),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1265),
.A2(n_1271),
.B1(n_1246),
.B2(n_1276),
.Y(n_1363)
);

CKINVDCx8_ASAP7_75t_R g1364 ( 
.A(n_1226),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1219),
.B(n_1279),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1251),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1191),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1216),
.B(n_1297),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1235),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1222),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_SL g1371 ( 
.A1(n_1305),
.A2(n_1296),
.B(n_1276),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1271),
.B(n_1267),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1294),
.Y(n_1373)
);

AOI22x1_ASAP7_75t_L g1374 ( 
.A1(n_1257),
.A2(n_1282),
.B1(n_1283),
.B2(n_1275),
.Y(n_1374)
);

OAI222xp33_ASAP7_75t_L g1375 ( 
.A1(n_1263),
.A2(n_1248),
.B1(n_1293),
.B2(n_1238),
.C1(n_1259),
.C2(n_1230),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1235),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1237),
.A2(n_1236),
.B(n_1231),
.Y(n_1377)
);

AOI221xp5_ASAP7_75t_L g1378 ( 
.A1(n_1230),
.A2(n_1258),
.B1(n_1240),
.B2(n_1223),
.C(n_1291),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1200),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1200),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1241),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1309),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1185),
.A2(n_1314),
.A3(n_1264),
.B(n_1261),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1240),
.A2(n_1194),
.B1(n_1269),
.B2(n_1272),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1295),
.A2(n_1273),
.B(n_1236),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1255),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1193),
.B(n_1255),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_SL g1388 ( 
.A1(n_1254),
.A2(n_1232),
.B(n_1260),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1288),
.B(n_1278),
.Y(n_1389)
);

AOI21xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1210),
.A2(n_1252),
.B(n_1247),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1255),
.B(n_1256),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1241),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1185),
.A2(n_1314),
.A3(n_1172),
.B(n_1266),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1185),
.A2(n_1314),
.B(n_1172),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1252),
.A2(n_1256),
.B(n_1224),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1256),
.B(n_1213),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1241),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1277),
.B(n_1172),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1250),
.A2(n_1247),
.B(n_1245),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1245),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1250),
.A2(n_1245),
.B(n_1247),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1250),
.B(n_1018),
.Y(n_1402)
);

OAI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1311),
.A2(n_982),
.B1(n_1018),
.B2(n_848),
.C(n_917),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1304),
.A2(n_1190),
.B(n_1087),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1174),
.A2(n_1114),
.B1(n_982),
.B2(n_1082),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1193),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1310),
.A2(n_1239),
.B(n_1244),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1210),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1311),
.A2(n_1018),
.B(n_982),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1309),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1211),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1171),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1304),
.A2(n_1244),
.B(n_1087),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1302),
.B(n_1308),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1304),
.A2(n_1244),
.B(n_1087),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1307),
.A2(n_917),
.B1(n_1018),
.B2(n_982),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1310),
.A2(n_1239),
.B(n_1244),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1304),
.A2(n_1244),
.B(n_1087),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1169),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1285),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1171),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1171),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1174),
.A2(n_1114),
.B1(n_982),
.B2(n_1082),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1311),
.A2(n_1018),
.B(n_982),
.Y(n_1429)
);

BUFx2_ASAP7_75t_R g1430 ( 
.A(n_1309),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_SL g1431 ( 
.A(n_1216),
.B(n_1203),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1171),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1304),
.A2(n_1190),
.B(n_1087),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1193),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1304),
.A2(n_1244),
.B(n_1087),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1285),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1171),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1171),
.Y(n_1439)
);

OAI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1311),
.A2(n_982),
.B1(n_1018),
.B2(n_848),
.C(n_917),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1262),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1302),
.B(n_1308),
.Y(n_1442)
);

INVxp33_ASAP7_75t_L g1443 ( 
.A(n_1299),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1307),
.B(n_1018),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1171),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1302),
.B(n_1308),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1196),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1171),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1262),
.B(n_1307),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1196),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1310),
.A2(n_1244),
.B(n_1239),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1302),
.B(n_1308),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1171),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1171),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1364),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1444),
.A2(n_1429),
.B(n_1411),
.C(n_1403),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1332),
.B(n_1326),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1406),
.A2(n_1428),
.B1(n_1440),
.B2(n_1420),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1406),
.A2(n_1428),
.B1(n_1443),
.B2(n_1444),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1322),
.B(n_1372),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1342),
.B(n_1321),
.Y(n_1463)
);

O2A1O1Ixp5_ASAP7_75t_L g1464 ( 
.A1(n_1402),
.A2(n_1375),
.B(n_1357),
.C(n_1340),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1341),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1328),
.A2(n_1442),
.B(n_1417),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1443),
.A2(n_1333),
.B1(n_1454),
.B2(n_1447),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1335),
.A2(n_1358),
.B(n_1366),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1336),
.A2(n_1316),
.B1(n_1363),
.B2(n_1384),
.Y(n_1469)
);

AOI21x1_ASAP7_75t_SL g1470 ( 
.A1(n_1398),
.A2(n_1355),
.B(n_1354),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1441),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1336),
.A2(n_1363),
.B1(n_1384),
.B2(n_1359),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1370),
.B(n_1402),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1342),
.B(n_1368),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1451),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1341),
.Y(n_1476)
);

AOI211xp5_ASAP7_75t_L g1477 ( 
.A1(n_1390),
.A2(n_1378),
.B(n_1373),
.C(n_1437),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1370),
.B(n_1330),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1323),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1382),
.B(n_1412),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1368),
.B(n_1431),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1346),
.A2(n_1360),
.B(n_1399),
.Y(n_1482)
);

O2A1O1Ixp5_ASAP7_75t_L g1483 ( 
.A1(n_1381),
.A2(n_1392),
.B(n_1400),
.C(n_1397),
.Y(n_1483)
);

AOI221x1_ASAP7_75t_SL g1484 ( 
.A1(n_1327),
.A2(n_1345),
.B1(n_1337),
.B2(n_1334),
.C(n_1456),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1330),
.B(n_1376),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1330),
.B(n_1351),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1359),
.A2(n_1339),
.B1(n_1424),
.B2(n_1349),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1369),
.B(n_1320),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1423),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1368),
.B(n_1351),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1351),
.A2(n_1365),
.B1(n_1325),
.B2(n_1374),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1318),
.B(n_1425),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1360),
.A2(n_1338),
.B(n_1329),
.Y(n_1493)
);

AOI21x1_ASAP7_75t_SL g1494 ( 
.A1(n_1367),
.A2(n_1389),
.B(n_1396),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1438),
.B(n_1446),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1387),
.A2(n_1404),
.B(n_1434),
.Y(n_1496)
);

A2O1A1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1377),
.A2(n_1350),
.B(n_1347),
.C(n_1343),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1315),
.A2(n_1427),
.B1(n_1319),
.B2(n_1414),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1371),
.B(n_1395),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1391),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1449),
.B(n_1455),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1353),
.Y(n_1502)
);

AOI21x1_ASAP7_75t_SL g1503 ( 
.A1(n_1385),
.A2(n_1388),
.B(n_1320),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1433),
.A2(n_1439),
.B1(n_1430),
.B2(n_1448),
.Y(n_1504)
);

AOI21x1_ASAP7_75t_SL g1505 ( 
.A1(n_1320),
.A2(n_1393),
.B(n_1348),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1452),
.A2(n_1356),
.B1(n_1362),
.B2(n_1352),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1369),
.B(n_1320),
.Y(n_1507)
);

BUFx4f_ASAP7_75t_SL g1508 ( 
.A(n_1410),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1352),
.A2(n_1362),
.B(n_1380),
.C(n_1379),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1338),
.A2(n_1329),
.B(n_1401),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1320),
.B(n_1350),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1407),
.A2(n_1435),
.B1(n_1410),
.B2(n_1331),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1407),
.B(n_1435),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1317),
.A2(n_1386),
.B1(n_1331),
.B2(n_1413),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1317),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_R g1516 ( 
.A(n_1413),
.B(n_1331),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1404),
.B(n_1434),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1386),
.B(n_1394),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1394),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1394),
.B(n_1393),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1361),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1393),
.B(n_1383),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1393),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1383),
.B(n_1348),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1383),
.B(n_1344),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1344),
.B(n_1383),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1344),
.A2(n_1418),
.B1(n_1416),
.B2(n_1422),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1348),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1348),
.B(n_1436),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1418),
.B(n_1324),
.Y(n_1530)
);

AOI21x1_ASAP7_75t_SL g1531 ( 
.A1(n_1324),
.A2(n_1421),
.B(n_1408),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1405),
.A2(n_1426),
.B(n_1409),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1405),
.B(n_1426),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1409),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1453),
.B(n_1415),
.Y(n_1535)
);

AOI211xp5_ASAP7_75t_L g1536 ( 
.A1(n_1415),
.A2(n_1419),
.B(n_1432),
.C(n_1445),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1432),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1445),
.A2(n_1450),
.B(n_1453),
.C(n_1361),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1450),
.B(n_1328),
.Y(n_1539)
);

CKINVDCx6p67_ASAP7_75t_R g1540 ( 
.A(n_1410),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1322),
.B(n_1372),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1328),
.B(n_1370),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1332),
.B(n_1326),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1441),
.Y(n_1544)
);

CKINVDCx12_ASAP7_75t_R g1545 ( 
.A(n_1332),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1406),
.A2(n_982),
.B1(n_917),
.B2(n_1428),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1322),
.B(n_1372),
.Y(n_1547)
);

NOR2xp67_ASAP7_75t_L g1548 ( 
.A(n_1326),
.B(n_1214),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1322),
.B(n_1372),
.Y(n_1549)
);

O2A1O1Ixp5_ASAP7_75t_L g1550 ( 
.A1(n_1411),
.A2(n_1429),
.B(n_1402),
.C(n_1018),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1441),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1406),
.A2(n_982),
.B1(n_917),
.B2(n_1428),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1403),
.A2(n_1018),
.B(n_1440),
.C(n_1429),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1322),
.B(n_1372),
.Y(n_1554)
);

O2A1O1Ixp5_ASAP7_75t_L g1555 ( 
.A1(n_1411),
.A2(n_1429),
.B(n_1402),
.C(n_1018),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1328),
.B(n_1370),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1328),
.B(n_1370),
.Y(n_1557)
);

O2A1O1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1403),
.A2(n_1018),
.B(n_1440),
.C(n_1429),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1342),
.B(n_1321),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1322),
.B(n_1372),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1382),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1406),
.A2(n_982),
.B1(n_917),
.B2(n_1428),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1441),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1322),
.B(n_1372),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1332),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1328),
.B(n_1370),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1518),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1490),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1509),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1509),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1553),
.A2(n_1558),
.B(n_1555),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1533),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1517),
.B(n_1525),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1519),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1565),
.B(n_1475),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1459),
.B(n_1543),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1517),
.B(n_1478),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1483),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1488),
.B(n_1507),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1478),
.B(n_1526),
.Y(n_1582)
);

NAND2x1p5_ASAP7_75t_L g1583 ( 
.A(n_1542),
.B(n_1566),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1545),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1499),
.B(n_1496),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1481),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1553),
.A2(n_1558),
.B(n_1550),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1488),
.B(n_1507),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_SL g1589 ( 
.A(n_1521),
.Y(n_1589)
);

AO21x1_ASAP7_75t_SL g1590 ( 
.A1(n_1542),
.A2(n_1566),
.B(n_1556),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1490),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1526),
.B(n_1528),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1510),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1486),
.B(n_1522),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1529),
.B(n_1556),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1535),
.A2(n_1527),
.B(n_1539),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1460),
.A2(n_1461),
.B1(n_1546),
.B2(n_1552),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1523),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1544),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1510),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1458),
.A2(n_1469),
.B(n_1562),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1499),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1464),
.A2(n_1530),
.B(n_1538),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1466),
.A2(n_1468),
.B(n_1467),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1506),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1463),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1557),
.B(n_1524),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1520),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1557),
.B(n_1524),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1492),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1482),
.B(n_1485),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1471),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1495),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1491),
.B(n_1472),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1501),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1485),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1484),
.Y(n_1618)
);

AOI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1537),
.A2(n_1534),
.B(n_1487),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1462),
.B(n_1554),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1541),
.B(n_1547),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1508),
.B(n_1551),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1548),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1500),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1493),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1563),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1498),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1532),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1489),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1479),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1474),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1576),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1574),
.B(n_1569),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1628),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1605),
.A2(n_1504),
.B1(n_1564),
.B2(n_1560),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1576),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1569),
.B(n_1536),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1598),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1573),
.B(n_1477),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1612),
.B(n_1549),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1603),
.B(n_1559),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1581),
.B(n_1588),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1580),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1625),
.A2(n_1531),
.B(n_1503),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1602),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1595),
.B(n_1513),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_SL g1647 ( 
.A1(n_1572),
.A2(n_1587),
.B1(n_1615),
.B2(n_1601),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1580),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1601),
.B(n_1512),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1585),
.B(n_1603),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1575),
.B(n_1582),
.Y(n_1651)
);

NOR4xp25_ASAP7_75t_SL g1652 ( 
.A(n_1602),
.B(n_1561),
.C(n_1494),
.D(n_1470),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1593),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1600),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1582),
.B(n_1514),
.Y(n_1655)
);

AOI211x1_ASAP7_75t_SL g1656 ( 
.A1(n_1597),
.A2(n_1480),
.B(n_1515),
.C(n_1465),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1583),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1595),
.B(n_1465),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1505),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1579),
.B(n_1617),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1583),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1592),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1647),
.A2(n_1618),
.B1(n_1597),
.B2(n_1617),
.C(n_1606),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1642),
.B(n_1624),
.Y(n_1664)
);

OAI33xp33_ASAP7_75t_L g1665 ( 
.A1(n_1639),
.A2(n_1579),
.A3(n_1577),
.B1(n_1627),
.B2(n_1578),
.B3(n_1610),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1633),
.B(n_1567),
.Y(n_1666)
);

OAI31xp33_ASAP7_75t_L g1667 ( 
.A1(n_1649),
.A2(n_1583),
.A3(n_1623),
.B(n_1603),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1649),
.A2(n_1615),
.B1(n_1639),
.B2(n_1650),
.Y(n_1668)
);

NOR4xp25_ASAP7_75t_SL g1669 ( 
.A(n_1657),
.B(n_1590),
.C(n_1568),
.D(n_1591),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1647),
.A2(n_1615),
.B1(n_1584),
.B2(n_1591),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1643),
.Y(n_1671)
);

OAI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1650),
.A2(n_1615),
.B1(n_1585),
.B2(n_1610),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1633),
.B(n_1642),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1632),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1635),
.A2(n_1615),
.B1(n_1568),
.B2(n_1631),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1635),
.A2(n_1631),
.B1(n_1608),
.B2(n_1607),
.Y(n_1676)
);

NAND2xp33_ASAP7_75t_R g1677 ( 
.A(n_1652),
.B(n_1516),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1634),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1643),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1633),
.B(n_1594),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1648),
.B(n_1604),
.C(n_1608),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1651),
.B(n_1596),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1655),
.A2(n_1626),
.B1(n_1585),
.B2(n_1627),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1636),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1648),
.Y(n_1685)
);

INVx5_ASAP7_75t_L g1686 ( 
.A(n_1650),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1638),
.Y(n_1687)
);

OAI33xp33_ASAP7_75t_L g1688 ( 
.A1(n_1660),
.A2(n_1614),
.A3(n_1616),
.B1(n_1611),
.B2(n_1570),
.B3(n_1571),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1585),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1637),
.A2(n_1613),
.B1(n_1630),
.B2(n_1629),
.C(n_1599),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1646),
.B(n_1611),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1657),
.A2(n_1619),
.B(n_1604),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1645),
.Y(n_1693)
);

OAI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1650),
.A2(n_1585),
.B1(n_1586),
.B2(n_1607),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1637),
.A2(n_1620),
.B1(n_1621),
.B2(n_1616),
.C(n_1614),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1640),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1658),
.B(n_1622),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1673),
.B(n_1637),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1667),
.B(n_1641),
.Y(n_1699)
);

OR2x6_ASAP7_75t_L g1700 ( 
.A(n_1681),
.B(n_1650),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1693),
.Y(n_1701)
);

OAI21xp33_ASAP7_75t_L g1702 ( 
.A1(n_1663),
.A2(n_1655),
.B(n_1659),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1671),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1690),
.B(n_1604),
.C(n_1652),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1684),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1684),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1682),
.B(n_1662),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1692),
.A2(n_1644),
.B(n_1625),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1678),
.A2(n_1654),
.B(n_1653),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1670),
.A2(n_1619),
.B(n_1661),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1693),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1687),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1679),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1693),
.B(n_1650),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1687),
.Y(n_1716)
);

NOR2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1664),
.B(n_1540),
.Y(n_1717)
);

INVxp67_ASAP7_75t_SL g1718 ( 
.A(n_1685),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1693),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1712),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1703),
.B(n_1674),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1700),
.B(n_1669),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1698),
.B(n_1696),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1704),
.A2(n_1668),
.B(n_1675),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1710),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1710),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1703),
.B(n_1718),
.Y(n_1727)
);

AOI22x1_ASAP7_75t_L g1728 ( 
.A1(n_1711),
.A2(n_1457),
.B1(n_1661),
.B2(n_1677),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1714),
.Y(n_1729)
);

INVx6_ASAP7_75t_L g1730 ( 
.A(n_1719),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1715),
.B(n_1686),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1714),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1715),
.B(n_1686),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1705),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1702),
.A2(n_1704),
.B1(n_1665),
.B2(n_1711),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1707),
.Y(n_1737)
);

AND4x1_ASAP7_75t_L g1738 ( 
.A(n_1702),
.B(n_1656),
.C(n_1676),
.D(n_1688),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1718),
.B(n_1698),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1710),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1698),
.B(n_1695),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1699),
.B(n_1694),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1719),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1706),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1715),
.B(n_1680),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1699),
.A2(n_1672),
.B1(n_1650),
.B2(n_1686),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1706),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1700),
.B(n_1693),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1713),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1700),
.B(n_1666),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1700),
.B(n_1666),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1713),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1707),
.A2(n_1683),
.B1(n_1697),
.B2(n_1502),
.C(n_1691),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1716),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1729),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1729),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1720),
.B(n_1707),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1720),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_SL g1761 ( 
.A(n_1728),
.B(n_1719),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1730),
.B(n_1719),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1701),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1720),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1730),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1736),
.B(n_1701),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1734),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1730),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1730),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1747),
.B(n_1719),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1734),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1738),
.B(n_1701),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1743),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1737),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1747),
.B(n_1712),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1723),
.B(n_1712),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1727),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1723),
.B(n_1712),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1738),
.B(n_1680),
.Y(n_1779)
);

NOR2xp67_ASAP7_75t_SL g1780 ( 
.A(n_1724),
.B(n_1730),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1739),
.B(n_1727),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1737),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1743),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1739),
.B(n_1708),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1746),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1732),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1746),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1731),
.B(n_1715),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1756),
.Y(n_1789)
);

NAND2x1p5_ASAP7_75t_L g1790 ( 
.A(n_1728),
.B(n_1709),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1742),
.B(n_1708),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1749),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1749),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1780),
.B(n_1724),
.C(n_1744),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1774),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1774),
.Y(n_1796)
);

BUFx2_ASAP7_75t_SL g1797 ( 
.A(n_1782),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1776),
.B(n_1745),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1786),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1757),
.B(n_1732),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1759),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1776),
.B(n_1745),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1777),
.B(n_1589),
.Y(n_1803)
);

INVx4_ASAP7_75t_L g1804 ( 
.A(n_1762),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1758),
.B(n_1742),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1772),
.A2(n_1755),
.B(n_1748),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1769),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1771),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1759),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1759),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1771),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1782),
.B(n_1721),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1778),
.B(n_1745),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1767),
.B(n_1721),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1778),
.B(n_1745),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_SL g1816 ( 
.A1(n_1779),
.A2(n_1761),
.B1(n_1763),
.B2(n_1766),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1775),
.B(n_1750),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1775),
.B(n_1750),
.Y(n_1818)
);

NOR3xp33_ASAP7_75t_L g1819 ( 
.A(n_1765),
.B(n_1722),
.C(n_1755),
.Y(n_1819)
);

OAI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1794),
.A2(n_1780),
.B1(n_1790),
.B2(n_1781),
.C(n_1765),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1817),
.B(n_1770),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1795),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1794),
.A2(n_1722),
.B1(n_1741),
.B2(n_1735),
.C1(n_1750),
.C2(n_1788),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1795),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1817),
.B(n_1770),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1816),
.A2(n_1790),
.B(n_1722),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1819),
.A2(n_1788),
.B1(n_1733),
.B2(n_1731),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1807),
.B(n_1781),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1803),
.B(n_1768),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1816),
.A2(n_1790),
.B(n_1733),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1818),
.B(n_1768),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1818),
.B(n_1762),
.Y(n_1832)
);

AOI21xp33_ASAP7_75t_SL g1833 ( 
.A1(n_1805),
.A2(n_1762),
.B(n_1791),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1796),
.Y(n_1834)
);

OAI222xp33_ASAP7_75t_L g1835 ( 
.A1(n_1806),
.A2(n_1700),
.B1(n_1762),
.B2(n_1791),
.C1(n_1735),
.C2(n_1741),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1806),
.A2(n_1735),
.B(n_1741),
.C(n_1731),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1807),
.A2(n_1733),
.B1(n_1731),
.B2(n_1715),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1796),
.B(n_1760),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1795),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1801),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1825),
.B(n_1798),
.Y(n_1841)
);

NAND2xp33_ASAP7_75t_R g1842 ( 
.A(n_1824),
.B(n_1799),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1840),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_R g1844 ( 
.A(n_1834),
.B(n_1799),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1825),
.B(n_1815),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1826),
.B(n_1804),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1840),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1831),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1821),
.B(n_1815),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1820),
.A2(n_1733),
.B1(n_1797),
.B2(n_1805),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1822),
.Y(n_1851)
);

O2A1O1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1846),
.A2(n_1830),
.B(n_1836),
.C(n_1833),
.Y(n_1852)
);

AOI21xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1842),
.A2(n_1828),
.B(n_1829),
.Y(n_1853)
);

OAI211xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1850),
.A2(n_1836),
.B(n_1827),
.C(n_1823),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1844),
.A2(n_1835),
.B1(n_1800),
.B2(n_1797),
.C(n_1838),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1841),
.B(n_1822),
.Y(n_1856)
);

AOI211xp5_ASAP7_75t_SL g1857 ( 
.A1(n_1848),
.A2(n_1829),
.B(n_1839),
.C(n_1800),
.Y(n_1857)
);

NOR4xp25_ASAP7_75t_L g1858 ( 
.A(n_1847),
.B(n_1839),
.C(n_1808),
.D(n_1811),
.Y(n_1858)
);

AOI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1849),
.A2(n_1814),
.B1(n_1812),
.B2(n_1808),
.C(n_1811),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1841),
.B(n_1801),
.Y(n_1860)
);

OAI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1851),
.A2(n_1837),
.B1(n_1804),
.B2(n_1814),
.C(n_1812),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1852),
.A2(n_1847),
.B(n_1843),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1856),
.Y(n_1863)
);

AOI222xp33_ASAP7_75t_L g1864 ( 
.A1(n_1855),
.A2(n_1845),
.B1(n_1849),
.B2(n_1843),
.C1(n_1832),
.C2(n_1804),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1860),
.Y(n_1865)
);

A2O1A1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1853),
.A2(n_1845),
.B(n_1832),
.C(n_1809),
.Y(n_1866)
);

AOI22x1_ASAP7_75t_L g1867 ( 
.A1(n_1857),
.A2(n_1804),
.B1(n_1810),
.B2(n_1809),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1867),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1863),
.B(n_1861),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1865),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1866),
.B(n_1858),
.Y(n_1871)
);

NAND3xp33_ASAP7_75t_L g1872 ( 
.A(n_1864),
.B(n_1854),
.C(n_1859),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1862),
.A2(n_1809),
.B(n_1801),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1866),
.B(n_1798),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1868),
.B(n_1810),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1873),
.B(n_1810),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1872),
.A2(n_1869),
.B1(n_1874),
.B2(n_1871),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1870),
.A2(n_1813),
.B1(n_1802),
.B2(n_1760),
.Y(n_1878)
);

OAI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1872),
.A2(n_1764),
.B1(n_1813),
.B2(n_1802),
.C(n_1773),
.Y(n_1879)
);

AOI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1872),
.A2(n_1764),
.B1(n_1792),
.B2(n_1789),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1875),
.B(n_1783),
.Y(n_1881)
);

XNOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1877),
.B(n_1717),
.Y(n_1882)
);

AO22x2_ASAP7_75t_L g1883 ( 
.A1(n_1876),
.A2(n_1787),
.B1(n_1793),
.B2(n_1785),
.Y(n_1883)
);

AOI32xp33_ASAP7_75t_L g1884 ( 
.A1(n_1882),
.A2(n_1878),
.A3(n_1879),
.B1(n_1880),
.B2(n_1793),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1884),
.A2(n_1881),
.B1(n_1883),
.B2(n_1773),
.C(n_1785),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1885),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1885),
.A2(n_1457),
.B1(n_1476),
.B2(n_1465),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1886),
.A2(n_1784),
.B1(n_1752),
.B2(n_1753),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1887),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1889),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1888),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1891),
.Y(n_1892)
);

AOI21xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1892),
.A2(n_1890),
.B(n_1784),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1893),
.A2(n_1752),
.B1(n_1753),
.B2(n_1756),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1894),
.Y(n_1895)
);

OA22x2_ASAP7_75t_L g1896 ( 
.A1(n_1895),
.A2(n_1726),
.B1(n_1725),
.B2(n_1740),
.Y(n_1896)
);

AOI211xp5_ASAP7_75t_L g1897 ( 
.A1(n_1896),
.A2(n_1476),
.B(n_1751),
.C(n_1754),
.Y(n_1897)
);


endmodule