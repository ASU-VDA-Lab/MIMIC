module fake_jpeg_21621_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_45),
.B(n_58),
.Y(n_132)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_33),
.CON(n_46),
.SN(n_46)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_54),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_55),
.B(n_75),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx12f_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_22),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_19),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_60),
.B(n_21),
.Y(n_144)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_1),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_17),
.B(n_14),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_67),
.B(n_39),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_1),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_3),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_4),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_86),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_30),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_40),
.B1(n_43),
.B2(n_24),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_92),
.A2(n_95),
.B1(n_122),
.B2(n_15),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_90),
.A2(n_40),
.B1(n_43),
.B2(n_24),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_40),
.B1(n_32),
.B2(n_29),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_27),
.B1(n_26),
.B2(n_83),
.Y(n_162)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_118),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_115),
.B(n_137),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_52),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_36),
.B1(n_32),
.B2(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_52),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_51),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_143),
.Y(n_182)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_SL g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_64),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_151),
.Y(n_206)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_60),
.C(n_61),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_148),
.B(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_63),
.B1(n_74),
.B2(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_150),
.A2(n_166),
.B1(n_116),
.B2(n_139),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_153),
.A2(n_179),
.B1(n_124),
.B2(n_96),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_46),
.A3(n_55),
.B1(n_35),
.B2(n_39),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_163),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_172),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_112),
.B(n_120),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_36),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_160),
.B(n_167),
.Y(n_218)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_79),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_170),
.Y(n_195)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_95),
.A2(n_47),
.B1(n_73),
.B2(n_76),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_132),
.B(n_27),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_84),
.B(n_85),
.C(n_91),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_168),
.A2(n_5),
.B(n_6),
.C(n_10),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_106),
.A2(n_82),
.B1(n_80),
.B2(n_72),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_169),
.A2(n_116),
.B1(n_114),
.B2(n_129),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_15),
.Y(n_170)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_38),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_106),
.A2(n_15),
.B1(n_38),
.B2(n_35),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_4),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_183),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_103),
.B(n_4),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_105),
.B(n_4),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_184),
.B(n_187),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_108),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_124),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_111),
.A2(n_52),
.B1(n_6),
.B2(n_9),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_119),
.B1(n_97),
.B2(n_101),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_100),
.B(n_5),
.CI(n_6),
.CON(n_190),
.SN(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_108),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_205),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_129),
.B1(n_111),
.B2(n_112),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_202),
.A2(n_213),
.B(n_156),
.C(n_177),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_186),
.B(n_163),
.Y(n_234)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_214),
.B1(n_217),
.B2(n_220),
.Y(n_230)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_165),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_168),
.A2(n_109),
.B1(n_128),
.B2(n_141),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_134),
.B1(n_130),
.B2(n_109),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_159),
.A2(n_170),
.B(n_190),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_184),
.B(n_175),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_155),
.A2(n_117),
.B1(n_108),
.B2(n_9),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_228),
.B1(n_189),
.B2(n_150),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_172),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_174),
.B(n_5),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_190),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_192),
.B1(n_221),
.B2(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_231),
.A2(n_243),
.B1(n_259),
.B2(n_229),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_232),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_233),
.B(n_239),
.Y(n_265)
);

OAI21x1_ASAP7_75t_SL g276 ( 
.A1(n_234),
.A2(n_239),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_236),
.A2(n_261),
.B1(n_199),
.B2(n_219),
.Y(n_267)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_192),
.C(n_148),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_242),
.C(n_258),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_183),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_195),
.C(n_212),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_209),
.B1(n_195),
.B2(n_153),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_152),
.A3(n_149),
.B1(n_180),
.B2(n_166),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_246),
.A2(n_222),
.B(n_226),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_249),
.B(n_218),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_182),
.B(n_158),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_193),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_216),
.B(n_173),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_255),
.Y(n_266)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_171),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_260),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_194),
.C(n_208),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_225),
.A2(n_188),
.B1(n_187),
.B2(n_178),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_200),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_220),
.A2(n_147),
.B1(n_181),
.B2(n_161),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_273),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_267),
.A2(n_272),
.B1(n_278),
.B2(n_257),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_206),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_275),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_214),
.B1(n_200),
.B2(n_229),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_218),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_247),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_226),
.B(n_211),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_245),
.B(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_230),
.A2(n_199),
.B1(n_210),
.B2(n_205),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_231),
.B(n_215),
.CI(n_226),
.CON(n_279),
.SN(n_279)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_279),
.B(n_273),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_235),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_233),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_246),
.B(n_259),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_215),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_289),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_222),
.B1(n_211),
.B2(n_157),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_261),
.B1(n_230),
.B2(n_255),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_204),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_249),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_238),
.C(n_251),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_291),
.A2(n_303),
.B(n_305),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_311),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_282),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_262),
.B(n_265),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_297),
.A2(n_284),
.B(n_274),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_267),
.B1(n_272),
.B2(n_278),
.Y(n_319)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_301),
.Y(n_327)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_304),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_314),
.B1(n_315),
.B2(n_266),
.Y(n_328)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_247),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_285),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_260),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_287),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_317),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_319),
.A2(n_322),
.B1(n_293),
.B2(n_297),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_262),
.B1(n_279),
.B2(n_246),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_303),
.A2(n_279),
.B1(n_246),
.B2(n_266),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_332),
.B1(n_294),
.B2(n_305),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_282),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_330),
.C(n_334),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_336),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_270),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_315),
.A2(n_246),
.B1(n_277),
.B2(n_250),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_290),
.C(n_263),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_276),
.C(n_274),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_337),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_284),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_351),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_336),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_319),
.A2(n_293),
.B1(n_314),
.B2(n_294),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_342),
.A2(n_346),
.B1(n_349),
.B2(n_325),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_311),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_344),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_335),
.B(n_291),
.CI(n_306),
.CON(n_344),
.SN(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_345),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_322),
.A2(n_313),
.B1(n_310),
.B2(n_309),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_332),
.A2(n_323),
.B1(n_320),
.B2(n_324),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_299),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_350),
.A2(n_337),
.B(n_318),
.Y(n_365)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_321),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_354),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_304),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_312),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

BUFx12f_ASAP7_75t_SL g360 ( 
.A(n_344),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_360),
.A2(n_363),
.B(n_353),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_366),
.Y(n_376)
);

A2O1A1O1Ixp25_ASAP7_75t_L g363 ( 
.A1(n_344),
.A2(n_325),
.B(n_316),
.C(n_330),
.D(n_326),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_367),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_355),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_338),
.Y(n_367)
);

AOI22x1_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_317),
.B1(n_308),
.B2(n_301),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_368),
.A2(n_349),
.B1(n_339),
.B2(n_340),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_292),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_347),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_368),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_372),
.B(n_380),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_358),
.A2(n_346),
.B1(n_342),
.B2(n_343),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_373),
.A2(n_253),
.B1(n_237),
.B2(n_196),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_292),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_378),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_363),
.Y(n_387)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_362),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_356),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_347),
.C(n_351),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_376),
.A2(n_359),
.B(n_364),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_381),
.A2(n_386),
.B(n_377),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_383),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g386 ( 
.A(n_376),
.B(n_367),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_11),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_388),
.A2(n_375),
.B1(n_377),
.B2(n_371),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_380),
.B(n_5),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_389),
.B(n_6),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_370),
.C(n_371),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_392),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_393),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_373),
.Y(n_392)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_394),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_395),
.A2(n_381),
.B(n_388),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_400),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_399),
.A2(n_396),
.B(n_392),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_402),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_387),
.C(n_383),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_397),
.Y(n_404)
);

OAI321xp33_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_157),
.C(n_176),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_405),
.B(n_12),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_12),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_13),
.Y(n_409)
);


endmodule