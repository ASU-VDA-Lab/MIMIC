module real_jpeg_2244_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_39),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_1),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_1),
.B(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_1),
.B(n_27),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_3),
.B(n_45),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_3),
.B(n_78),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_3),
.B(n_50),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_3),
.B(n_106),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_3),
.B(n_36),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_4),
.B(n_27),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_4),
.B(n_32),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_4),
.B(n_39),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_4),
.B(n_45),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_4),
.B(n_50),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_5),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_5),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_5),
.B(n_45),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_5),
.B(n_78),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_5),
.B(n_50),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_6),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_6),
.B(n_78),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_6),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_8),
.B(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_8),
.B(n_39),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_8),
.B(n_45),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_8),
.B(n_32),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_8),
.B(n_50),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_78),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_8),
.B(n_106),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_8),
.B(n_36),
.Y(n_305)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_13),
.B(n_32),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_13),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_13),
.B(n_27),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_13),
.B(n_39),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_13),
.B(n_45),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_14),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_14),
.B(n_78),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_14),
.B(n_106),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_19),
.B(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.C(n_81),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_20),
.A2(n_21),
.B1(n_61),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_42),
.B2(n_60),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_22),
.B(n_43),
.C(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_31),
.C(n_34),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_25),
.A2(n_26),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_25),
.A2(n_26),
.B1(n_107),
.B2(n_360),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_26),
.B(n_101),
.C(n_107),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_26),
.B(n_331),
.C(n_334),
.Y(n_356)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_27),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.C(n_40),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_35),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_35),
.Y(n_98)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_36),
.Y(n_145)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_38),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_38),
.A2(n_97),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_38),
.B(n_297),
.C(n_301),
.Y(n_331)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_39),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_52),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.C(n_51),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_44),
.A2(n_55),
.B1(n_89),
.B2(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_44),
.B(n_89),
.C(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_45),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_74),
.C(n_76),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_49),
.B1(n_76),
.B2(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_48),
.A2(n_49),
.B1(n_168),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_49),
.B(n_168),
.C(n_169),
.Y(n_167)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_50),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_57),
.C(n_58),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_56),
.A2(n_57),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_56),
.A2(n_57),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_57),
.B(n_70),
.C(n_197),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_61),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.C(n_73),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_62),
.A2(n_63),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_65),
.B(n_73),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.C(n_71),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_92),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_67),
.B(n_153),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_69),
.A2(n_70),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_75),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_76),
.A2(n_77),
.B1(n_207),
.B2(n_210),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_76),
.A2(n_77),
.B1(n_105),
.B2(n_231),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_103),
.C(n_105),
.Y(n_102)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_79),
.B(n_212),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_81),
.B(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_95),
.C(n_100),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_82),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_91),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_83),
.A2(n_84),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_87),
.B(n_91),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_88),
.B(n_90),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_89),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_89),
.A2(n_147),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_95),
.B(n_100),
.Y(n_379)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_101),
.A2(n_102),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_103),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_103),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_105),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_105),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_105),
.A2(n_135),
.B1(n_165),
.B2(n_231),
.Y(n_304)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_106),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_107),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_122),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_120),
.A2(n_121),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_121),
.B(n_317),
.C(n_318),
.Y(n_329)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_372),
.B(n_387),
.Y(n_125)
);

OAI31xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_321),
.A3(n_361),
.B(n_366),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_289),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_213),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_181),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_130),
.B(n_181),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_148),
.C(n_171),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_131),
.B(n_286),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_131),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_138),
.CI(n_142),
.CON(n_131),
.SN(n_131)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_132),
.B(n_138),
.C(n_142),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_137),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_133),
.A2(n_134),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_134),
.A2(n_165),
.B(n_231),
.C(n_305),
.Y(n_344)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_162),
.B1(n_165),
.B2(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_136),
.B(n_137),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_141),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_141),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_144),
.B(n_163),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_144),
.B(n_192),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_148),
.B(n_171),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_159),
.B2(n_170),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_160),
.C(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_156),
.C(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_155),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_167),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_164),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_168),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_179),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_172),
.B(n_175),
.CI(n_179),
.CON(n_276),
.SN(n_276)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_178),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_224),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_181),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_199),
.CI(n_200),
.CON(n_181),
.SN(n_181)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_182),
.B(n_199),
.C(n_200),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_183),
.B(n_186),
.C(n_193),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_193),
.B2(n_194),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_187),
.B(n_189),
.C(n_191),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_197),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_202),
.B(n_203),
.C(n_205),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_207),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_284),
.B(n_288),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_272),
.B(n_283),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_244),
.B(n_271),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_235),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_235),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_227),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.C(n_222),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_221),
.CI(n_222),
.CON(n_236),
.SN(n_236)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_225),
.C(n_227),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_233),
.C(n_234),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.C(n_243),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_268),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_236),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_238),
.B1(n_243),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_265),
.B(n_270),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_256),
.B(n_264),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_252),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_259),
.B(n_263),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_261),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_274),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_279),
.C(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_276),
.Y(n_392)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_290),
.A2(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_320),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_291),
.B(n_320),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_292),
.B(n_294),
.C(n_307),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_306),
.B2(n_307),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_295),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_302),
.CI(n_303),
.CON(n_295),
.SN(n_295)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_302),
.C(n_303),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_312),
.C(n_313),
.Y(n_336)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g366 ( 
.A1(n_322),
.A2(n_362),
.B(n_367),
.C(n_370),
.D(n_371),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_348),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_323),
.B(n_348),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_336),
.C(n_337),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_325),
.B1(n_337),
.B2(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_335),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_329),
.C(n_330),
.Y(n_349)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_344),
.C(n_345),
.Y(n_355)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_346),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_351),
.C(n_354),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_354),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_356),
.CI(n_357),
.CON(n_354),
.SN(n_354)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_356),
.C(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_365),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_384),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_373),
.A2(n_388),
.B(n_389),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_377),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_377),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.C(n_383),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g385 ( 
.A(n_378),
.B(n_380),
.CI(n_383),
.CON(n_385),
.SN(n_385)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_381),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_386),
.Y(n_388)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_385),
.Y(n_394)
);


endmodule