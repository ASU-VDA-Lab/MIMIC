module fake_jpeg_26232_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_38),
.Y(n_69)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_32),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_18),
.B1(n_17),
.B2(n_32),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_53)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_40),
.B1(n_37),
.B2(n_41),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_18),
.B1(n_30),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_19),
.B1(n_30),
.B2(n_29),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_28),
.B1(n_19),
.B2(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_44),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_66),
.B1(n_36),
.B2(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_42),
.Y(n_64)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_41),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_75),
.Y(n_95)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_22),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_40),
.C(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_85),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_89),
.B1(n_57),
.B2(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_27),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_47),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_43),
.B1(n_37),
.B2(n_40),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_66),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_61),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_73),
.B(n_91),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_69),
.C(n_47),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_73),
.Y(n_122)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_106),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_50),
.B(n_67),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_76),
.B(n_97),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_105),
.Y(n_130)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_112),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_53),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_117),
.B(n_125),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_95),
.B(n_110),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_132),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_126),
.B1(n_131),
.B2(n_138),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_124),
.A2(n_25),
.B(n_16),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_70),
.B1(n_76),
.B2(n_85),
.Y(n_126)
);

OAI22x1_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_81),
.B1(n_80),
.B2(n_53),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_115),
.B(n_74),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_82),
.B1(n_79),
.B2(n_53),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_79),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_77),
.B1(n_62),
.B2(n_63),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_74),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_141),
.B(n_142),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_151),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_122),
.C(n_119),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_148),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_109),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_109),
.B(n_95),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_152),
.B(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_95),
.B(n_110),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_112),
.C(n_98),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_164),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_158),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_106),
.C(n_96),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_106),
.B1(n_100),
.B2(n_115),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_77),
.B1(n_140),
.B2(n_104),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_105),
.B(n_111),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_160),
.B(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_24),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_131),
.B1(n_136),
.B2(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_169),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_177),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_134),
.B1(n_129),
.B2(n_135),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_183),
.B1(n_187),
.B2(n_143),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_176),
.B1(n_181),
.B2(n_62),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_104),
.B1(n_93),
.B2(n_114),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_157),
.Y(n_177)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_178),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_25),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_165),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_42),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_188),
.B(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_93),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_192),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_165),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_204),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_147),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_148),
.C(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_201),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_152),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_202),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_144),
.C(n_146),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_143),
.C(n_161),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_64),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_62),
.B1(n_54),
.B2(n_46),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_46),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_208),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_185),
.B1(n_188),
.B2(n_167),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_184),
.B(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_68),
.C(n_54),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_40),
.B1(n_24),
.B2(n_16),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_168),
.B1(n_181),
.B2(n_167),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_214),
.B(n_226),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_174),
.B(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_208),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_183),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_201),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_168),
.B(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_68),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_0),
.B(n_1),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_228),
.B(n_1),
.Y(n_230)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_240),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_213),
.A2(n_220),
.B1(n_207),
.B2(n_216),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_238),
.B1(n_215),
.B2(n_3),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_198),
.C(n_205),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_235),
.C(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_227),
.C(n_225),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_211),
.B1(n_3),
.B2(n_4),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_211),
.C(n_42),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_2),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_223),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_235),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_236),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_248),
.B(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_25),
.C(n_26),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_2),
.B(n_4),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_5),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_229),
.B1(n_239),
.B2(n_234),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_232),
.C(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_244),
.C(n_251),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_248),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_5),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_5),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_26),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_258),
.A3(n_253),
.B1(n_255),
.B2(n_26),
.C1(n_14),
.C2(n_6),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_269),
.B(n_263),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_7),
.A3(n_10),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_261),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_271),
.B(n_268),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_13),
.B(n_15),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_13),
.Y(n_274)
);


endmodule