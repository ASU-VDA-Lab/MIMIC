module fake_jpeg_15085_n_163 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_33),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_18),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_21),
.C(n_27),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_20),
.C(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_15),
.B(n_2),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_16),
.A2(n_18),
.B1(n_25),
.B2(n_14),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_16),
.B(n_6),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_6),
.Y(n_70)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_7),
.B1(n_8),
.B2(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_66),
.B(n_70),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_7),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_76),
.C(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_19),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_89),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_32),
.B1(n_44),
.B2(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_35),
.C(n_32),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_90),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_19),
.C(n_8),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_95),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_9),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_97),
.Y(n_116)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_101),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_68),
.C(n_67),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_52),
.C(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_79),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_106),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_96),
.B1(n_94),
.B2(n_99),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_59),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_117),
.B1(n_118),
.B2(n_115),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_52),
.C(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_79),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_125),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_83),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_123),
.C(n_129),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.C(n_107),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_81),
.B1(n_88),
.B2(n_101),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_97),
.B1(n_95),
.B2(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_131),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_114),
.B(n_102),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_90),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_60),
.B1(n_78),
.B2(n_63),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_67),
.B1(n_98),
.B2(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_104),
.B1(n_117),
.B2(n_105),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_143),
.B1(n_124),
.B2(n_128),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_140),
.C(n_121),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_129),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_142),
.C(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_139),
.A2(n_125),
.B1(n_126),
.B2(n_132),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_150),
.B1(n_138),
.B2(n_135),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_136),
.B1(n_135),
.B2(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_155),
.C(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_154),
.B1(n_148),
.B2(n_145),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_127),
.A3(n_144),
.B1(n_151),
.B2(n_152),
.C1(n_156),
.C2(n_162),
.Y(n_163)
);


endmodule