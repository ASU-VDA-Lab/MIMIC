module fake_netlist_1_7582_n_934 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_934);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_934;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_285;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_504;
wire n_170;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g109 ( .A(n_21), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_11), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_41), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_71), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_94), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_97), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_6), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_58), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_57), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_42), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_31), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_4), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_8), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_65), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_5), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_90), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g129 ( .A(n_20), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_40), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_35), .Y(n_131) );
INVx1_ASAP7_75t_SL g132 ( .A(n_2), .Y(n_132) );
INVx2_ASAP7_75t_SL g133 ( .A(n_89), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_35), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_37), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_98), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_78), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_25), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_100), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_68), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_80), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_24), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_101), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_105), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_7), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_28), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_61), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_93), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_49), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_54), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_130), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_109), .B(n_0), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_126), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_125), .B(n_1), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_129), .B(n_1), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_129), .B(n_2), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_133), .B(n_4), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_125), .B(n_5), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_110), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_109), .B(n_6), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_152), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_115), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_110), .B(n_38), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_115), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
BUFx12f_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_165), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_156), .A2(n_135), .B1(n_123), .B2(n_111), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_160), .A2(n_126), .B1(n_144), .B2(n_112), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_160), .A2(n_134), .B1(n_127), .B2(n_147), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_160), .A2(n_148), .B1(n_118), .B2(n_138), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_159), .B(n_111), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_160), .A2(n_142), .B1(n_122), .B2(n_124), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_161), .A2(n_142), .B1(n_122), .B2(n_124), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_176), .B(n_138), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
OA22x2_ASAP7_75t_L g192 ( .A1(n_159), .A2(n_113), .B1(n_132), .B2(n_153), .Y(n_192) );
OAI22xp33_ASAP7_75t_SL g193 ( .A1(n_157), .A2(n_113), .B1(n_132), .B2(n_153), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_141), .B1(n_110), .B2(n_128), .Y(n_195) );
OAI22xp33_ASAP7_75t_SL g196 ( .A1(n_157), .A2(n_119), .B1(n_128), .B2(n_143), .Y(n_196) );
AO22x2_ASAP7_75t_L g197 ( .A1(n_161), .A2(n_145), .B1(n_143), .B2(n_119), .Y(n_197) );
AO22x2_ASAP7_75t_L g198 ( .A1(n_161), .A2(n_145), .B1(n_152), .B2(n_140), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_176), .A2(n_110), .B1(n_140), .B2(n_149), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_176), .B(n_110), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_151), .B1(n_150), .B2(n_139), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_163), .A2(n_137), .B1(n_136), .B2(n_121), .Y(n_204) );
OAI22xp33_ASAP7_75t_SL g205 ( .A1(n_156), .A2(n_120), .B1(n_117), .B2(n_116), .Y(n_205) );
XOR2xp5_ASAP7_75t_L g206 ( .A(n_159), .B(n_7), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_163), .A2(n_114), .B1(n_9), .B2(n_10), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_163), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_159), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_212) );
OAI22xp33_ASAP7_75t_SL g213 ( .A1(n_169), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_175), .B(n_14), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_167), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
OAI22xp5_ASAP7_75t_SL g217 ( .A1(n_169), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_175), .B(n_15), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_164), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_169), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_175), .B(n_173), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_173), .A2(n_19), .B1(n_22), .B2(n_23), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_164), .B(n_39), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_186), .B(n_164), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_179), .A2(n_173), .B(n_172), .Y(n_229) );
BUFx6f_ASAP7_75t_SL g230 ( .A(n_227), .Y(n_230) );
XNOR2x2_ASAP7_75t_L g231 ( .A(n_198), .B(n_162), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_223), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_197), .B(n_164), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_200), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_194), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_191), .Y(n_237) );
XOR2xp5_ASAP7_75t_L g238 ( .A(n_206), .B(n_197), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_181), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_190), .B(n_177), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_186), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_204), .B(n_177), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
XNOR2xp5_ASAP7_75t_L g244 ( .A(n_180), .B(n_173), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_186), .B(n_162), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_197), .B(n_154), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_224), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_225), .A2(n_172), .B(n_166), .Y(n_250) );
XOR2xp5_ASAP7_75t_L g251 ( .A(n_198), .B(n_22), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
INVxp67_ASAP7_75t_SL g253 ( .A(n_218), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_192), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_187), .B(n_162), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_205), .B(n_177), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_202), .B(n_177), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_192), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_189), .B(n_154), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_227), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_185), .B(n_154), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_219), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_207), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_183), .B(n_195), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_227), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_227), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_202), .B(n_177), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_199), .Y(n_272) );
NAND2xp33_ASAP7_75t_R g273 ( .A(n_180), .B(n_23), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_178), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_178), .A2(n_172), .B(n_166), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_217), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_182), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_182), .B(n_166), .Y(n_278) );
XOR2xp5_ASAP7_75t_L g279 ( .A(n_196), .B(n_24), .Y(n_279) );
OR2x6_ASAP7_75t_L g280 ( .A(n_226), .B(n_166), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_184), .B(n_154), .Y(n_281) );
OR2x6_ASAP7_75t_L g282 ( .A(n_226), .B(n_166), .Y(n_282) );
XOR2xp5_ASAP7_75t_L g283 ( .A(n_193), .B(n_26), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_213), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_184), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_188), .B(n_154), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_188), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_201), .Y(n_288) );
XOR2xp5_ASAP7_75t_L g289 ( .A(n_221), .B(n_26), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_201), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_203), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_203), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_244), .B(n_168), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_267), .B(n_208), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_261), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_238), .B(n_154), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_247), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_241), .Y(n_301) );
BUFx4_ASAP7_75t_SL g302 ( .A(n_280), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_287), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_247), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_241), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_244), .B(n_168), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_287), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_264), .A2(n_220), .B(n_215), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_233), .B(n_154), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_233), .B(n_168), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_228), .Y(n_312) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_248), .B(n_172), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_228), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_249), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_249), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_248), .B(n_172), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_253), .B(n_154), .Y(n_318) );
OR2x2_ASAP7_75t_SL g319 ( .A(n_254), .B(n_155), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_228), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_278), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_245), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_251), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_260), .B(n_158), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_263), .B(n_208), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_288), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_230), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_251), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_260), .B(n_158), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_245), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_235), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_264), .A2(n_220), .B(n_215), .Y(n_332) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_231), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_262), .B(n_158), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_278), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
AND2x2_ASAP7_75t_SL g337 ( .A(n_290), .B(n_158), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_240), .B(n_168), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_262), .B(n_168), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_265), .B(n_158), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_284), .B(n_158), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_269), .A2(n_270), .B(n_229), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_250), .A2(n_211), .B(n_158), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_278), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_236), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_280), .B(n_158), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_266), .B(n_168), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_245), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_346), .B(n_237), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_299), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_297), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_297), .Y(n_353) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_327), .B(n_280), .Y(n_354) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_327), .B(n_230), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_301), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_300), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_346), .B(n_243), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_300), .B(n_268), .Y(n_360) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_313), .B(n_231), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_299), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_346), .B(n_246), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_300), .B(n_268), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_305), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_312), .B(n_320), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_312), .Y(n_368) );
AND2x6_ASAP7_75t_L g369 ( .A(n_346), .B(n_230), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_301), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_297), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_312), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_327), .B(n_255), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_302), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_305), .B(n_252), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_323), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_305), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_299), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_303), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_315), .B(n_252), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_315), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_346), .B(n_232), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_369), .Y(n_383) );
BUFx5_ASAP7_75t_L g384 ( .A(n_382), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_369), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_369), .Y(n_386) );
BUFx12f_ASAP7_75t_L g387 ( .A(n_374), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_349), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_349), .B(n_346), .Y(n_391) );
INVx4_ASAP7_75t_L g392 ( .A(n_369), .Y(n_392) );
INVx3_ASAP7_75t_L g393 ( .A(n_351), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_357), .B(n_315), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_358), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_358), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_369), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_357), .B(n_316), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
INVx5_ASAP7_75t_L g403 ( .A(n_369), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
INVx3_ASAP7_75t_SL g405 ( .A(n_374), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_358), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_362), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_357), .B(n_313), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_362), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_362), .Y(n_411) );
BUFx12f_ASAP7_75t_L g412 ( .A(n_369), .Y(n_412) );
INVx4_ASAP7_75t_L g413 ( .A(n_403), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_238), .B1(n_323), .B2(n_328), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_389), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_384), .A2(n_323), .B1(n_328), .B2(n_361), .Y(n_416) );
BUFx12f_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
BUFx8_ASAP7_75t_SL g418 ( .A(n_387), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_409), .A2(n_273), .B1(n_289), .B2(n_361), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_389), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_405), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_389), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_389), .Y(n_423) );
CKINVDCx11_ASAP7_75t_R g424 ( .A(n_387), .Y(n_424) );
CKINVDCx10_ASAP7_75t_R g425 ( .A(n_387), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_402), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_396), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
INVx2_ASAP7_75t_SL g430 ( .A(n_384), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_384), .A2(n_361), .B1(n_289), .B2(n_276), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_390), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
INVx6_ASAP7_75t_L g434 ( .A(n_384), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_384), .A2(n_361), .B1(n_276), .B2(n_280), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_384), .A2(n_282), .B1(n_376), .B2(n_354), .Y(n_437) );
BUFx2_ASAP7_75t_SL g438 ( .A(n_403), .Y(n_438) );
INVx4_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_384), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_384), .A2(n_282), .B1(n_376), .B2(n_354), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_384), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_390), .Y(n_443) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_392), .A2(n_298), .B1(n_282), .B2(n_302), .Y(n_444) );
BUFx4f_ASAP7_75t_SL g445 ( .A(n_387), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_412), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_405), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g448 ( .A(n_403), .B(n_356), .Y(n_448) );
AOI21xp5_ASAP7_75t_SL g449 ( .A1(n_392), .A2(n_302), .B(n_333), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g450 ( .A(n_403), .B(n_356), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
BUFx2_ASAP7_75t_SL g452 ( .A(n_403), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
CKINVDCx11_ASAP7_75t_R g454 ( .A(n_405), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_412), .A2(n_337), .B1(n_333), .B2(n_313), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_394), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_402), .Y(n_458) );
CKINVDCx6p67_ASAP7_75t_R g459 ( .A(n_425), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
BUFx5_ASAP7_75t_L g461 ( .A(n_427), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_419), .A2(n_283), .B(n_279), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_433), .B(n_402), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_430), .B(n_409), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_444), .A2(n_384), .B1(n_282), .B2(n_412), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_424), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_419), .A2(n_403), .B1(n_392), .B2(n_386), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_414), .B(n_283), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_430), .B(n_409), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_435), .A2(n_384), .B1(n_412), .B2(n_346), .Y(n_470) );
BUFx4f_ASAP7_75t_SL g471 ( .A(n_417), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_456), .A2(n_384), .B1(n_412), .B2(n_404), .Y(n_472) );
NOR2x1p5_ASAP7_75t_L g473 ( .A(n_413), .B(n_383), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_454), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_429), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_434), .A2(n_384), .B1(n_386), .B2(n_404), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_446), .A2(n_383), .B1(n_386), .B2(n_404), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_434), .A2(n_384), .B1(n_386), .B2(n_404), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_431), .B(n_239), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_434), .A2(n_384), .B1(n_386), .B2(n_404), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_434), .B(n_239), .Y(n_482) );
OAI21xp5_ASAP7_75t_SL g483 ( .A1(n_437), .A2(n_279), .B(n_298), .Y(n_483) );
BUFx8_ASAP7_75t_SL g484 ( .A(n_418), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_425), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_429), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_440), .A2(n_384), .B1(n_386), .B2(n_404), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_433), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_420), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_420), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_440), .A2(n_384), .B1(n_383), .B2(n_409), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_442), .A2(n_383), .B1(n_385), .B2(n_400), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_446), .A2(n_383), .B1(n_400), .B2(n_385), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_433), .B(n_436), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_441), .A2(n_385), .B1(n_400), .B2(n_392), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_416), .A2(n_400), .B1(n_385), .B2(n_417), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_438), .A2(n_400), .B1(n_385), .B2(n_392), .Y(n_497) );
BUFx12f_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_458), .B(n_394), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_445), .A2(n_392), .B1(n_337), .B2(n_298), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_432), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_432), .B(n_394), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_438), .A2(n_392), .B1(n_337), .B2(n_298), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_452), .A2(n_392), .B1(n_403), .B2(n_333), .Y(n_504) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_448), .A2(n_307), .B(n_294), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_436), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_452), .A2(n_337), .B1(n_382), .B2(n_391), .Y(n_507) );
OAI222xp33_ASAP7_75t_L g508 ( .A1(n_458), .A2(n_388), .B1(n_406), .B2(n_401), .C1(n_397), .C2(n_403), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_413), .A2(n_337), .B1(n_382), .B2(n_391), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_436), .B(n_406), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_455), .Y(n_512) );
BUFx12f_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_443), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g515 ( .A1(n_443), .A2(n_256), .B1(n_307), .B2(n_294), .C1(n_364), .C2(n_360), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_449), .A2(n_257), .B(n_258), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_453), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_413), .A2(n_382), .B1(n_391), .B2(n_363), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_453), .A2(n_313), .B1(n_364), .B2(n_360), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_413), .A2(n_382), .B1(n_391), .B2(n_350), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_421), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_439), .A2(n_382), .B1(n_391), .B2(n_350), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_449), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_415), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g525 ( .A1(n_457), .A2(n_256), .B1(n_307), .B2(n_294), .C1(n_340), .C2(n_341), .Y(n_525) );
AOI222xp33_ASAP7_75t_L g526 ( .A1(n_457), .A2(n_256), .B1(n_340), .B2(n_341), .C1(n_347), .C2(n_334), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g527 ( .A1(n_439), .A2(n_405), .B1(n_403), .B2(n_313), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_455), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_426), .Y(n_529) );
AOI211xp5_ASAP7_75t_L g530 ( .A1(n_422), .A2(n_405), .B(n_340), .C(n_341), .Y(n_530) );
OAI21xp5_ASAP7_75t_SL g531 ( .A1(n_448), .A2(n_334), .B(n_373), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_439), .A2(n_391), .B1(n_350), .B2(n_359), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_439), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_465), .A2(n_423), .B1(n_388), .B2(n_399), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_462), .A2(n_391), .B1(n_403), .B2(n_359), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_523), .A2(n_451), .B1(n_426), .B2(n_403), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_474), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_467), .A2(n_391), .B1(n_403), .B2(n_359), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_488), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_527), .A2(n_350), .B1(n_359), .B2(n_363), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_527), .A2(n_350), .B1(n_359), .B2(n_363), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_519), .A2(n_388), .B1(n_399), .B2(n_410), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_468), .A2(n_350), .B1(n_359), .B2(n_363), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_476), .B(n_428), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_515), .A2(n_363), .B1(n_451), .B2(n_426), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_530), .A2(n_451), .B1(n_426), .B2(n_450), .Y(n_546) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_523), .A2(n_405), .B1(n_450), .B2(n_426), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_480), .A2(n_363), .B1(n_451), .B2(n_367), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_525), .A2(n_451), .B1(n_367), .B2(n_365), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_470), .A2(n_451), .B1(n_367), .B2(n_365), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_476), .B(n_406), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_503), .A2(n_381), .B1(n_377), .B2(n_365), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_513), .A2(n_450), .B1(n_388), .B2(n_406), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_513), .A2(n_388), .B1(n_408), .B2(n_393), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_486), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_500), .A2(n_377), .B1(n_381), .B2(n_369), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_519), .A2(n_411), .B1(n_410), .B2(n_399), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_483), .A2(n_401), .B1(n_397), .B2(n_408), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_533), .A2(n_408), .B1(n_393), .B2(n_395), .Y(n_559) );
OAI211xp5_ASAP7_75t_L g560 ( .A1(n_531), .A2(n_259), .B(n_340), .C(n_341), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_516), .A2(n_380), .B1(n_375), .B2(n_295), .C(n_339), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_526), .A2(n_381), .B1(n_377), .B2(n_369), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_533), .A2(n_397), .B1(n_401), .B2(n_411), .Y(n_563) );
OAI222xp33_ASAP7_75t_L g564 ( .A1(n_478), .A2(n_411), .B1(n_410), .B2(n_396), .C1(n_407), .C2(n_398), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_486), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_521), .B(n_27), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_475), .A2(n_369), .B1(n_174), .B2(n_373), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_475), .A2(n_174), .B1(n_373), .B2(n_317), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_501), .B(n_398), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_482), .A2(n_347), .B1(n_334), .B2(n_295), .C(n_325), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_471), .A2(n_408), .B1(n_395), .B2(n_393), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_496), .A2(n_347), .B(n_375), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_475), .A2(n_174), .B1(n_373), .B2(n_317), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_501), .B(n_398), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_514), .B(n_398), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_507), .A2(n_398), .B1(n_407), .B2(n_408), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_463), .B(n_407), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_495), .A2(n_174), .B1(n_373), .B2(n_317), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_509), .A2(n_174), .B1(n_317), .B2(n_395), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_459), .A2(n_380), .B1(n_347), .B2(n_334), .C(n_339), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_514), .B(n_407), .Y(n_581) );
AOI222xp33_ASAP7_75t_L g582 ( .A1(n_466), .A2(n_317), .B1(n_324), .B2(n_329), .C1(n_310), .C2(n_318), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_472), .A2(n_174), .B1(n_317), .B2(n_408), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_461), .A2(n_408), .B1(n_395), .B2(n_393), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_473), .A2(n_174), .B1(n_317), .B2(n_393), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_473), .A2(n_174), .B1(n_395), .B2(n_393), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_491), .A2(n_174), .B1(n_395), .B2(n_393), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_493), .A2(n_407), .B1(n_319), .B2(n_378), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_532), .A2(n_174), .B1(n_372), .B2(n_368), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_488), .Y(n_590) );
BUFx8_ASAP7_75t_SL g591 ( .A(n_484), .Y(n_591) );
OAI222xp33_ASAP7_75t_L g592 ( .A1(n_497), .A2(n_379), .B1(n_378), .B2(n_310), .C1(n_339), .C2(n_311), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_518), .A2(n_174), .B1(n_372), .B2(n_368), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_520), .A2(n_174), .B1(n_372), .B2(n_368), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_461), .A2(n_355), .B1(n_310), .B2(n_318), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_522), .A2(n_174), .B1(n_372), .B2(n_316), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_459), .A2(n_174), .B1(n_316), .B2(n_329), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_477), .A2(n_324), .B1(n_329), .B2(n_379), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_517), .B(n_378), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_479), .A2(n_324), .B1(n_329), .B2(n_379), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_510), .B(n_379), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_481), .A2(n_324), .B1(n_370), .B2(n_356), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_487), .A2(n_370), .B1(n_356), .B2(n_310), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_464), .A2(n_370), .B1(n_356), .B2(n_338), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_469), .A2(n_370), .B1(n_338), .B2(n_366), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_508), .A2(n_325), .B(n_311), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_461), .A2(n_485), .B1(n_489), .B2(n_490), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_463), .B(n_155), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_461), .A2(n_370), .B1(n_338), .B2(n_366), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_505), .A2(n_345), .B1(n_331), .B2(n_355), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_461), .A2(n_345), .B1(n_331), .B2(n_171), .Y(n_611) );
NAND3xp33_ASAP7_75t_SL g612 ( .A(n_485), .B(n_242), .C(n_318), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_461), .A2(n_331), .B1(n_345), .B2(n_318), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_504), .A2(n_319), .B1(n_311), .B2(n_330), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_510), .B(n_27), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_461), .A2(n_155), .B1(n_170), .B2(n_171), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_499), .B(n_28), .Y(n_617) );
AOI221xp5_ASAP7_75t_SL g618 ( .A1(n_502), .A2(n_155), .B1(n_170), .B2(n_171), .C(n_319), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_461), .A2(n_155), .B1(n_170), .B2(n_171), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_498), .A2(n_327), .B1(n_353), .B2(n_352), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_492), .A2(n_498), .B1(n_524), .B2(n_499), .Y(n_621) );
OAI222xp33_ASAP7_75t_L g622 ( .A1(n_528), .A2(n_168), .B1(n_327), .B2(n_271), .C1(n_314), .C2(n_234), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_528), .A2(n_319), .B1(n_330), .B2(n_348), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_494), .A2(n_155), .B1(n_171), .B2(n_170), .C(n_167), .Y(n_624) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_529), .A2(n_327), .B1(n_353), .B2(n_352), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_506), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_506), .A2(n_348), .B1(n_322), .B2(n_314), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_529), .A2(n_155), .B1(n_171), .B2(n_170), .Y(n_628) );
OAI22xp5_ASAP7_75t_SL g629 ( .A1(n_511), .A2(n_327), .B1(n_348), .B2(n_322), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_511), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_529), .A2(n_155), .B1(n_170), .B2(n_171), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_512), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_494), .B(n_29), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_608), .B(n_537), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_547), .B(n_512), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_608), .B(n_460), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_537), .B(n_555), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_607), .B(n_460), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_566), .A2(n_155), .B(n_170), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_577), .B(n_460), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_555), .B(n_460), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_577), .B(n_460), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_540), .A2(n_308), .B1(n_326), .B2(n_303), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_612), .A2(n_155), .B1(n_171), .B2(n_170), .Y(n_644) );
OA21x2_ASAP7_75t_L g645 ( .A1(n_564), .A2(n_275), .B(n_342), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_610), .A2(n_168), .B(n_167), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_565), .B(n_155), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_626), .B(n_155), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_580), .A2(n_170), .B1(n_171), .B2(n_167), .C(n_168), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_563), .B(n_170), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_621), .B(n_170), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_617), .B(n_170), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_551), .B(n_171), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_572), .A2(n_171), .B1(n_167), .B2(n_168), .C(n_321), .Y(n_654) );
OA211x2_ASAP7_75t_L g655 ( .A1(n_541), .A2(n_29), .B(n_30), .C(n_31), .Y(n_655) );
OA211x2_ASAP7_75t_L g656 ( .A1(n_545), .A2(n_30), .B(n_32), .C(n_33), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_630), .B(n_632), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_630), .B(n_171), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_601), .B(n_32), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_633), .B(n_33), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_632), .B(n_34), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_582), .A2(n_335), .B1(n_344), .B2(n_321), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_546), .B(n_34), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_539), .B(n_36), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_535), .A2(n_312), .B(n_320), .C(n_343), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_615), .B(n_36), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_584), .B(n_168), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_539), .B(n_37), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_549), .A2(n_308), .B1(n_326), .B2(n_303), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_590), .B(n_167), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_590), .B(n_167), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_597), .A2(n_168), .B1(n_286), .B2(n_343), .C(n_272), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_588), .A2(n_168), .B1(n_353), .B2(n_352), .Y(n_673) );
AOI221x1_ASAP7_75t_SL g674 ( .A1(n_542), .A2(n_336), .B1(n_326), .B2(n_308), .C(n_304), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_542), .A2(n_321), .B1(n_344), .B2(n_335), .C(n_343), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g676 ( .A1(n_610), .A2(n_342), .B(n_332), .Y(n_676) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_568), .B(n_281), .C(n_342), .D(n_344), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_536), .B(n_352), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_624), .B(n_309), .C(n_332), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_544), .B(n_303), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_569), .B(n_304), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_574), .B(n_304), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_573), .B(n_309), .C(n_332), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_595), .B(n_309), .C(n_304), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_575), .B(n_304), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_553), .B(n_308), .C(n_326), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_581), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_559), .B(n_554), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_562), .A2(n_336), .B1(n_321), .B2(n_335), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_567), .B(n_336), .C(n_353), .Y(n_690) );
AND2x2_ASAP7_75t_SL g691 ( .A(n_613), .B(n_352), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_534), .B(n_43), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_548), .A2(n_336), .B1(n_321), .B2(n_335), .Y(n_693) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_583), .A2(n_281), .B(n_335), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_599), .B(n_321), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_586), .B(n_371), .C(n_353), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_613), .B(n_335), .Y(n_697) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_543), .A2(n_344), .B1(n_322), .B2(n_320), .C(n_312), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_534), .B(n_344), .Y(n_699) );
AOI221xp5_ASAP7_75t_SL g700 ( .A1(n_585), .A2(n_344), .B1(n_320), .B2(n_312), .C(n_292), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_576), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_556), .A2(n_344), .B1(n_353), .B2(n_352), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_557), .B(n_44), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_571), .B(n_371), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_557), .B(n_45), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_609), .B(n_46), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_561), .A2(n_322), .B1(n_312), .B2(n_320), .C(n_306), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_576), .B(n_47), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_552), .B(n_48), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_605), .B(n_50), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_538), .A2(n_371), .B1(n_353), .B2(n_352), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_550), .B(n_51), .Y(n_712) );
OA21x2_ASAP7_75t_L g713 ( .A1(n_618), .A2(n_292), .B(n_293), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_596), .A2(n_320), .B1(n_306), .B2(n_285), .C(n_301), .Y(n_714) );
NAND4xp25_ASAP7_75t_L g715 ( .A(n_579), .B(n_320), .C(n_291), .D(n_301), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_588), .B(n_52), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_627), .B(n_53), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_627), .B(n_55), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_604), .B(n_56), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_606), .B(n_59), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_570), .B(n_60), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_620), .A2(n_371), .B1(n_353), .B2(n_352), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_560), .B(n_62), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_606), .B(n_63), .Y(n_724) );
OAI21xp33_ASAP7_75t_L g725 ( .A1(n_589), .A2(n_285), .B(n_301), .Y(n_725) );
OAI21xp5_ASAP7_75t_SL g726 ( .A1(n_592), .A2(n_306), .B(n_371), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_629), .B(n_64), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_578), .A2(n_296), .B1(n_291), .B2(n_371), .C(n_277), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_611), .B(n_66), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_618), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_587), .B(n_371), .C(n_296), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_602), .B(n_67), .Y(n_732) );
AOI21xp5_ASAP7_75t_SL g733 ( .A1(n_614), .A2(n_371), .B(n_297), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_582), .B(n_69), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_616), .B(n_70), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_629), .A2(n_296), .B1(n_297), .B2(n_291), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_730), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_726), .B(n_631), .C(n_628), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_640), .B(n_625), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_691), .A2(n_594), .B1(n_593), .B2(n_603), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_642), .B(n_619), .Y(n_741) );
AND2x4_ASAP7_75t_L g742 ( .A(n_687), .B(n_600), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_687), .B(n_598), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_657), .B(n_623), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_662), .A2(n_591), .B1(n_622), .B2(n_296), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_691), .B(n_72), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_636), .B(n_73), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_634), .B(n_74), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_701), .B(n_75), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_730), .B(n_591), .C(n_297), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_713), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_639), .B(n_296), .C(n_77), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_688), .B(n_76), .Y(n_753) );
AND2x2_ASAP7_75t_SL g754 ( .A(n_645), .B(n_297), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_637), .B(n_79), .Y(n_755) );
NOR2x1_ASAP7_75t_L g756 ( .A(n_663), .B(n_296), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_662), .A2(n_296), .B1(n_297), .B2(n_277), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_638), .B(n_81), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_638), .B(n_297), .Y(n_759) );
NOR4xp75_ASAP7_75t_L g760 ( .A(n_678), .B(n_82), .C(n_83), .D(n_84), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_678), .B(n_297), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_635), .B(n_297), .C(n_85), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_635), .B(n_87), .C(n_88), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_641), .B(n_91), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_666), .B(n_660), .C(n_734), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_648), .B(n_92), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_647), .Y(n_767) );
AND2x6_ASAP7_75t_L g768 ( .A(n_716), .B(n_95), .Y(n_768) );
AND2x4_ASAP7_75t_L g769 ( .A(n_647), .B(n_96), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_674), .B(n_99), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_651), .B(n_102), .C(n_104), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_656), .A2(n_106), .B1(n_107), .B2(n_108), .Y(n_772) );
NOR3xp33_ASAP7_75t_SL g773 ( .A(n_667), .B(n_211), .C(n_677), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g774 ( .A(n_733), .B(n_644), .C(n_650), .Y(n_774) );
NAND4xp75_ASAP7_75t_L g775 ( .A(n_655), .B(n_667), .C(n_700), .D(n_646), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_658), .B(n_664), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_658), .B(n_668), .Y(n_777) );
AO21x2_ASAP7_75t_L g778 ( .A1(n_661), .A2(n_703), .B(n_705), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_692), .B(n_720), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_699), .B(n_659), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_720), .B(n_733), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_644), .B(n_686), .C(n_673), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_720), .B(n_645), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_676), .B(n_653), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_645), .B(n_671), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g786 ( .A(n_727), .B(n_649), .C(n_704), .D(n_724), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_670), .B(n_704), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_675), .B(n_680), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_681), .B(n_682), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_685), .Y(n_790) );
NAND3xp33_ASAP7_75t_L g791 ( .A(n_652), .B(n_727), .C(n_654), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_723), .B(n_665), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_698), .B(n_715), .C(n_725), .D(n_721), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_693), .A2(n_672), .B1(n_694), .B2(n_732), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_696), .B(n_713), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_710), .B(n_706), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g797 ( .A1(n_714), .A2(n_717), .B(n_718), .C(n_708), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_707), .A2(n_697), .B1(n_689), .B2(n_695), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_713), .Y(n_799) );
INVx3_ASAP7_75t_L g800 ( .A(n_712), .Y(n_800) );
AO21x2_ASAP7_75t_L g801 ( .A1(n_709), .A2(n_719), .B(n_690), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_722), .Y(n_802) );
AOI211xp5_ASAP7_75t_L g803 ( .A1(n_736), .A2(n_669), .B(n_711), .C(n_728), .Y(n_803) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_731), .B(n_683), .C(n_729), .Y(n_804) );
NOR3xp33_ASAP7_75t_L g805 ( .A(n_729), .B(n_679), .C(n_735), .Y(n_805) );
AO21x2_ASAP7_75t_L g806 ( .A1(n_684), .A2(n_735), .B(n_702), .Y(n_806) );
OA211x2_ASAP7_75t_L g807 ( .A1(n_643), .A2(n_638), .B(n_678), .C(n_635), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_726), .B(n_730), .C(n_638), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_726), .A2(n_558), .B1(n_688), .B2(n_656), .Y(n_809) );
AO21x2_ASAP7_75t_L g810 ( .A1(n_635), .A2(n_650), .B(n_638), .Y(n_810) );
INVxp67_ASAP7_75t_L g811 ( .A(n_730), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_634), .B(n_687), .Y(n_812) );
NAND4xp75_ASAP7_75t_L g813 ( .A(n_663), .B(n_638), .C(n_656), .D(n_688), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_662), .A2(n_558), .B1(n_612), .B2(n_462), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_809), .A2(n_813), .B1(n_765), .B2(n_805), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_812), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_737), .B(n_811), .Y(n_817) );
NAND4xp75_ASAP7_75t_L g818 ( .A(n_807), .B(n_753), .C(n_773), .D(n_756), .Y(n_818) );
INVx5_ASAP7_75t_L g819 ( .A(n_751), .Y(n_819) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_737), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_811), .B(n_790), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_744), .B(n_784), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_739), .B(n_781), .Y(n_823) );
NOR2x1_ASAP7_75t_L g824 ( .A(n_808), .B(n_750), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_799), .Y(n_825) );
XOR2x2_ASAP7_75t_L g826 ( .A(n_765), .B(n_775), .Y(n_826) );
NOR2xp33_ASAP7_75t_SL g827 ( .A(n_768), .B(n_793), .Y(n_827) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_770), .B(n_791), .C(n_763), .Y(n_828) );
XOR2xp5_ASAP7_75t_L g829 ( .A(n_776), .B(n_777), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_805), .A2(n_814), .B1(n_792), .B2(n_796), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_742), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_787), .Y(n_832) );
XNOR2xp5_ASAP7_75t_L g833 ( .A(n_779), .B(n_814), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_742), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_742), .Y(n_835) );
INVxp67_ASAP7_75t_L g836 ( .A(n_810), .Y(n_836) );
NAND4xp75_ASAP7_75t_SL g837 ( .A(n_783), .B(n_792), .C(n_758), .D(n_746), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_789), .B(n_767), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_743), .Y(n_839) );
INVx1_ASAP7_75t_SL g840 ( .A(n_769), .Y(n_840) );
XOR2x2_ASAP7_75t_L g841 ( .A(n_760), .B(n_786), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_802), .B(n_785), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_802), .B(n_800), .Y(n_843) );
AND3x1_ASAP7_75t_L g844 ( .A(n_773), .B(n_745), .C(n_800), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_741), .B(n_810), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_743), .Y(n_846) );
NAND4xp75_ASAP7_75t_SL g847 ( .A(n_796), .B(n_749), .C(n_768), .D(n_806), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_743), .Y(n_848) );
XOR2xp5_ASAP7_75t_L g849 ( .A(n_780), .B(n_740), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_774), .A2(n_759), .B1(n_745), .B2(n_761), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g851 ( .A(n_795), .B(n_754), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_797), .B(n_788), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_806), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_778), .Y(n_854) );
AND2x4_ASAP7_75t_L g855 ( .A(n_778), .B(n_801), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_755), .Y(n_856) );
NAND4xp75_ASAP7_75t_L g857 ( .A(n_794), .B(n_772), .C(n_748), .D(n_747), .Y(n_857) );
XOR2x2_ASAP7_75t_L g858 ( .A(n_826), .B(n_804), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_815), .A2(n_803), .B1(n_762), .B2(n_782), .Y(n_859) );
BUFx2_ASAP7_75t_L g860 ( .A(n_832), .Y(n_860) );
INVx1_ASAP7_75t_SL g861 ( .A(n_840), .Y(n_861) );
XOR2x2_ASAP7_75t_L g862 ( .A(n_826), .B(n_804), .Y(n_862) );
XOR2x2_ASAP7_75t_L g863 ( .A(n_833), .B(n_738), .Y(n_863) );
XNOR2x1_ASAP7_75t_L g864 ( .A(n_830), .B(n_769), .Y(n_864) );
NOR2xp33_ASAP7_75t_SL g865 ( .A(n_827), .B(n_818), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_842), .B(n_801), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g867 ( .A(n_852), .B(n_849), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_831), .Y(n_868) );
INVxp67_ASAP7_75t_L g869 ( .A(n_852), .Y(n_869) );
XNOR2xp5_ASAP7_75t_L g870 ( .A(n_841), .B(n_798), .Y(n_870) );
INVx6_ASAP7_75t_L g871 ( .A(n_819), .Y(n_871) );
XOR2xp5_ASAP7_75t_L g872 ( .A(n_837), .B(n_798), .Y(n_872) );
INVx1_ASAP7_75t_SL g873 ( .A(n_821), .Y(n_873) );
BUFx2_ASAP7_75t_L g874 ( .A(n_832), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_834), .Y(n_875) );
INVx1_ASAP7_75t_SL g876 ( .A(n_838), .Y(n_876) );
OAI22xp33_ASAP7_75t_R g877 ( .A1(n_853), .A2(n_768), .B1(n_752), .B2(n_771), .Y(n_877) );
XNOR2xp5_ASAP7_75t_L g878 ( .A(n_841), .B(n_764), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_835), .Y(n_879) );
XNOR2xp5_ASAP7_75t_L g880 ( .A(n_844), .B(n_766), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_843), .B(n_845), .Y(n_881) );
INVx5_ASAP7_75t_L g882 ( .A(n_819), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_822), .B(n_768), .Y(n_883) );
AO22x1_ASAP7_75t_L g884 ( .A1(n_824), .A2(n_768), .B1(n_752), .B2(n_757), .Y(n_884) );
XNOR2xp5_ASAP7_75t_L g885 ( .A(n_858), .B(n_857), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_868), .Y(n_886) );
OA22x2_ASAP7_75t_L g887 ( .A1(n_870), .A2(n_820), .B1(n_817), .B2(n_855), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_875), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_879), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_860), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_858), .A2(n_828), .B1(n_850), .B2(n_823), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_864), .A2(n_851), .B1(n_820), .B2(n_829), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_876), .Y(n_893) );
INVxp67_ASAP7_75t_L g894 ( .A(n_867), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_874), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_882), .Y(n_896) );
XOR2x2_ASAP7_75t_SL g897 ( .A(n_859), .B(n_847), .Y(n_897) );
INVx1_ASAP7_75t_SL g898 ( .A(n_861), .Y(n_898) );
OA22x2_ASAP7_75t_L g899 ( .A1(n_869), .A2(n_855), .B1(n_836), .B2(n_851), .Y(n_899) );
OA22x2_ASAP7_75t_L g900 ( .A1(n_872), .A2(n_855), .B1(n_836), .B2(n_839), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_893), .Y(n_901) );
OAI322xp33_ASAP7_75t_L g902 ( .A1(n_887), .A2(n_867), .A3(n_865), .B1(n_864), .B2(n_873), .C1(n_862), .C2(n_878), .Y(n_902) );
AOI322xp5_ASAP7_75t_L g903 ( .A1(n_894), .A2(n_883), .A3(n_881), .B1(n_862), .B2(n_866), .C1(n_863), .C2(n_846), .Y(n_903) );
INVx2_ASAP7_75t_L g904 ( .A(n_898), .Y(n_904) );
INVx2_ASAP7_75t_SL g905 ( .A(n_890), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_898), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_895), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_886), .Y(n_908) );
OAI322xp33_ASAP7_75t_L g909 ( .A1(n_887), .A2(n_880), .A3(n_883), .B1(n_863), .B2(n_866), .C1(n_854), .C2(n_848), .Y(n_909) );
NOR4xp25_ASAP7_75t_L g910 ( .A(n_902), .B(n_894), .C(n_892), .D(n_897), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_906), .A2(n_892), .B1(n_885), .B2(n_891), .Y(n_911) );
INVx1_ASAP7_75t_SL g912 ( .A(n_904), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_904), .Y(n_913) );
NAND2x1_ASAP7_75t_SL g914 ( .A(n_901), .B(n_896), .Y(n_914) );
OAI22xp33_ASAP7_75t_L g915 ( .A1(n_911), .A2(n_900), .B1(n_899), .B2(n_905), .Y(n_915) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_912), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_913), .A2(n_900), .B1(n_905), .B2(n_907), .Y(n_917) );
NAND2xp5_ASAP7_75t_SL g918 ( .A(n_915), .B(n_910), .Y(n_918) );
AO22x2_ASAP7_75t_L g919 ( .A1(n_917), .A2(n_901), .B1(n_907), .B2(n_908), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_916), .B(n_903), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_919), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_919), .Y(n_922) );
OR2x2_ASAP7_75t_L g923 ( .A(n_921), .B(n_918), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_922), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_924), .Y(n_925) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_923), .A2(n_920), .B1(n_899), .B2(n_909), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_925), .A2(n_871), .B1(n_914), .B2(n_882), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_927), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_928), .A2(n_926), .B1(n_877), .B2(n_828), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_929), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_930), .A2(n_888), .B1(n_889), .B2(n_914), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_931), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_932), .A2(n_884), .B1(n_881), .B2(n_854), .C(n_882), .Y(n_933) );
AOI211xp5_ASAP7_75t_L g934 ( .A1(n_933), .A2(n_816), .B(n_856), .C(n_825), .Y(n_934) );
endmodule