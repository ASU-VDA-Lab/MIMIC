module fake_jpeg_30524_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_16),
.Y(n_61)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_5),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_29),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_30),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_50),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_55),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_64),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_21),
.B1(n_18),
.B2(n_24),
.Y(n_58)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_24),
.B1(n_26),
.B2(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_23),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_66),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_78),
.Y(n_100)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_20),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_34),
.A3(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_51),
.B(n_1),
.C(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_5),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_10),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_11),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_89),
.A2(n_59),
.B1(n_50),
.B2(n_58),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_53),
.C(n_56),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_102),
.C(n_103),
.Y(n_121)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_68),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_51),
.B(n_1),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_91),
.B(n_106),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_51),
.B1(n_1),
.B2(n_0),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_71),
.B1(n_86),
.B2(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_13),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_92),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_85),
.B1(n_89),
.B2(n_69),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_76),
.B1(n_69),
.B2(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_51),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_124),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_104),
.C(n_90),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_93),
.B(n_104),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_133),
.C(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_110),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_142),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_128),
.C(n_122),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_145),
.B(n_138),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_151),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_140),
.B(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_112),
.C(n_133),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.C(n_157),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_158),
.B(n_152),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_115),
.B(n_124),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_131),
.B(n_117),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_131),
.B1(n_117),
.B2(n_147),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_161),
.Y(n_164)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_110),
.B1(n_118),
.B2(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_162),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_167),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_164),
.Y(n_170)
);


endmodule