module fake_jpeg_10319_n_229 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_25),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_22),
.B1(n_33),
.B2(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_30),
.B1(n_28),
.B2(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_73),
.B1(n_26),
.B2(n_28),
.Y(n_79)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_70),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_24),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_9),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_75),
.B(n_66),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_53),
.B1(n_16),
.B2(n_15),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_35),
.B1(n_20),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_89),
.B1(n_74),
.B2(n_103),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_34),
.B1(n_17),
.B2(n_19),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_90),
.B1(n_66),
.B2(n_80),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_2),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_97),
.B(n_103),
.C(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_96),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_30),
.B1(n_17),
.B2(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_17),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_104),
.B1(n_56),
.B2(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_12),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_81),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_13),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_10),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_117),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_106),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_49),
.B1(n_53),
.B2(n_62),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_112),
.B1(n_119),
.B2(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_116),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_16),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_92),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_90),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_85),
.C(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_88),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_139),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_120),
.B1(n_127),
.B2(n_109),
.C(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_149),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_99),
.C(n_98),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_144),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_85),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_112),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_82),
.B(n_124),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_84),
.C(n_85),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_113),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_148),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_164),
.B(n_147),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_166),
.B(n_130),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_123),
.B1(n_119),
.B2(n_122),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_169),
.B1(n_170),
.B2(n_142),
.Y(n_184)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_161),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_168),
.B1(n_149),
.B2(n_131),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_133),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_165),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_82),
.B(n_128),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_151),
.B1(n_139),
.B2(n_134),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_128),
.B1(n_86),
.B2(n_84),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_86),
.B1(n_115),
.B2(n_116),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_176),
.B(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_141),
.C(n_136),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_159),
.C(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_116),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_164),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_182),
.B(n_162),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_143),
.B1(n_145),
.B2(n_115),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_168),
.B1(n_155),
.B2(n_153),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_170),
.B1(n_169),
.B2(n_142),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_150),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_175),
.B1(n_179),
.B2(n_172),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_152),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_182),
.Y(n_207)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_193),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_171),
.C(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_178),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_189),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_185),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_203),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_174),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_207),
.C(n_192),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_191),
.B1(n_176),
.B2(n_193),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g208 ( 
.A(n_199),
.B(n_195),
.C(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_204),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_187),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_188),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_201),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_218),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_197),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_211),
.B(n_213),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_210),
.C(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_225),
.B1(n_222),
.B2(n_220),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_227),
.B(n_143),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_184),
.B1(n_208),
.B2(n_156),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_161),
.Y(n_229)
);


endmodule