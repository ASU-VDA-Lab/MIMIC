module real_jpeg_33737_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_0),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_0),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_1),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_3),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_4),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_4),
.Y(n_199)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_4),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_5),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_5),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_183),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g410 ( 
.A1(n_5),
.A2(n_183),
.B1(n_411),
.B2(n_414),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_5),
.A2(n_183),
.B1(n_454),
.B2(n_457),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_8),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

AO22x2_ASAP7_75t_L g135 ( 
.A1(n_8),
.A2(n_25),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_8),
.A2(n_25),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_25),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_56),
.B1(n_102),
.B2(n_105),
.Y(n_101)
);

AOI22x1_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_56),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g233 ( 
.A1(n_10),
.A2(n_56),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g431 ( 
.A(n_10),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_10),
.B(n_111),
.Y(n_449)
);

OAI32xp33_ASAP7_75t_L g468 ( 
.A1(n_10),
.A2(n_200),
.A3(n_469),
.B1(n_473),
.B2(n_480),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_11),
.B(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_12),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_13),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_13),
.A2(n_67),
.B1(n_196),
.B2(n_200),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_13),
.A2(n_67),
.B1(n_220),
.B2(n_224),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_13),
.A2(n_67),
.B1(n_311),
.B2(n_315),
.Y(n_310)
);

OAI31xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_165),
.A3(n_538),
.B(n_541),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

OAI31xp33_ASAP7_75t_L g545 ( 
.A1(n_16),
.A2(n_537),
.A3(n_538),
.B(n_543),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_164),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_58),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_18),
.B(n_58),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_20),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_21),
.B(n_50),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_23),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_24),
.Y(n_182)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_56),
.Y(n_57)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_28),
.Y(n_252)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_31),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_31),
.B(n_178),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_SL g325 ( 
.A1(n_31),
.A2(n_52),
.B(n_61),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_31),
.B(n_52),
.Y(n_351)
);

NOR2x1p5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_41),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_35),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_41),
.B(n_178),
.Y(n_177)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_42),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_43),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_44),
.Y(n_146)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_45),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_46),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_46),
.Y(n_427)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_49),
.B(n_247),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_49),
.B(n_247),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_51),
.B(n_56),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_56),
.B(n_57),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI32xp33_ASAP7_75t_L g423 ( 
.A1(n_56),
.A2(n_424),
.A3(n_428),
.B1(n_430),
.B2(n_431),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_56),
.B(n_481),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_56),
.B(n_74),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_56),
.B(n_499),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_57),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_156),
.C(n_160),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_59),
.B(n_532),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.C(n_108),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_60),
.B(n_363),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B(n_70),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_63),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_71),
.B(n_352),
.C(n_360),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_72),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_72),
.A2(n_109),
.B1(n_346),
.B2(n_364),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_72),
.B(n_382),
.C(n_384),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_72),
.A2(n_346),
.B1(n_382),
.B2(n_391),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_86),
.B(n_101),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_73),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_73),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_73),
.B(n_101),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_73),
.B(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_87),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_81),
.B2(n_84),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_76),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_79),
.Y(n_497)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_80),
.Y(n_235)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_85),
.Y(n_213)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_85),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_86),
.B(n_101),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_86),
.B(n_189),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_86),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_86),
.B(n_410),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_94),
.B2(n_99),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_90),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_98),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_103),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_109),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_134),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_110),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_125),
.Y(n_110)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_111),
.B(n_135),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_111),
.Y(n_319)
);

NAND2xp33_ASAP7_75t_SL g383 ( 
.A(n_111),
.B(n_242),
.Y(n_383)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AO21x2_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_143),
.B(n_150),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_123),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_124),
.Y(n_226)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21x1_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_142),
.B(n_163),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g291 ( 
.A(n_126),
.B(n_142),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_129),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_130),
.Y(n_318)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_134),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_134),
.B(n_383),
.Y(n_382)
);

NAND2x1_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_141),
.B(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_142),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_150),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_156),
.A2(n_160),
.B1(n_161),
.B2(n_533),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_156),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_159),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_159),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_161),
.B(n_272),
.C(n_274),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_529),
.B(n_537),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI31xp33_ASAP7_75t_SL g541 ( 
.A1(n_167),
.A2(n_542),
.A3(n_544),
.B(n_545),
.Y(n_541)
);

AOI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_372),
.B(n_524),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_335),
.B(n_338),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_295),
.B(n_297),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_270),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_172),
.B(n_270),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_216),
.C(n_238),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_174),
.B(n_216),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_185),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_177),
.B(n_351),
.Y(n_384)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_194),
.Y(n_185)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_186),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_187),
.B(n_409),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_188),
.A2(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_188),
.B(n_437),
.Y(n_447)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_191),
.Y(n_413)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_192),
.Y(n_429)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g385 ( 
.A(n_194),
.B(n_386),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_202),
.B(n_206),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_195),
.A2(n_229),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_201),
.Y(n_456)
);

AO21x2_ASAP7_75t_L g282 ( 
.A1(n_202),
.A2(n_204),
.B(n_283),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g502 ( 
.A1(n_202),
.A2(n_283),
.B(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_211),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_203),
.A2(n_233),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_203),
.B(n_453),
.Y(n_452)
);

INVx4_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_206),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_206),
.B(n_452),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx2_ASAP7_75t_SL g458 ( 
.A(n_213),
.Y(n_458)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2x2_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_228),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_227),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_218),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_287)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_226),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_227),
.B(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_229),
.B(n_503),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_230),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_238),
.B(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.C(n_248),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_239),
.A2(n_240),
.B1(n_246),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_241),
.B(n_349),
.Y(n_397)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_246),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_248),
.B(n_379),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_259),
.B(n_267),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_250),
.B(n_260),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.C(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_264),
.B(n_266),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_267),
.B(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_275),
.Y(n_270)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_281),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g421 ( 
.A1(n_281),
.A2(n_282),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_282),
.A2(n_356),
.B(n_357),
.Y(n_355)
);

NOR2x1_ASAP7_75t_SL g438 ( 
.A(n_282),
.B(n_423),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_285),
.Y(n_301)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

AOI22x1_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_288)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_291),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_294),
.Y(n_333)
);

NOR4xp25_ASAP7_75t_L g518 ( 
.A(n_295),
.B(n_336),
.C(n_519),
.D(n_522),
.Y(n_518)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_303),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_303),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.C(n_302),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_330),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_304)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_305),
.B(n_331),
.C(n_368),
.Y(n_367)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_308),
.B(n_321),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_308),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_307),
.B(n_437),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_319),
.B(n_320),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_310),
.A2(n_348),
.B(n_349),
.Y(n_347)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_326),
.B2(n_327),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_325),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.C(n_334),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_366),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_358),
.Y(n_340)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_341),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_353),
.C(n_355),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_342),
.A2(n_343),
.B1(n_353),
.B2(n_354),
.Y(n_371)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_350),
.B2(n_352),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_350),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_350),
.A2(n_352),
.B1(n_362),
.B2(n_365),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_352),
.B(n_359),
.C(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_358),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_362),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_365),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_367),
.B(n_369),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_402),
.B(n_518),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_387),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_374),
.B(n_521),
.Y(n_520)
);

NAND2x1_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_375),
.B(n_377),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_385),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_401),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_385),
.Y(n_401)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_390),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_400),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_388),
.B(n_400),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.C(n_398),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_389),
.B(n_516),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_392),
.B(n_398),
.Y(n_516)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_397),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_393),
.A2(n_395),
.B1(n_396),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

AO21x1_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_513),
.B(n_517),
.Y(n_403)
);

OAI21x1_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_443),
.B(n_512),
.Y(n_404)
);

NOR2x1_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_434),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_406),
.B(n_434),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_417),
.C(n_420),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_408),
.B(n_418),
.Y(n_460)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_460),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_439),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_438),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_436),
.B(n_438),
.C(n_439),
.Y(n_514)
);

XOR2x2_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.Y(n_439)
);

AOI21x1_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_461),
.B(n_511),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_459),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_SL g511 ( 
.A(n_445),
.B(n_459),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.C(n_450),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_448),
.B1(n_449),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_500),
.Y(n_503)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_488),
.B(n_510),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_463),
.B(n_466),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_486),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_467),
.B(n_487),
.Y(n_507)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_468),
.B(n_486),
.Y(n_508)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AOI21x1_ASAP7_75t_SL g488 ( 
.A1(n_489),
.A2(n_505),
.B(n_509),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_493),
.B(n_504),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_492),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_502),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_498),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NAND3xp33_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_507),
.C(n_508),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_506),
.A2(n_507),
.B(n_508),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_515),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

BUFx2_ASAP7_75t_SL g524 ( 
.A(n_525),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_527),
.C(n_528),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_529),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_534),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_535),
.Y(n_537)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_539),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_539),
.B(n_540),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_543),
.Y(n_542)
);


endmodule