module fake_jpeg_19_n_42 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_42);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_0),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_14),
.B(n_13),
.C(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_20),
.B1(n_19),
.B2(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

AND2x6_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_2),
.Y(n_26)
);

XOR2x2_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_26),
.B(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_34),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_30),
.C(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_32),
.B1(n_34),
.B2(n_27),
.Y(n_38)
);

OAI21x1_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_35),
.B(n_7),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_39),
.A3(n_38),
.B1(n_9),
.B2(n_10),
.C1(n_8),
.C2(n_4),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_8),
.Y(n_42)
);


endmodule