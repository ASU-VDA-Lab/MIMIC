module fake_jpeg_10786_n_610 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_610);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_610;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_64),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_9),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_66),
.Y(n_170)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_68),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_70),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_73),
.Y(n_181)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_74),
.Y(n_168)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_79),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_8),
.B1(n_17),
.B2(n_2),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_80),
.A2(n_31),
.B1(n_59),
.B2(n_49),
.Y(n_182)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_82),
.Y(n_179)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g202 ( 
.A(n_84),
.Y(n_202)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_94),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_40),
.B(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_100),
.B(n_126),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_112),
.Y(n_191)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_27),
.B(n_7),
.Y(n_122)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_43),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_127),
.Y(n_148)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_43),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_40),
.B(n_7),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_31),
.B(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_34),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_50),
.B1(n_28),
.B2(n_21),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_130),
.A2(n_136),
.B1(n_137),
.B2(n_145),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_62),
.A2(n_21),
.B1(n_28),
.B2(n_52),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_135),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_68),
.A2(n_28),
.B1(n_48),
.B2(n_33),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_68),
.A2(n_33),
.B1(n_48),
.B2(n_56),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_117),
.B1(n_123),
.B2(n_48),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_151),
.B(n_157),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_34),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_185),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_61),
.C(n_60),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_192),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_73),
.A2(n_60),
.B1(n_56),
.B2(n_45),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_162),
.A2(n_182),
.B1(n_200),
.B2(n_203),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_44),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_174),
.B(n_175),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_44),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_111),
.A2(n_37),
.B1(n_59),
.B2(n_49),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_196),
.B1(n_198),
.B2(n_101),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_66),
.B(n_61),
.C(n_45),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_125),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_79),
.A2(n_58),
.B1(n_41),
.B2(n_2),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_71),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_107),
.A2(n_12),
.B1(n_18),
.B2(n_2),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_84),
.B(n_12),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_204),
.B(n_207),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_86),
.B(n_13),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_88),
.B(n_10),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_210),
.B(n_10),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_0),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_211),
.B(n_227),
.Y(n_290)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_212),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_78),
.B1(n_120),
.B2(n_90),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g317 ( 
.A1(n_213),
.A2(n_221),
.B1(n_267),
.B2(n_275),
.Y(n_317)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_145),
.B1(n_162),
.B2(n_130),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_216),
.A2(n_250),
.B1(n_265),
.B2(n_273),
.Y(n_292)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_148),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_220),
.B(n_243),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_159),
.A2(n_119),
.B1(n_105),
.B2(n_102),
.Y(n_221)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_222),
.Y(n_313)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_223),
.Y(n_299)
);

BUFx8_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

BUFx2_ASAP7_75t_SL g338 ( 
.A(n_224),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_225),
.A2(n_211),
.B1(n_266),
.B2(n_230),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_131),
.A2(n_18),
.B(n_16),
.C(n_3),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_149),
.A2(n_97),
.B(n_95),
.C(n_94),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g306 ( 
.A1(n_228),
.A2(n_229),
.B1(n_176),
.B2(n_209),
.Y(n_306)
);

AO22x1_ASAP7_75t_SL g229 ( 
.A1(n_139),
.A2(n_93),
.B1(n_91),
.B2(n_0),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_201),
.B1(n_169),
.B2(n_154),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_230),
.A2(n_225),
.B1(n_232),
.B2(n_252),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_133),
.B(n_0),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_231),
.B(n_233),
.C(n_277),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_155),
.Y(n_232)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_232),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_138),
.B(n_1),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_141),
.Y(n_234)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_236),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_168),
.B(n_3),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_238),
.B(n_252),
.Y(n_304)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_129),
.Y(n_240)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

AO22x1_ASAP7_75t_L g241 ( 
.A1(n_142),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_241),
.A2(n_246),
.B(n_255),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_208),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_242),
.B(n_263),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_183),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_244),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_146),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_246),
.B(n_262),
.Y(n_323)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_132),
.Y(n_248)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_203),
.A2(n_136),
.B1(n_137),
.B2(n_181),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_41),
.Y(n_252)
);

BUFx4f_ASAP7_75t_SL g253 ( 
.A(n_156),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_253),
.Y(n_284)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_132),
.Y(n_254)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_156),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_257),
.Y(n_326)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_259),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_134),
.B(n_4),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_260),
.B(n_270),
.Y(n_305)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_191),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_191),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_264),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_181),
.A2(n_202),
.B1(n_140),
.B2(n_179),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_206),
.B(n_10),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_215),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_159),
.A2(n_41),
.B1(n_58),
.B2(n_18),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_147),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_269),
.Y(n_328)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_271),
.A2(n_281),
.B1(n_282),
.B2(n_242),
.Y(n_311)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_161),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_274),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_140),
.A2(n_14),
.B1(n_58),
.B2(n_202),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_164),
.Y(n_274)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_188),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_153),
.A2(n_14),
.B1(n_58),
.B2(n_180),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_276),
.A2(n_279),
.B1(n_236),
.B2(n_235),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_171),
.B(n_187),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_153),
.A2(n_180),
.B1(n_197),
.B2(n_190),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_144),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_280),
.B(n_283),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_164),
.Y(n_281)
);

BUFx4f_ASAP7_75t_SL g282 ( 
.A(n_208),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_146),
.B(n_166),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_219),
.A2(n_165),
.B1(n_166),
.B2(n_209),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_285),
.A2(n_322),
.B1(n_332),
.B2(n_274),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_215),
.B(n_165),
.C(n_188),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_286),
.B(n_302),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_309),
.B1(n_314),
.B2(n_319),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_229),
.A2(n_176),
.B1(n_190),
.B2(n_197),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_295),
.A2(n_289),
.B1(n_284),
.B2(n_334),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_164),
.C(n_188),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g372 ( 
.A1(n_306),
.A2(n_307),
.B(n_317),
.C(n_286),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g307 ( 
.A1(n_216),
.A2(n_258),
.B1(n_229),
.B2(n_250),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_310),
.B(n_241),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_311),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_251),
.A2(n_215),
.B1(n_278),
.B2(n_247),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g319 ( 
.A1(n_228),
.A2(n_237),
.B1(n_271),
.B2(n_222),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_265),
.A2(n_233),
.B1(n_231),
.B2(n_277),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_320),
.A2(n_214),
.B(n_217),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_232),
.B1(n_257),
.B2(n_259),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_245),
.A2(n_254),
.B1(n_261),
.B2(n_263),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_325),
.A2(n_281),
.B1(n_218),
.B2(n_269),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_301),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_231),
.B(n_233),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_301),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_249),
.B(n_268),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_335),
.B(n_298),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_256),
.A2(n_239),
.B1(n_234),
.B2(n_212),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_336),
.B1(n_293),
.B2(n_297),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_342),
.B(n_353),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_373),
.Y(n_387)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_227),
.B(n_253),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_345),
.A2(n_371),
.B(n_374),
.Y(n_401)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_328),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_328),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_240),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_369),
.Y(n_392)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_292),
.A2(n_253),
.B1(n_282),
.B2(n_224),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_357),
.A2(n_370),
.B1(n_372),
.B2(n_383),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_290),
.A2(n_282),
.B(n_224),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_358),
.A2(n_368),
.B(n_303),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_359),
.A2(n_364),
.B(n_386),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_362),
.B(n_365),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_307),
.A2(n_292),
.B1(n_319),
.B2(n_290),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_363),
.A2(n_375),
.B1(n_378),
.B2(n_380),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_328),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_304),
.A2(n_323),
.B(n_330),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_299),
.B(n_305),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_307),
.A2(n_320),
.B1(n_310),
.B2(n_332),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_302),
.A2(n_307),
.B(n_339),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_296),
.B(n_306),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_306),
.A2(n_317),
.B1(n_299),
.B2(n_341),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_300),
.Y(n_377)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_377),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_306),
.A2(n_300),
.B1(n_293),
.B2(n_318),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_338),
.Y(n_379)
);

NAND2x1_ASAP7_75t_SL g418 ( 
.A(n_379),
.B(n_381),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_300),
.A2(n_318),
.B1(n_297),
.B2(n_340),
.Y(n_380)
);

XOR2x1_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_296),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_288),
.Y(n_391)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_294),
.Y(n_382)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_333),
.A2(n_313),
.B1(n_331),
.B2(n_316),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_313),
.B1(n_331),
.B2(n_321),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_384),
.A2(n_347),
.B1(n_344),
.B2(n_356),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_327),
.B(n_312),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_303),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_315),
.B(n_312),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_380),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_390),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_379),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_364),
.A2(n_337),
.B(n_315),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_396),
.A2(n_406),
.B(n_419),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_415),
.B1(n_342),
.B2(n_357),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_379),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_410),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_287),
.C(n_288),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_376),
.C(n_353),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_402),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_384),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_405),
.B(n_409),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_287),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_346),
.B(n_316),
.Y(n_410)
);

OA21x2_ASAP7_75t_SL g412 ( 
.A1(n_373),
.A2(n_364),
.B(n_376),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_420),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_363),
.A2(n_294),
.B1(n_346),
.B2(n_371),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_418),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_345),
.A2(n_374),
.B(n_343),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_358),
.A2(n_365),
.B(n_351),
.Y(n_420)
);

OAI32xp33_ASAP7_75t_L g425 ( 
.A1(n_395),
.A2(n_372),
.A3(n_369),
.B1(n_352),
.B2(n_362),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_430),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_426),
.A2(n_448),
.B1(n_453),
.B2(n_406),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_418),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_431),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_434),
.C(n_447),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_368),
.C(n_372),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_418),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_435),
.B(n_437),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_366),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_436),
.B(n_424),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_395),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_422),
.A2(n_375),
.B1(n_378),
.B2(n_359),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_438),
.A2(n_441),
.B1(n_450),
.B2(n_393),
.Y(n_483)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_394),
.Y(n_439)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_372),
.B1(n_359),
.B2(n_349),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_442),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_409),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_444),
.B(n_449),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_389),
.B(n_350),
.Y(n_446)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_446),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_400),
.B(n_372),
.C(n_381),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_417),
.A2(n_372),
.B1(n_361),
.B2(n_354),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_355),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_406),
.A2(n_360),
.B1(n_348),
.B2(n_386),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_398),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_451),
.Y(n_464)
);

OAI32xp33_ASAP7_75t_L g452 ( 
.A1(n_416),
.A2(n_385),
.A3(n_377),
.B1(n_367),
.B2(n_382),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_417),
.A2(n_382),
.B1(n_383),
.B2(n_415),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_387),
.B(n_396),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_402),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_391),
.C(n_420),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_392),
.Y(n_473)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_457),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_460),
.A2(n_477),
.B1(n_488),
.B2(n_433),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_401),
.B(n_388),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_468),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_463),
.B(n_440),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_392),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_465),
.B(n_475),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_449),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_467),
.B(n_446),
.Y(n_502)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_428),
.Y(n_468)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_453),
.A2(n_410),
.B1(n_416),
.B2(n_390),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_471),
.A2(n_478),
.B1(n_458),
.B2(n_433),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_SL g472 ( 
.A1(n_441),
.A2(n_401),
.B(n_388),
.C(n_419),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_472),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_476),
.C(n_455),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_425),
.B(n_399),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_432),
.B(n_454),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_448),
.A2(n_416),
.B1(n_405),
.B2(n_421),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_456),
.A2(n_393),
.B(n_399),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_485),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_483),
.A2(n_484),
.B1(n_426),
.B2(n_427),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_450),
.A2(n_393),
.B1(n_404),
.B2(n_423),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_429),
.B(n_456),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_451),
.A2(n_404),
.B1(n_423),
.B2(n_408),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_486),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_503),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_434),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_491),
.B(n_492),
.Y(n_526)
);

AOI21xp33_ASAP7_75t_L g493 ( 
.A1(n_486),
.A2(n_445),
.B(n_428),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_501),
.C(n_466),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_474),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_496),
.B(n_517),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_497),
.B(n_484),
.Y(n_528)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_478),
.Y(n_500)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_500),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_444),
.Y(n_501)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_502),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_469),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_487),
.Y(n_504)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_504),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_487),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_509),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_506),
.A2(n_510),
.B1(n_511),
.B2(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_508),
.Y(n_530)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_440),
.C(n_447),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_512),
.B(n_514),
.C(n_515),
.Y(n_527)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_489),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_463),
.B(n_429),
.C(n_458),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_424),
.C(n_457),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_459),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_516),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_461),
.B(n_431),
.Y(n_517)
);

XNOR2x1_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_483),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_519),
.B(n_528),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_492),
.B(n_479),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_529),
.B(n_533),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_534),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_481),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_496),
.B(n_472),
.C(n_477),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_512),
.B(n_481),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_537),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_472),
.C(n_488),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_536),
.B(n_539),
.C(n_494),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_472),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_507),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_538),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_515),
.B(n_472),
.C(n_464),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_517),
.B(n_452),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_540),
.B(n_506),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_536),
.A2(n_534),
.B(n_527),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_541),
.A2(n_548),
.B(n_556),
.Y(n_562)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_518),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_549),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_545),
.B(n_555),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_520),
.A2(n_500),
.B1(n_508),
.B2(n_504),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_546),
.A2(n_522),
.B1(n_540),
.B2(n_532),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_524),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_539),
.A2(n_499),
.B(n_502),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_513),
.C(n_510),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_464),
.C(n_467),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_551),
.B(n_557),
.Y(n_563)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_521),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_554),
.B(n_533),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_523),
.B(n_509),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_525),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_516),
.C(n_466),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_480),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_558),
.B(n_528),
.Y(n_566)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_559),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_560),
.B(n_561),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_529),
.C(n_530),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_519),
.C(n_537),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_565),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_566),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_558),
.B(n_480),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_567),
.B(n_570),
.C(n_572),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_495),
.C(n_459),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_551),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_571),
.A2(n_495),
.B(n_408),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_547),
.B(n_555),
.Y(n_572)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_556),
.B(n_439),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_573),
.A2(n_548),
.B(n_553),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_552),
.B(n_442),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_552),
.C(n_550),
.Y(n_582)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_575),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_564),
.A2(n_561),
.B1(n_562),
.B2(n_570),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_578),
.B(n_582),
.Y(n_591)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_579),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_563),
.A2(n_568),
.B(n_544),
.Y(n_581)
);

AOI21xp33_ASAP7_75t_L g588 ( 
.A1(n_581),
.A2(n_583),
.B(n_572),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_574),
.A2(n_544),
.B(n_550),
.Y(n_583)
);

AOI21xp33_ASAP7_75t_L g585 ( 
.A1(n_569),
.A2(n_414),
.B(n_470),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_585),
.B(n_567),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_586),
.B(n_569),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_587),
.B(n_594),
.Y(n_601)
);

OAI21xp33_ASAP7_75t_SL g596 ( 
.A1(n_588),
.A2(n_575),
.B(n_576),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_560),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_582),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_592),
.A2(n_595),
.B1(n_581),
.B2(n_583),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_584),
.B(n_413),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_414),
.Y(n_595)
);

INVxp33_ASAP7_75t_SL g602 ( 
.A(n_596),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_598),
.C(n_599),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_590),
.A2(n_578),
.B(n_577),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_589),
.Y(n_600)
);

AOI21xp33_ASAP7_75t_L g603 ( 
.A1(n_600),
.A2(n_595),
.B(n_593),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_603),
.B(n_601),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_605),
.A2(n_606),
.B1(n_604),
.B2(n_462),
.Y(n_607)
);

OAI321xp33_ASAP7_75t_L g606 ( 
.A1(n_602),
.A2(n_596),
.A3(n_591),
.B1(n_462),
.B2(n_443),
.C(n_407),
.Y(n_606)
);

BUFx24_ASAP7_75t_SL g608 ( 
.A(n_607),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_591),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_SL g610 ( 
.A1(n_609),
.A2(n_407),
.B(n_411),
.C(n_605),
.Y(n_610)
);


endmodule