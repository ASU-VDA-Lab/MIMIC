module fake_jpeg_21811_n_303 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_294;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_10),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_18),
.B(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_22),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_66),
.B1(n_32),
.B2(n_29),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_61),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_30),
.B1(n_22),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_27),
.B1(n_34),
.B2(n_28),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_58),
.B1(n_52),
.B2(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_19),
.B1(n_31),
.B2(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_2),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_12),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_57),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_36),
.A2(n_26),
.B1(n_17),
.B2(n_32),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_43),
.C(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_79),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_78),
.B(n_98),
.Y(n_125)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_80),
.Y(n_109)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_83),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_94),
.B1(n_61),
.B2(n_45),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_36),
.C(n_40),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_24),
.C(n_3),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_17),
.B(n_29),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_69),
.B(n_49),
.Y(n_107)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_102),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_12),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_11),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_49),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_124),
.B(n_101),
.Y(n_140)
);

OA22x2_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_60),
.B1(n_45),
.B2(n_46),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_97),
.A3(n_84),
.B1(n_83),
.B2(n_88),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_93),
.B1(n_76),
.B2(n_91),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_45),
.B1(n_47),
.B2(n_68),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_90),
.B1(n_96),
.B2(n_81),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_85),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_3),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_107),
.B(n_126),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_32),
.B(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_24),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_95),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_130),
.Y(n_148)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_88),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_24),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_9),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_13),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_138),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_136),
.A2(n_137),
.B(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_149),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_140),
.A2(n_111),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_133),
.B(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_146),
.B(n_150),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_98),
.B(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_152),
.B(n_164),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_160),
.B1(n_155),
.B2(n_138),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_160),
.B1(n_132),
.B2(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_71),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_163),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_161),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_77),
.B(n_75),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_124),
.B(n_108),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_97),
.B1(n_74),
.B2(n_100),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_79),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_112),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_11),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_4),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_182),
.B1(n_184),
.B2(n_191),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_158),
.B(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_136),
.C(n_140),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_186),
.C(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_131),
.B1(n_112),
.B2(n_108),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_121),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_192),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_111),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_151),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_122),
.B1(n_88),
.B2(n_72),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_3),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_181),
.B(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_196),
.B(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_207),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_212),
.B(n_218),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_187),
.A2(n_137),
.B1(n_139),
.B2(n_154),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_179),
.B1(n_177),
.B2(n_195),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_157),
.CI(n_165),
.CON(n_202),
.SN(n_202)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_202),
.B(n_204),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_114),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_214),
.C(n_178),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_122),
.B1(n_163),
.B2(n_114),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_208),
.B(n_193),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_189),
.A2(n_163),
.B1(n_5),
.B2(n_7),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_182),
.B1(n_191),
.B2(n_171),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_172),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_5),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_8),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_194),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_175),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_224),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_189),
.B(n_192),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_231),
.B(n_234),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_188),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_194),
.B(n_176),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_239),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_199),
.B(n_195),
.C(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_197),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_236),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_179),
.B1(n_173),
.B2(n_170),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_216),
.C(n_210),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_168),
.C(n_173),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_240),
.C(n_211),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_168),
.B(n_174),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_207),
.B1(n_220),
.B2(n_201),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_181),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_16),
.C(n_13),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_232),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_229),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_217),
.C(n_216),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_252),
.C(n_256),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_229),
.B1(n_13),
.B2(n_14),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_202),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_209),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_241),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_233),
.B(n_227),
.C(n_230),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_236),
.B(n_218),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_210),
.C(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_219),
.C(n_220),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_225),
.C(n_240),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_255),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_262),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_233),
.B1(n_228),
.B2(n_222),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_249),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_226),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_225),
.B(n_223),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_269),
.B(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_266),
.C(n_242),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_276),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_249),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

INVx11_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_8),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_281),
.B(n_8),
.Y(n_287)
);

OAI321xp33_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_275),
.A3(n_279),
.B1(n_273),
.B2(n_264),
.C(n_271),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_266),
.B(n_15),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_14),
.C(n_15),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_268),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_280),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_289),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_286),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_282),
.C(n_289),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_16),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_16),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_299),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_294),
.B(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_298),
.C(n_288),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_301),
.Y(n_303)
);


endmodule