module fake_ariane_2285_n_259 (n_8, n_24, n_7, n_22, n_43, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_45, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_259);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_259;

wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_221;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_242;
wire n_115;
wire n_133;
wire n_66;
wire n_205;
wire n_236;
wire n_71;
wire n_109;
wire n_208;
wire n_245;
wire n_96;
wire n_156;
wire n_209;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_235;
wire n_225;
wire n_200;
wire n_51;
wire n_166;
wire n_253;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_244;
wire n_246;
wire n_226;
wire n_46;
wire n_220;
wire n_84;
wire n_247;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_224;
wire n_217;
wire n_240;
wire n_82;
wire n_178;
wire n_57;
wire n_131;
wire n_201;
wire n_229;
wire n_70;
wire n_250;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_256;
wire n_214;
wire n_227;
wire n_48;
wire n_101;
wire n_94;
wire n_243;
wire n_134;
wire n_188;
wire n_185;
wire n_249;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_255;
wire n_122;
wire n_257;
wire n_198;
wire n_148;
wire n_232;
wire n_164;
wire n_52;
wire n_248;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_258;
wire n_73;
wire n_77;
wire n_171;
wire n_228;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_241;
wire n_254;
wire n_238;
wire n_219;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_252;
wire n_142;
wire n_251;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_63;
wire n_59;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_54;

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_4),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

INVxp33_ASAP7_75t_SL g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_1),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_2),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_3),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_46),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_6),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_6),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_7),
.B(n_8),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_8),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_10),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_11),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_15),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_75),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_79),
.C(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

O2A1O1Ixp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_70),
.B(n_47),
.C(n_67),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_59),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_73),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_58),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_23),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_26),
.Y(n_119)
);

NOR2x1p5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_93),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_92),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_95),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_120),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_88),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_107),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_90),
.B(n_121),
.C(n_137),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_124),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_107),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_106),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_108),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_113),
.B(n_108),
.C(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_88),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_119),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_83),
.B1(n_91),
.B2(n_101),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_85),
.B(n_92),
.C(n_119),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_118),
.B(n_77),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_109),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_91),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_129),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g164 ( 
.A(n_145),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_133),
.B(n_94),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_101),
.B1(n_133),
.B2(n_87),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_148),
.B(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_129),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_156),
.B1(n_144),
.B2(n_154),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_149),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_172),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_173),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_147),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_179),
.B(n_164),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_145),
.B1(n_159),
.B2(n_149),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND4xp25_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_158),
.C(n_139),
.D(n_85),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_162),
.Y(n_197)
);

OAI33xp33_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_151),
.A3(n_170),
.B1(n_152),
.B2(n_94),
.B3(n_140),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_165),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_179),
.A2(n_94),
.B1(n_167),
.B2(n_171),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_186),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_168),
.B(n_180),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_183),
.B1(n_189),
.B2(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_200),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_186),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_183),
.Y(n_210)
);

NAND2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_187),
.Y(n_211)
);

NAND2x1p5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_187),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_183),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_182),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_198),
.C(n_180),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_184),
.Y(n_216)
);

AOI31xp33_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_197),
.A3(n_201),
.B(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_189),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_187),
.Y(n_220)
);

NOR2x1_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

NAND2x1_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_189),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_168),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_175),
.Y(n_228)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_187),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_189),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_187),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_184),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

NOR3xp33_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_217),
.C(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_228),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_233),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_242),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_241),
.Y(n_249)
);

OAI211xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_226),
.B(n_230),
.C(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_217),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_182),
.B1(n_180),
.B2(n_165),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_157),
.C(n_35),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

NOR3xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_166),
.C(n_36),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_257),
.B(n_255),
.Y(n_259)
);


endmodule