module fake_jpeg_637_n_209 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_209);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_7),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_6),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_0),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_84),
.Y(n_98)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_51),
.Y(n_82)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_54),
.B1(n_61),
.B2(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_87),
.B1(n_81),
.B2(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_54),
.B1(n_80),
.B2(n_76),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_50),
.B(n_69),
.C(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_62),
.B1(n_63),
.B2(n_75),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_55),
.B1(n_51),
.B2(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_61),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_83),
.B1(n_80),
.B2(n_76),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_100),
.A2(n_108),
.B1(n_111),
.B2(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_106),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_89),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_81),
.B1(n_75),
.B2(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_109),
.B1(n_52),
.B2(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_73),
.B1(n_72),
.B2(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_113),
.Y(n_129)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_58),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_55),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_97),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_117),
.Y(n_122)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_57),
.C(n_67),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_130),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_126),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_57),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_0),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_135),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_97),
.C(n_24),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_104),
.C(n_117),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_1),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_1),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_147)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_151),
.A2(n_161),
.B1(n_36),
.B2(n_46),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_32),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_12),
.B(n_14),
.Y(n_157)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_159),
.B(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_34),
.B1(n_47),
.B2(n_20),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_136),
.B1(n_123),
.B2(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_171),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_31),
.C(n_44),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_15),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_163),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_29),
.C(n_22),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_162),
.B(n_152),
.C(n_155),
.D(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_183),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_175),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_158),
.B(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_16),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_179),
.B(n_167),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_168),
.B(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_194),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_181),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_197),
.A2(n_190),
.B1(n_170),
.B2(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_192),
.B(n_199),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_204),
.A2(n_202),
.B(n_195),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_200),
.B(n_193),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_187),
.A3(n_16),
.B1(n_25),
.B2(n_27),
.C1(n_28),
.C2(n_39),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_23),
.C(n_41),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_43),
.Y(n_209)
);


endmodule