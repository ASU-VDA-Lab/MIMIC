module fake_netlist_6_4793_n_15 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_15);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;

output n_15;

wire n_14;
wire n_13;
wire n_10;
wire n_9;
wire n_11;
wire n_8;
wire n_12;

INVxp67_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

AOI332xp33_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_8),
.A3(n_0),
.B1(n_3),
.B2(n_4),
.B3(n_2),
.C1(n_6),
.C2(n_7),
.Y(n_12)
);

AND2x4_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);


endmodule