module fake_aes_12587_n_629 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_629);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_629;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_17), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_14), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_58), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_82), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_6), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_32), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_28), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_22), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_23), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_68), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_0), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_73), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_11), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_65), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_33), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_47), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_24), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_56), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_5), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_20), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_44), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_49), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_66), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_79), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_67), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_64), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_71), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_9), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_7), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_63), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_46), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_18), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_61), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_17), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_54), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_89), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_70), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_19), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_26), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_98), .B(n_0), .Y(n_135) );
BUFx12f_ASAP7_75t_L g136 ( .A(n_98), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_123), .B(n_1), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_99), .B(n_1), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_101), .B(n_25), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_101), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_104), .B(n_2), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_99), .B(n_2), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_104), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_106), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_123), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_129), .Y(n_146) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_134), .A2(n_3), .B(n_4), .Y(n_147) );
BUFx8_ASAP7_75t_L g148 ( .A(n_106), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_106), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_134), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_133), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_151) );
BUFx12f_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_115), .B(n_6), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_106), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_136), .B(n_111), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_136), .B(n_94), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_136), .B(n_96), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_146), .B(n_92), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_147), .Y(n_159) );
OAI21xp33_ASAP7_75t_L g160 ( .A1(n_140), .A2(n_129), .B(n_103), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_147), .Y(n_161) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
OR2x2_ASAP7_75t_L g165 ( .A(n_146), .B(n_91), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
AND2x6_ASAP7_75t_L g169 ( .A(n_137), .B(n_93), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_137), .B(n_127), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_148), .Y(n_171) );
INVxp67_ASAP7_75t_SL g172 ( .A(n_135), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_140), .B(n_91), .Y(n_173) );
INVxp33_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_151), .B(n_100), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_143), .B(n_102), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_148), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_172), .B(n_152), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_170), .B(n_153), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_169), .A2(n_137), .B1(n_139), .B2(n_153), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_174), .A2(n_125), .B1(n_121), .B2(n_131), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_143), .B(n_135), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_171), .B(n_152), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_155), .B(n_137), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_169), .A2(n_137), .B1(n_139), .B2(n_141), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_173), .B(n_138), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_165), .B(n_138), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_180), .B(n_142), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_171), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_169), .B(n_142), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_181), .B(n_96), .Y(n_200) );
INVx5_ASAP7_75t_L g201 ( .A(n_181), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_169), .B(n_112), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_179), .Y(n_204) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_162), .B(n_97), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_178), .B(n_150), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_169), .B(n_112), .Y(n_208) );
INVxp67_ASAP7_75t_R g209 ( .A(n_169), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_169), .A2(n_139), .B1(n_141), .B2(n_150), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_158), .B(n_130), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_177), .A2(n_151), .B1(n_139), .B2(n_100), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_170), .B(n_145), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_170), .B(n_150), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_190), .A2(n_162), .B(n_176), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_193), .A2(n_160), .B(n_170), .C(n_163), .Y(n_218) );
AOI21x1_ASAP7_75t_L g219 ( .A1(n_190), .A2(n_167), .B(n_176), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_184), .B(n_156), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_194), .B(n_177), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_188), .A2(n_167), .B(n_139), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_194), .B(n_177), .Y(n_223) );
AND2x2_ASAP7_75t_SL g224 ( .A(n_205), .B(n_103), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_185), .A2(n_177), .B1(n_90), .B2(n_105), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_216), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_206), .B(n_157), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g228 ( .A1(n_197), .A2(n_107), .B(n_108), .C(n_109), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_213), .A2(n_160), .B1(n_102), .B2(n_133), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_191), .A2(n_150), .B(n_145), .C(n_114), .Y(n_230) );
NOR2x1_ASAP7_75t_L g231 ( .A(n_182), .B(n_95), .Y(n_231) );
NOR2x1_ASAP7_75t_L g232 ( .A(n_195), .B(n_113), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_216), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_215), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_198), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_183), .B(n_211), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_197), .A2(n_164), .B(n_168), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_202), .A2(n_164), .B(n_168), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_212), .A2(n_124), .B(n_122), .C(n_127), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_202), .A2(n_164), .B(n_175), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_183), .B(n_130), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_204), .A2(n_175), .B(n_166), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_183), .A2(n_139), .B1(n_148), .B2(n_116), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_204), .A2(n_166), .B(n_126), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_187), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_214), .A2(n_120), .B(n_110), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_183), .B(n_132), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_214), .A2(n_128), .B(n_117), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_223), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_239), .A2(n_199), .B(n_189), .C(n_207), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_217), .A2(n_196), .B(n_186), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_235), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_222), .A2(n_196), .B(n_186), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_236), .A2(n_212), .B(n_192), .C(n_210), .Y(n_255) );
NOR4xp25_ASAP7_75t_L g256 ( .A(n_239), .B(n_118), .C(n_119), .D(n_154), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_235), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_196), .B(n_186), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_234), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g260 ( .A(n_224), .B(n_198), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_238), .A2(n_200), .B(n_154), .Y(n_261) );
AO22x2_ASAP7_75t_L g262 ( .A1(n_225), .A2(n_215), .B1(n_207), .B2(n_208), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_235), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_223), .B(n_215), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_230), .A2(n_215), .B(n_203), .C(n_154), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_218), .A2(n_205), .B(n_139), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_218), .A2(n_154), .A3(n_198), .B(n_139), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_221), .B(n_209), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_233), .B(n_205), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_230), .A2(n_201), .B(n_132), .C(n_106), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_240), .A2(n_198), .B(n_201), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_232), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_258), .A2(n_228), .B(n_244), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_250), .A2(n_243), .B(n_246), .Y(n_276) );
OR2x6_ASAP7_75t_L g277 ( .A(n_262), .B(n_248), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_253), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_254), .Y(n_279) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_263), .B(n_241), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_255), .A2(n_242), .B(n_231), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_267), .B(n_201), .Y(n_282) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_252), .A2(n_247), .B(n_245), .Y(n_283) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_252), .A2(n_245), .B(n_228), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_259), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_267), .B(n_224), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_260), .B(n_201), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_270), .B(n_220), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_262), .B(n_227), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_264), .B(n_249), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_254), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_253), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_263), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_250), .A2(n_229), .B(n_139), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_253), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_275), .B(n_262), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_285), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_289), .B(n_262), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_274), .A2(n_266), .B(n_256), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_292), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_281), .A2(n_256), .B(n_265), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_292), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_289), .B(n_273), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_274), .A2(n_266), .B(n_250), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_295), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_289), .B(n_268), .Y(n_313) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_291), .A2(n_271), .B(n_261), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_268), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_289), .B(n_268), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_289), .B(n_268), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_289), .B(n_268), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_313), .B(n_277), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_313), .B(n_283), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_318), .B(n_286), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_296), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_313), .B(n_277), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_315), .B(n_283), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_315), .B(n_283), .Y(n_331) );
NOR2x1_ASAP7_75t_SL g332 ( .A(n_299), .B(n_277), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_315), .B(n_283), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_301), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_298), .B(n_283), .Y(n_336) );
NOR2x1_ASAP7_75t_SL g337 ( .A(n_299), .B(n_277), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_298), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_309), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_301), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_318), .B(n_286), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_299), .A2(n_260), .B1(n_288), .B2(n_290), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_300), .B(n_283), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_309), .B(n_277), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_307), .B(n_277), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_316), .B(n_277), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_316), .B(n_284), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_303), .B(n_288), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_310), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_316), .B(n_284), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_317), .B(n_284), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_312), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_303), .B(n_284), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_305), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_306), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_307), .B(n_284), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_299), .A2(n_280), .B1(n_269), .B2(n_273), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_307), .B(n_273), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_306), .B(n_281), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_312), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_332), .B(n_299), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_324), .B(n_317), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_347), .B(n_297), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_327), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_340), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_358), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_358), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_359), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_352), .B(n_311), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_325), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_349), .B(n_317), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_347), .B(n_297), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_363), .B(n_321), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_332), .B(n_321), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_324), .B(n_321), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_329), .B(n_322), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_329), .B(n_322), .Y(n_384) );
NAND2xp67_ASAP7_75t_L g385 ( .A(n_352), .B(n_312), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_331), .B(n_319), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_331), .B(n_319), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_333), .B(n_319), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_340), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_350), .B(n_320), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_325), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_350), .B(n_320), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_335), .B(n_287), .Y(n_394) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_349), .B(n_311), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_330), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_338), .B(n_304), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_338), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_346), .B(n_308), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_354), .B(n_308), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_354), .B(n_308), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_339), .B(n_304), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_335), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_355), .B(n_308), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_339), .B(n_302), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_355), .B(n_302), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_323), .B(n_302), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_346), .B(n_302), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_334), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_334), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_334), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_326), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_341), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_342), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_364), .B(n_302), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_341), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_361), .B(n_314), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_341), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_323), .B(n_314), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_344), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_344), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_361), .B(n_314), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_323), .B(n_314), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_323), .B(n_314), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_367), .B(n_343), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_368), .B(n_328), .Y(n_428) );
NOR2xp33_ASAP7_75t_SL g429 ( .A(n_395), .B(n_280), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_414), .A2(n_328), .B1(n_348), .B2(n_362), .C(n_336), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_368), .B(n_328), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_416), .B(n_343), .Y(n_432) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_403), .B(n_336), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_397), .A2(n_348), .B1(n_345), .B2(n_357), .C(n_149), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_393), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_379), .B(n_351), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_382), .B(n_348), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_366), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_369), .B(n_351), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_389), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_407), .B(n_337), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_383), .B(n_357), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_367), .B(n_337), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_376), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_407), .B(n_351), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_408), .B(n_353), .Y(n_447) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_381), .B(n_353), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_383), .B(n_365), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_384), .B(n_353), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_370), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_385), .Y(n_452) );
NOR2x1p5_ASAP7_75t_L g453 ( .A(n_403), .B(n_356), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_386), .B(n_365), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_387), .B(n_365), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_387), .B(n_8), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_375), .B(n_8), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_381), .B(n_287), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_381), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_396), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_402), .B(n_9), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_396), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_372), .B(n_10), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_398), .Y(n_464) );
OR2x6_ASAP7_75t_L g465 ( .A(n_377), .B(n_293), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_398), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_388), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_373), .B(n_12), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_394), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_400), .B(n_149), .Y(n_471) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_377), .B(n_282), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_376), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_371), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_394), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_400), .B(n_149), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_411), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_374), .B(n_13), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_380), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_401), .B(n_149), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_385), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_401), .B(n_15), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_378), .B(n_15), .Y(n_484) );
INVx4_ASAP7_75t_L g485 ( .A(n_394), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_377), .B(n_16), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_380), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_405), .B(n_16), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_413), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_415), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_391), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_378), .B(n_390), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_467), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_438), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_446), .B(n_406), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
AOI222xp33_ASAP7_75t_L g497 ( .A1(n_484), .A2(n_405), .B1(n_417), .B2(n_426), .C1(n_425), .C2(n_421), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_446), .B(n_409), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_428), .B(n_421), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_428), .B(n_425), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_448), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_443), .B(n_409), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_492), .B(n_390), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_431), .B(n_426), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_448), .Y(n_506) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_465), .A2(n_424), .B1(n_419), .B2(n_399), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_490), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_465), .A2(n_391), .B(n_410), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_486), .A2(n_392), .B1(n_399), .B2(n_420), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_462), .Y(n_512) );
OAI21xp33_ASAP7_75t_L g513 ( .A1(n_442), .A2(n_423), .B(n_422), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_471), .B(n_418), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_441), .B(n_420), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_490), .Y(n_516) );
OAI21xp5_ASAP7_75t_SL g517 ( .A1(n_472), .A2(n_423), .B(n_422), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_464), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_466), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_482), .B(n_18), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_469), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_453), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_450), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_477), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_488), .B(n_484), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_430), .A2(n_412), .B1(n_290), .B2(n_293), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_452), .Y(n_527) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_465), .B(n_282), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_437), .B(n_149), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_449), .B(n_149), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_441), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_481), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_476), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_427), .A2(n_293), .B1(n_276), .B2(n_282), .Y(n_534) );
AOI322xp5_ASAP7_75t_L g535 ( .A1(n_456), .A2(n_20), .A3(n_21), .B1(n_22), .B2(n_23), .C1(n_269), .C2(n_282), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_459), .B(n_21), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_459), .B(n_276), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_480), .B(n_276), .Y(n_538) );
NOR2xp67_ASAP7_75t_L g539 ( .A(n_459), .B(n_27), .Y(n_539) );
NAND2x1_ASAP7_75t_L g540 ( .A(n_444), .B(n_282), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_491), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_480), .B(n_276), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_461), .B(n_29), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g544 ( .A(n_485), .B(n_30), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_447), .B(n_268), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_491), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_483), .B(n_294), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_540), .A2(n_429), .B(n_433), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_497), .B(n_474), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_497), .B(n_474), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_517), .A2(n_526), .B1(n_513), .B2(n_511), .C(n_532), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_531), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_525), .A2(n_432), .B1(n_458), .B2(n_434), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_515), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_515), .Y(n_555) );
AOI31xp33_ASAP7_75t_L g556 ( .A1(n_536), .A2(n_435), .A3(n_458), .B(n_470), .Y(n_556) );
AOI21xp33_ASAP7_75t_SL g557 ( .A1(n_507), .A2(n_475), .B(n_436), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_494), .B(n_457), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_496), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_536), .B(n_485), .Y(n_560) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_510), .A2(n_473), .B(n_445), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_530), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_520), .A2(n_478), .B1(n_463), .B2(n_468), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_499), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_541), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_500), .B(n_454), .Y(n_566) );
AOI32xp33_ASAP7_75t_L g567 ( .A1(n_493), .A2(n_455), .A3(n_489), .B1(n_440), .B2(n_487), .Y(n_567) );
AOI22x1_ASAP7_75t_SL g568 ( .A1(n_502), .A2(n_473), .B1(n_445), .B2(n_479), .Y(n_568) );
AO221x1_ASAP7_75t_L g569 ( .A1(n_507), .A2(n_479), .B1(n_257), .B2(n_294), .C(n_35), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_533), .A2(n_294), .B1(n_257), .B2(n_148), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_501), .B(n_31), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_527), .A2(n_251), .B(n_272), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_546), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_505), .B(n_34), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_506), .A2(n_36), .B1(n_37), .B2(n_38), .C(n_40), .Y(n_575) );
OAI221xp5_ASAP7_75t_SL g576 ( .A1(n_535), .A2(n_41), .B1(n_42), .B2(n_45), .C(n_48), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_522), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_529), .Y(n_578) );
OAI221xp5_ASAP7_75t_L g579 ( .A1(n_549), .A2(n_503), .B1(n_495), .B2(n_498), .C(n_509), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_550), .A2(n_495), .B1(n_523), .B2(n_534), .C(n_521), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_557), .A2(n_534), .B1(n_508), .B2(n_512), .C(n_518), .Y(n_581) );
OAI32xp33_ASAP7_75t_L g582 ( .A1(n_560), .A2(n_504), .A3(n_516), .B1(n_498), .B2(n_514), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_578), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_551), .A2(n_543), .B(n_519), .C(n_524), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g585 ( .A1(n_556), .A2(n_537), .B(n_545), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_568), .A2(n_542), .B1(n_538), .B2(n_547), .Y(n_586) );
OAI222xp33_ASAP7_75t_L g587 ( .A1(n_567), .A2(n_539), .B1(n_544), .B2(n_53), .C1(n_55), .C2(n_57), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_560), .A2(n_59), .B(n_60), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_558), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_559), .Y(n_590) );
OAI31xp33_ASAP7_75t_L g591 ( .A1(n_548), .A2(n_72), .A3(n_74), .B(n_75), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_566), .B(n_76), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_569), .A2(n_77), .B1(n_78), .B2(n_80), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_553), .A2(n_81), .B1(n_83), .B2(n_84), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_558), .A2(n_85), .B1(n_86), .B2(n_87), .C(n_88), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_561), .A2(n_575), .B(n_562), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_564), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_561), .A2(n_562), .B(n_576), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_553), .A2(n_554), .B1(n_555), .B2(n_563), .C(n_552), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_561), .A2(n_574), .B(n_571), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_565), .A2(n_573), .B1(n_572), .B2(n_577), .C(n_570), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_565), .B(n_557), .C(n_550), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_573), .A2(n_550), .B(n_549), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_549), .A2(n_550), .B(n_557), .C(n_551), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_549), .B(n_550), .Y(n_605) );
AND4x1_ASAP7_75t_L g606 ( .A(n_548), .B(n_549), .C(n_550), .D(n_528), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_597), .Y(n_607) );
NOR2x1_ASAP7_75t_L g608 ( .A(n_587), .B(n_584), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_604), .B(n_605), .C(n_603), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_599), .A2(n_580), .B1(n_602), .B2(n_582), .C(n_579), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_596), .A2(n_587), .B(n_585), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_590), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_609), .B(n_591), .C(n_593), .D(n_588), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_608), .B(n_595), .C(n_581), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_611), .B(n_583), .Y(n_615) );
NOR2x1p5_ASAP7_75t_L g616 ( .A(n_607), .B(n_606), .Y(n_616) );
XOR2xp5_ASAP7_75t_L g617 ( .A(n_613), .B(n_592), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_615), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_614), .B(n_612), .Y(n_619) );
XNOR2xp5_ASAP7_75t_L g620 ( .A(n_617), .B(n_616), .Y(n_620) );
INVx2_ASAP7_75t_SL g621 ( .A(n_618), .Y(n_621) );
OA21x2_ASAP7_75t_L g622 ( .A1(n_620), .A2(n_619), .B(n_610), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_621), .Y(n_623) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_623), .Y(n_624) );
XOR2xp5_ASAP7_75t_L g625 ( .A(n_622), .B(n_594), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_624), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_626), .A2(n_625), .B(n_622), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_627), .A2(n_589), .B(n_598), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_628), .A2(n_586), .B1(n_601), .B2(n_600), .Y(n_629) );
endmodule