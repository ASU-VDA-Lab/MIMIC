module fake_jpeg_24872_n_319 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_23),
.B1(n_20),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_36),
.B1(n_23),
.B2(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_23),
.B1(n_26),
.B2(n_20),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_36),
.B1(n_26),
.B2(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_26),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_69),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_67),
.B1(n_52),
.B2(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_36),
.B1(n_20),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_66),
.B1(n_72),
.B2(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2x1p5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_16),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_16),
.C(n_42),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_32),
.B1(n_37),
.B2(n_34),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_33),
.B(n_37),
.C(n_31),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_90),
.B1(n_96),
.B2(n_94),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_87),
.B1(n_91),
.B2(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_90),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_69),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_67),
.C(n_61),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_29),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_115),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_107),
.B1(n_34),
.B2(n_33),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_108),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_59),
.B(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_65),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_79),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_73),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_119),
.B(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_120),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_117),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_85),
.B(n_86),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_125),
.B(n_141),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_89),
.B1(n_73),
.B2(n_51),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_136),
.B1(n_34),
.B2(n_54),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_53),
.B(n_55),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_35),
.B1(n_41),
.B2(n_50),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_130),
.B1(n_62),
.B2(n_63),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_41),
.B1(n_49),
.B2(n_29),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_135),
.Y(n_153)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_99),
.C(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_44),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_29),
.B(n_51),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_101),
.B(n_14),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_151),
.C(n_171),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_62),
.B1(n_54),
.B2(n_93),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_149),
.B(n_167),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_31),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_115),
.C(n_110),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_168),
.B1(n_130),
.B2(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_165),
.Y(n_176)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_169),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_126),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_124),
.A2(n_110),
.B1(n_107),
.B2(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_107),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_80),
.B(n_70),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_119),
.C(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_170),
.B1(n_171),
.B2(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_137),
.C(n_142),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_186),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_145),
.B1(n_123),
.B2(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_187),
.B1(n_195),
.B2(n_199),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_125),
.C(n_144),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_192),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_131),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_189),
.B(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_136),
.B1(n_144),
.B2(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_165),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_158),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_121),
.B1(n_117),
.B2(n_93),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_54),
.B1(n_148),
.B2(n_80),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_195),
.B1(n_196),
.B2(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_103),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_155),
.B(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_217),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_187),
.B1(n_184),
.B2(n_190),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_219),
.B1(n_177),
.B2(n_191),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_155),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_209),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_215),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_157),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_158),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_188),
.C(n_176),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_182),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_218),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_31),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_31),
.C(n_17),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_230),
.B1(n_219),
.B2(n_211),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_229),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_176),
.C(n_188),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_232),
.C(n_236),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_182),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_181),
.B1(n_183),
.B2(n_197),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_220),
.C(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_210),
.C(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_95),
.C(n_58),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_241),
.C(n_242),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_34),
.B1(n_21),
.B2(n_27),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_240),
.B1(n_224),
.B2(n_235),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_28),
.C(n_22),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_21),
.B1(n_27),
.B2(n_95),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_68),
.C(n_44),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_68),
.C(n_44),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_247),
.B(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_28),
.B1(n_22),
.B2(n_17),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_246),
.A2(n_239),
.B1(n_25),
.B2(n_15),
.Y(n_275)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_10),
.B(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_242),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_254),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_10),
.B(n_12),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_0),
.B(n_2),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_24),
.Y(n_256)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_11),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_10),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_0),
.C(n_1),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_259),
.C(n_222),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_0),
.C(n_1),
.Y(n_259)
);

NOR2x1_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_11),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_3),
.B(n_4),
.Y(n_277)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_251),
.C(n_253),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_273),
.C(n_276),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_251),
.C(n_222),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_28),
.B1(n_22),
.B2(n_17),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_285),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_259),
.C(n_246),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_286),
.C(n_287),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_243),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_273),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_268),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_248),
.B1(n_247),
.B2(n_255),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_276),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_25),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_3),
.Y(n_296)
);

AOI31xp67_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_265),
.A3(n_274),
.B(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_298),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_267),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_294),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_4),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_15),
.B(n_25),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_300),
.B(n_4),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_3),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_287),
.C(n_284),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_5),
.C(n_7),
.Y(n_308)
);

NAND4xp25_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_305),
.B(n_301),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_5),
.B(n_6),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_299),
.B(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_304),
.C(n_302),
.Y(n_313)
);

NAND2x1p5_ASAP7_75t_SL g315 ( 
.A(n_313),
.B(n_309),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_314),
.B(n_7),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_7),
.B(n_8),
.C(n_307),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_7),
.B1(n_8),
.B2(n_265),
.Y(n_319)
);


endmodule