module fake_jpeg_17429_n_164 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_32),
.B(n_35),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_33),
.A2(n_45),
.B1(n_20),
.B2(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_15),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_34),
.A2(n_31),
.B(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_42),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_6),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_8),
.B1(n_11),
.B2(n_25),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_29),
.B1(n_31),
.B2(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_48),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_17),
.A2(n_11),
.B1(n_27),
.B2(n_25),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.Y(n_58)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_64),
.Y(n_102)
);

AO21x2_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_14),
.B(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_74),
.B1(n_39),
.B2(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_71),
.Y(n_83)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_56),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_78),
.B(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_79),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_22),
.B(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_88),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_41),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_86),
.B1(n_70),
.B2(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_71),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_76),
.C(n_60),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_75),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_103),
.B(n_85),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_54),
.B1(n_82),
.B2(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_59),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_73),
.B1(n_69),
.B2(n_67),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_69),
.B(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_114),
.B1(n_115),
.B2(n_121),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_64),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_117),
.B(n_118),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_70),
.B1(n_67),
.B2(n_75),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_83),
.B1(n_86),
.B2(n_103),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_70),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_87),
.C(n_88),
.Y(n_119)
);

NOR4xp25_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_97),
.C(n_90),
.D(n_93),
.Y(n_126)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_90),
.B(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_99),
.B1(n_100),
.B2(n_89),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_130),
.B1(n_132),
.B2(n_114),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_129),
.C(n_107),
.Y(n_136)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_119),
.B1(n_121),
.B2(n_115),
.C(n_117),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_97),
.Y(n_129)
);

AO21x2_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_104),
.B(n_95),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.C(n_122),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_141),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_144),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_130),
.B(n_132),
.C(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_113),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_130),
.B1(n_113),
.B2(n_124),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_130),
.B1(n_125),
.B2(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_147),
.B1(n_136),
.B2(n_137),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_152),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_144),
.C(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_148),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_156),
.B1(n_149),
.B2(n_152),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_131),
.B1(n_120),
.B2(n_110),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_131),
.B(n_139),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_146),
.C(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.C(n_155),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_151),
.C(n_153),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.Y(n_164)
);


endmodule