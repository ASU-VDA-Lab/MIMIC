module fake_netlist_5_2133_n_2373 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2373);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2373;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_901;
wire n_553;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_604;
wire n_368;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_331;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_378;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2340;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_1138;
wire n_364;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_92),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_124),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_70),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_40),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_94),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_108),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_133),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_84),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_43),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_67),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_145),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_109),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_146),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_82),
.Y(n_244)
);

INVx4_ASAP7_75t_R g245 ( 
.A(n_113),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_102),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_207),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_135),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_198),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_216),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_68),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_174),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_181),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_69),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_10),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_5),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_121),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_96),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_52),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_191),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_1),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_3),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_139),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_103),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_67),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_152),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_88),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_137),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_128),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_21),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_95),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_98),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_160),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_100),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_28),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_78),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_76),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_48),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_116),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_47),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_16),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_31),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_61),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_123),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_81),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_51),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_212),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_150),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_7),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_193),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_50),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_136),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_166),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_84),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_177),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_114),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_49),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_39),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_132),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_184),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_220),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_125),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_28),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_129),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_223),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_26),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_96),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_70),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_187),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_37),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_119),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_57),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_47),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_13),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_143),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_41),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_189),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_115),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_205),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_213),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_61),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_24),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_211),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_208),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_105),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_37),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_176),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_56),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_7),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_200),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_44),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_110),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_78),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_30),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_42),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_16),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_48),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_83),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_88),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_89),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_173),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_131),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_161),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_162),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_86),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_134),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_65),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_202),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_74),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_83),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_195),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_42),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_12),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_81),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_8),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_55),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_43),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_50),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_117),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_27),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_126),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_33),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_141),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_23),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_91),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_66),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_217),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_4),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_54),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_107),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_199),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_45),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_20),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_151),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_169),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_178),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_112),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_77),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_26),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_165),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_46),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_196),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_53),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_39),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_10),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_164),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_192),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_122),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_73),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_167),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_27),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_46),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_140),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_18),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_2),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_19),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_186),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_95),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_5),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_98),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_77),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_2),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_35),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_75),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_73),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_82),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_111),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_120),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_30),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_156),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_197),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_17),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_62),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_8),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_203),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_19),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_59),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_13),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_18),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_185),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_190),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_127),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_53),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_32),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_4),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_180),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_94),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_215),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_159),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_72),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_72),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_62),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_63),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_25),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_64),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_69),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_71),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_236),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_228),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_292),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_232),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_292),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_246),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_292),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_234),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_292),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_249),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_240),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_299),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_292),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_242),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_243),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_316),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_292),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_230),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_229),
.B(n_261),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_316),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_230),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_230),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_0),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_231),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_231),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_254),
.Y(n_472)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_237),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_247),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_248),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_231),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_250),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_332),
.B(n_0),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_332),
.B(n_1),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_436),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_255),
.B(n_3),
.Y(n_482)
);

BUFx2_ASAP7_75t_SL g483 ( 
.A(n_320),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_253),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_431),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_296),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_436),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_229),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_261),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_296),
.Y(n_490)
);

BUFx6f_ASAP7_75t_SL g491 ( 
.A(n_235),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_263),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_263),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_421),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_266),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_L g497 ( 
.A(n_359),
.B(n_6),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_266),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_268),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_305),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_443),
.B(n_6),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_333),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_268),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_271),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_415),
.Y(n_505)
);

BUFx2_ASAP7_75t_SL g506 ( 
.A(n_349),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_427),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_257),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_271),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_280),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_258),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_276),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_276),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_251),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_432),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_262),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_281),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_235),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_281),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_280),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_265),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_251),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_282),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_235),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_272),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_279),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_235),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_282),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_285),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_283),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_283),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_251),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_284),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_233),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_291),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_284),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_290),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_290),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_302),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_267),
.B(n_9),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_304),
.Y(n_542)
);

CKINVDCx14_ASAP7_75t_R g543 ( 
.A(n_360),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_308),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_309),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_334),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_294),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_233),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_294),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_310),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_311),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_313),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_300),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_314),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_300),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_303),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_267),
.B(n_9),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_303),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_318),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_324),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_306),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_269),
.B(n_11),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_326),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_328),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_306),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_L g566 ( 
.A(n_446),
.B(n_11),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_449),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_510),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_449),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_451),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_R g571 ( 
.A(n_543),
.B(n_329),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_448),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_514),
.B(n_334),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_453),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_453),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_455),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_510),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_483),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_455),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_483),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_533),
.B(n_334),
.Y(n_583)
);

NOR2x1_ASAP7_75t_L g584 ( 
.A(n_459),
.B(n_402),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_459),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_546),
.B(n_339),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_463),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_450),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_515),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_R g590 ( 
.A(n_478),
.B(n_227),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_463),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_454),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_521),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_522),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_535),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_521),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_457),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_488),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_489),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_489),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_464),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_516),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_535),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_492),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_467),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_479),
.B(n_252),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_530),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_492),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_493),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_505),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_535),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_462),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_467),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_468),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_R g617 ( 
.A(n_460),
.B(n_341),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_548),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_493),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_496),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_480),
.B(n_350),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_461),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_496),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_480),
.B(n_353),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_507),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_474),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_498),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_548),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_482),
.B(n_252),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_540),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_468),
.Y(n_631)
);

OA21x2_ASAP7_75t_L g632 ( 
.A1(n_470),
.A2(n_270),
.B(n_241),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_481),
.B(n_402),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_559),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_466),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_470),
.A2(n_270),
.B(n_241),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_498),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_447),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_471),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_486),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_471),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_519),
.B(n_238),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_481),
.B(n_402),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_456),
.Y(n_645)
);

CKINVDCx8_ASAP7_75t_R g646 ( 
.A(n_525),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_487),
.B(n_355),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_476),
.B(n_241),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_476),
.B(n_270),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_458),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_500),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_502),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_485),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_475),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_548),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_477),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_490),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_499),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_503),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_491),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_548),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_633),
.B(n_487),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_568),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_618),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_574),
.B(n_523),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_593),
.Y(n_666)
);

AND3x2_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_557),
.C(n_541),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_633),
.B(n_523),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_633),
.B(n_269),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_644),
.B(n_274),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_593),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_586),
.B(n_484),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_593),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_596),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_596),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_567),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_574),
.B(n_497),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_574),
.B(n_506),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_569),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_618),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_608),
.B(n_629),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_586),
.B(n_508),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_598),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_618),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_583),
.B(n_506),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_567),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_618),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_618),
.Y(n_690)
);

INVxp67_ASAP7_75t_SL g691 ( 
.A(n_655),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_570),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_618),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_570),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_644),
.B(n_274),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_569),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_608),
.B(n_511),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_657),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_570),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_629),
.B(n_517),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_572),
.Y(n_701)
);

AO22x2_ASAP7_75t_L g702 ( 
.A1(n_589),
.A2(n_495),
.B1(n_494),
.B2(n_349),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_583),
.B(n_526),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_583),
.B(n_644),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_655),
.B(n_527),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_618),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_584),
.B(n_275),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_573),
.B(n_536),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_618),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_572),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_584),
.B(n_275),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_657),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_578),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_590),
.A2(n_472),
.B1(n_452),
.B2(n_542),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_655),
.B(n_544),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_621),
.B(n_503),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_568),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_621),
.B(n_504),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_568),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_632),
.A2(n_562),
.B1(n_566),
.B2(n_501),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_598),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_599),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

BUFx6f_ASAP7_75t_SL g724 ( 
.A(n_660),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_600),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_600),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_571),
.B(n_528),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_588),
.B(n_545),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_646),
.B(n_406),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_601),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_577),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_605),
.B(n_550),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_568),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_575),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_648),
.B(n_649),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_568),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_624),
.B(n_504),
.Y(n_738)
);

BUFx4f_ASAP7_75t_L g739 ( 
.A(n_632),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_601),
.Y(n_740)
);

INVxp33_ASAP7_75t_L g741 ( 
.A(n_614),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_624),
.B(n_509),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_568),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_575),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_605),
.B(n_613),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_592),
.B(n_551),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_606),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_605),
.B(n_552),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_606),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_597),
.B(n_554),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_622),
.B(n_560),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_614),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_647),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_647),
.B(n_509),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_635),
.B(n_473),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_605),
.B(n_563),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_635),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_628),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_605),
.B(n_564),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_589),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_568),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_575),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_578),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_587),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_604),
.B(n_465),
.Y(n_765)
);

AND2x6_ASAP7_75t_L g766 ( 
.A(n_613),
.B(n_352),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_571),
.B(n_360),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_648),
.B(n_297),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_604),
.B(n_465),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_587),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_610),
.B(n_512),
.Y(n_771)
);

BUFx4_ASAP7_75t_L g772 ( 
.A(n_646),
.Y(n_772)
);

AO22x2_ASAP7_75t_L g773 ( 
.A1(n_643),
.A2(n_352),
.B1(n_370),
.B2(n_238),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_576),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_613),
.B(n_233),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_576),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_579),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_617),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_579),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_628),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_576),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_626),
.B(n_491),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_579),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_610),
.B(n_512),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_628),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_617),
.B(n_654),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_612),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_632),
.Y(n_788)
);

OAI21xp33_ASAP7_75t_L g789 ( 
.A1(n_611),
.A2(n_426),
.B(n_381),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_590),
.A2(n_491),
.B1(n_406),
.B2(n_438),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_613),
.B(n_438),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_579),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_632),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_611),
.B(n_513),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_579),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_581),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_656),
.B(n_357),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_581),
.Y(n_798)
);

INVxp33_ASAP7_75t_SL g799 ( 
.A(n_580),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_656),
.A2(n_582),
.B1(n_580),
.B2(n_469),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_613),
.B(n_376),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_581),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_640),
.B(n_381),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_582),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_661),
.B(n_595),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_661),
.B(n_380),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_632),
.Y(n_807)
);

AO22x2_ASAP7_75t_L g808 ( 
.A1(n_648),
.A2(n_370),
.B1(n_352),
.B2(n_426),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_577),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_648),
.B(n_297),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_628),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_595),
.B(n_239),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_585),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_628),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_640),
.B(n_439),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_595),
.B(n_244),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_660),
.B(n_360),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_660),
.B(n_360),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_636),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_661),
.B(n_383),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_628),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_651),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_660),
.B(n_384),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_636),
.Y(n_824)
);

INVxp33_ASAP7_75t_L g825 ( 
.A(n_755),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_678),
.B(n_640),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_682),
.A2(n_704),
.B1(n_753),
.B2(n_773),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_680),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_771),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_L g830 ( 
.A(n_700),
.B(n_646),
.C(n_259),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_680),
.Y(n_831)
);

BUFx8_ASAP7_75t_L g832 ( 
.A(n_724),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_822),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_696),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_736),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_753),
.B(n_661),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_679),
.B(n_660),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_788),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_697),
.B(n_594),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_716),
.B(n_595),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_752),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_704),
.A2(n_619),
.B(n_623),
.C(n_620),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_696),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_701),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_679),
.B(n_661),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_822),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_716),
.B(n_595),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_771),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_701),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_718),
.B(n_577),
.Y(n_850)
);

NAND3xp33_ASAP7_75t_SL g851 ( 
.A(n_790),
.B(n_652),
.C(n_651),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_718),
.B(n_577),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_686),
.B(n_788),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_698),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_686),
.B(n_788),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_752),
.Y(n_856)
);

NOR2x1p5_ASAP7_75t_L g857 ( 
.A(n_755),
.B(n_652),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_738),
.B(n_648),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_738),
.B(n_742),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_773),
.A2(n_370),
.B1(n_636),
.B2(n_649),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_788),
.B(n_628),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_784),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_784),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_736),
.B(n_668),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_742),
.B(n_754),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_754),
.B(n_649),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_791),
.B(n_649),
.Y(n_867)
);

INVxp33_ASAP7_75t_L g868 ( 
.A(n_741),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_672),
.B(n_594),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_794),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_788),
.B(n_628),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_757),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_691),
.B(n_649),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_683),
.B(n_301),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_703),
.A2(n_619),
.B(n_623),
.C(n_620),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_793),
.B(n_233),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_668),
.B(n_627),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_819),
.A2(n_319),
.B(n_330),
.C(n_323),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_736),
.Y(n_879)
);

NOR2x2_ASAP7_75t_L g880 ( 
.A(n_769),
.B(n_295),
.Y(n_880)
);

OR2x2_ASAP7_75t_SL g881 ( 
.A(n_803),
.B(n_815),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_720),
.B(n_301),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_794),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_710),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_773),
.A2(n_636),
.B1(n_327),
.B2(n_351),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_819),
.A2(n_323),
.B(n_330),
.C(n_319),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_665),
.B(n_327),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_665),
.B(n_812),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_824),
.A2(n_343),
.B(n_347),
.C(n_344),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_SL g890 ( 
.A(n_705),
.B(n_317),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_678),
.A2(n_668),
.B1(n_662),
.B2(n_816),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_732),
.B(n_748),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_756),
.B(n_336),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_684),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_757),
.B(n_609),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_759),
.B(n_336),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_797),
.B(n_708),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_793),
.B(n_351),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_760),
.B(n_609),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_765),
.B(n_630),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_773),
.A2(n_636),
.B1(n_368),
.B2(n_385),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_793),
.B(n_233),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_760),
.B(n_630),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_710),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_793),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_793),
.B(n_368),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_801),
.A2(n_591),
.B(n_585),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_807),
.B(n_379),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_807),
.B(n_379),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_807),
.B(n_233),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_807),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_807),
.B(n_385),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_715),
.B(n_721),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_664),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_722),
.B(n_395),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_723),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_725),
.B(n_395),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_669),
.A2(n_397),
.B1(n_437),
.B2(n_416),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_726),
.B(n_397),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_769),
.B(n_634),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_678),
.A2(n_386),
.B1(n_391),
.B2(n_389),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_739),
.B(n_372),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_728),
.B(n_634),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_739),
.B(n_664),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_730),
.B(n_416),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_740),
.B(n_437),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_747),
.B(n_627),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_669),
.A2(n_435),
.B1(n_372),
.B2(n_356),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_669),
.A2(n_372),
.B1(n_435),
.B2(n_280),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_749),
.B(n_637),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_739),
.B(n_372),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_664),
.B(n_372),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_678),
.A2(n_396),
.B1(n_417),
.B2(n_399),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_664),
.B(n_372),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_662),
.B(n_637),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_824),
.B(n_641),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_662),
.A2(n_714),
.B1(n_695),
.B2(n_670),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_713),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_713),
.B(n_641),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_763),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_765),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_763),
.B(n_764),
.Y(n_942)
);

NAND2x1_ASAP7_75t_L g943 ( 
.A(n_664),
.B(n_245),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_764),
.B(n_658),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_770),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_770),
.B(n_658),
.Y(n_946)
);

BUFx8_ASAP7_75t_L g947 ( 
.A(n_724),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_670),
.B(n_659),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_768),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_670),
.B(n_659),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_695),
.B(n_585),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_695),
.B(n_707),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_SL g953 ( 
.A(n_681),
.B(n_435),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_681),
.B(n_435),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_768),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_746),
.B(n_638),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_L g957 ( 
.A(n_681),
.B(n_280),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_707),
.B(n_591),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_707),
.B(n_591),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_731),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_769),
.B(n_513),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_674),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_778),
.B(n_786),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_769),
.Y(n_964)
);

BUFx5_ASAP7_75t_L g965 ( 
.A(n_766),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_768),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_681),
.B(n_435),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_789),
.A2(n_344),
.B(n_347),
.C(n_343),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_SL g969 ( 
.A1(n_712),
.A2(n_645),
.B1(n_650),
.B2(n_638),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_711),
.B(n_602),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_681),
.B(n_435),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_667),
.A2(n_420),
.B1(n_424),
.B2(n_419),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_674),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_675),
.Y(n_974)
);

AND2x6_ASAP7_75t_L g975 ( 
.A(n_711),
.B(n_348),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_711),
.B(n_602),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_810),
.B(n_602),
.Y(n_977)
);

BUFx5_ASAP7_75t_L g978 ( 
.A(n_766),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_810),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_750),
.B(n_645),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_751),
.B(n_650),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_810),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_690),
.B(n_603),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_690),
.B(n_603),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_690),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_690),
.B(n_603),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_690),
.B(n_709),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_808),
.A2(n_280),
.B1(n_375),
.B2(n_392),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_L g989 ( 
.A(n_709),
.B(n_280),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_709),
.B(n_607),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_778),
.B(n_518),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_803),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_777),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_808),
.A2(n_280),
.B1(n_375),
.B2(n_392),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_804),
.B(n_518),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_709),
.B(n_607),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_709),
.B(n_280),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_731),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_806),
.B(n_607),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_828),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_838),
.B(n_685),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_838),
.B(n_685),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_R g1003 ( 
.A(n_833),
.B(n_653),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_859),
.A2(n_799),
.B1(n_729),
.B2(n_800),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_865),
.B(n_809),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_828),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_831),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_838),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_838),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_960),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_897),
.A2(n_799),
.B1(n_820),
.B2(n_766),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_SL g1012 ( 
.A(n_851),
.B(n_260),
.C(n_256),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_834),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_834),
.Y(n_1014)
);

AO21x1_ASAP7_75t_L g1015 ( 
.A1(n_882),
.A2(n_775),
.B(n_745),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_843),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_888),
.A2(n_766),
.B1(n_818),
.B2(n_817),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_892),
.B(n_809),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_843),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_846),
.B(n_653),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_844),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_844),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_960),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_975),
.A2(n_808),
.B1(n_766),
.B2(n_779),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_849),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_877),
.B(n_727),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_995),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_911),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_832),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_849),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_911),
.B(n_685),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_841),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_960),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_884),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_854),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_960),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_913),
.B(n_782),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_829),
.B(n_808),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_904),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_998),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_911),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_827),
.B(n_724),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_975),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_998),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_864),
.Y(n_1045)
);

AND2x6_ASAP7_75t_L g1046 ( 
.A(n_837),
.B(n_805),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_856),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_904),
.Y(n_1048)
);

CKINVDCx8_ASAP7_75t_R g1049 ( 
.A(n_826),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_914),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_940),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_940),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_835),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_991),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_895),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_877),
.B(n_823),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_864),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_914),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_848),
.B(n_862),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_992),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_945),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_SL g1062 ( 
.A(n_890),
.B(n_969),
.C(n_830),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_945),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_R g1064 ( 
.A(n_854),
.B(n_612),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_835),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_962),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_935),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_877),
.B(n_767),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_890),
.B(n_273),
.C(n_264),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_962),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_914),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_935),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_935),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_993),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_952),
.A2(n_766),
.B1(n_804),
.B2(n_775),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_899),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_891),
.A2(n_804),
.B1(n_717),
.B2(n_733),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_835),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_850),
.B(n_663),
.Y(n_1079)
);

AO22x1_ASAP7_75t_L g1080 ( 
.A1(n_839),
.A2(n_439),
.B1(n_787),
.B2(n_277),
.Y(n_1080)
);

CKINVDCx8_ASAP7_75t_R g1081 ( 
.A(n_826),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_832),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_985),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_964),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_973),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_863),
.B(n_702),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_879),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_879),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_879),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_SL g1090 ( 
.A(n_900),
.B(n_625),
.C(n_815),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_840),
.B(n_689),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_826),
.B(n_702),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_938),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_870),
.B(n_663),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_852),
.B(n_905),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_883),
.B(n_663),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_973),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_949),
.Y(n_1098)
);

INVxp67_ASAP7_75t_SL g1099 ( 
.A(n_853),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_955),
.B(n_717),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_832),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_985),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_966),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_847),
.B(n_689),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_979),
.B(n_717),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_982),
.B(n_733),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_894),
.B(n_916),
.Y(n_1107)
);

BUFx4f_ASAP7_75t_SL g1108 ( 
.A(n_947),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_903),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_874),
.B(n_733),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_974),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_974),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_858),
.B(n_735),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_975),
.Y(n_1114)
);

AND2x6_ASAP7_75t_SL g1115 ( 
.A(n_956),
.B(n_348),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_951),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_942),
.Y(n_1117)
);

BUFx2_ASAP7_75t_SL g1118 ( 
.A(n_872),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_948),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_977),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_SL g1121 ( 
.A(n_869),
.B(n_286),
.C(n_278),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_826),
.B(n_702),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_961),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_868),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_950),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_866),
.B(n_735),
.Y(n_1126)
);

OA22x2_ASAP7_75t_L g1127 ( 
.A1(n_941),
.A2(n_937),
.B1(n_963),
.B2(n_920),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_963),
.B(n_735),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_SL g1129 ( 
.A(n_868),
.B(n_625),
.C(n_337),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_985),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_975),
.A2(n_777),
.B1(n_783),
.B2(n_779),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_939),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_853),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_855),
.B(n_761),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_944),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_946),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_855),
.B(n_761),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_924),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_927),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_898),
.B(n_761),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_845),
.B(n_783),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_930),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_970),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_845),
.B(n_792),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_947),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_976),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_907),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_975),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_958),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_980),
.B(n_772),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_936),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_975),
.Y(n_1152)
);

INVxp67_ASAP7_75t_SL g1153 ( 
.A(n_924),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_893),
.B(n_792),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_959),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_947),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_842),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_881),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_885),
.A2(n_795),
.B1(n_702),
.B2(n_671),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_915),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_983),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_825),
.B(n_335),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_836),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_981),
.Y(n_1164)
);

AO22x1_ASAP7_75t_L g1165 ( 
.A1(n_825),
.A2(n_287),
.B1(n_289),
.B2(n_288),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_987),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_887),
.B(n_675),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_896),
.B(n_795),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_963),
.B(n_666),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_963),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_836),
.B(n_867),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_965),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_873),
.B(n_666),
.Y(n_1173)
);

INVx3_ASAP7_75t_SL g1174 ( 
.A(n_880),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_906),
.B(n_671),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_917),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_857),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_984),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_919),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_880),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_925),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_965),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_965),
.B(n_689),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_878),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_901),
.B(n_676),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_972),
.Y(n_1186)
);

BUFx4f_ASAP7_75t_L g1187 ( 
.A(n_875),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_908),
.B(n_673),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_986),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_860),
.B(n_676),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_926),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_SL g1192 ( 
.A(n_933),
.B(n_298),
.C(n_293),
.Y(n_1192)
);

NOR2x1_ASAP7_75t_L g1193 ( 
.A(n_1040),
.B(n_923),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1147),
.A2(n_987),
.B(n_912),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1117),
.B(n_909),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1124),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1008),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1139),
.B(n_988),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1187),
.A2(n_931),
.B(n_922),
.C(n_943),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1132),
.A2(n_968),
.B(n_994),
.C(n_878),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1135),
.A2(n_1136),
.B(n_1151),
.C(n_1125),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1099),
.A2(n_931),
.B(n_922),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1058),
.A2(n_706),
.B(n_693),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1014),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1134),
.A2(n_996),
.B(n_990),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_1163),
.A2(n_999),
.B(n_918),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1142),
.B(n_921),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1164),
.B(n_876),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1058),
.B(n_965),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1067),
.B(n_886),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1037),
.B(n_928),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1119),
.B(n_1054),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1054),
.B(n_876),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1058),
.A2(n_706),
.B(n_693),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1058),
.A2(n_706),
.B(n_693),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1147),
.A2(n_910),
.B(n_902),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1147),
.A2(n_910),
.B(n_902),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1058),
.A2(n_871),
.B(n_861),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1163),
.A2(n_929),
.B(n_367),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1095),
.A2(n_871),
.B(n_861),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1008),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1076),
.B(n_1109),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1050),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1137),
.A2(n_997),
.B(n_934),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1047),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1151),
.B(n_886),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1160),
.B(n_889),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1187),
.A2(n_889),
.B(n_367),
.C(n_371),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1018),
.A2(n_934),
.B1(n_954),
.B2(n_932),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1176),
.B(n_673),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1102),
.A2(n_737),
.B(n_719),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1091),
.A2(n_1104),
.B(n_1172),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1171),
.A2(n_997),
.B(n_954),
.Y(n_1233)
);

OA22x2_ASAP7_75t_L g1234 ( 
.A1(n_1055),
.A2(n_772),
.B1(n_371),
.B2(n_393),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1001),
.A2(n_967),
.B(n_932),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1181),
.B(n_965),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1001),
.A2(n_1002),
.B(n_1079),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1008),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1015),
.A2(n_971),
.B(n_967),
.Y(n_1239)
);

INVx3_ASAP7_75t_SL g1240 ( 
.A(n_1029),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1190),
.A2(n_971),
.B(n_957),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1191),
.B(n_965),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1123),
.A2(n_989),
.B1(n_957),
.B2(n_430),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1190),
.A2(n_989),
.B(n_687),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1146),
.B(n_978),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1002),
.A2(n_1183),
.B(n_1104),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1032),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1015),
.A2(n_1184),
.A3(n_1157),
.B(n_1133),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1153),
.A2(n_409),
.B1(n_358),
.B2(n_373),
.Y(n_1249)
);

OA22x2_ASAP7_75t_L g1250 ( 
.A1(n_1004),
.A2(n_354),
.B1(n_393),
.B2(n_398),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1183),
.A2(n_687),
.B(n_677),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_SL g1252 ( 
.A1(n_1041),
.A2(n_398),
.B(n_354),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1027),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1035),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1133),
.A2(n_688),
.B(n_677),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_SL g1256 ( 
.A1(n_1041),
.A2(n_403),
.B(n_400),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1017),
.A2(n_390),
.B1(n_408),
.B2(n_410),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1149),
.B(n_965),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1155),
.B(n_978),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1091),
.A2(n_692),
.B(n_688),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1172),
.A2(n_694),
.B(n_692),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_SL g1262 ( 
.A1(n_1041),
.A2(n_403),
.B(n_400),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1027),
.B(n_411),
.Y(n_1263)
);

AND2x6_ASAP7_75t_SL g1264 ( 
.A(n_1162),
.B(n_407),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1185),
.A2(n_699),
.B(n_694),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1172),
.A2(n_780),
.B(n_758),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1143),
.B(n_978),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1182),
.A2(n_734),
.B(n_699),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1182),
.A2(n_744),
.B(n_734),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1040),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1162),
.B(n_520),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1185),
.A2(n_762),
.B(n_744),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1123),
.B(n_520),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1113),
.A2(n_774),
.B(n_762),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1182),
.A2(n_776),
.B(n_774),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1014),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1029),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1019),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1143),
.B(n_978),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1175),
.A2(n_781),
.B(n_776),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1008),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1188),
.A2(n_781),
.A3(n_796),
.B(n_802),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1090),
.B(n_524),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1031),
.A2(n_780),
.B(n_758),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1064),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1126),
.A2(n_953),
.B(n_802),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1019),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1005),
.B(n_978),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1116),
.A2(n_813),
.B(n_796),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1022),
.Y(n_1290)
);

AND3x1_ASAP7_75t_L g1291 ( 
.A(n_1062),
.B(n_412),
.C(n_407),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1031),
.A2(n_813),
.B(n_798),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1080),
.B(n_312),
.C(n_307),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1187),
.A2(n_428),
.B(n_412),
.C(n_414),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1141),
.A2(n_798),
.B(n_978),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1022),
.Y(n_1296)
);

INVx5_ASAP7_75t_L g1297 ( 
.A(n_1102),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1116),
.A2(n_798),
.B(n_616),
.Y(n_1298)
);

NOR3xp33_ASAP7_75t_L g1299 ( 
.A(n_1129),
.B(n_321),
.C(n_315),
.Y(n_1299)
);

NOR3xp33_ASAP7_75t_L g1300 ( 
.A(n_1165),
.B(n_325),
.C(n_322),
.Y(n_1300)
);

OAI21xp33_ASAP7_75t_L g1301 ( 
.A1(n_1059),
.A2(n_445),
.B(n_338),
.Y(n_1301)
);

O2A1O1Ixp5_ASAP7_75t_SL g1302 ( 
.A1(n_1000),
.A2(n_565),
.B(n_561),
.C(n_558),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1144),
.A2(n_978),
.B(n_616),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1010),
.Y(n_1304)
);

AOI221x1_ASAP7_75t_L g1305 ( 
.A1(n_1042),
.A2(n_547),
.B1(n_565),
.B2(n_556),
.C(n_555),
.Y(n_1305)
);

NOR2x1_ASAP7_75t_L g1306 ( 
.A(n_1044),
.B(n_414),
.Y(n_1306)
);

AOI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1127),
.A2(n_340),
.B(n_331),
.Y(n_1307)
);

AO21x2_ASAP7_75t_L g1308 ( 
.A1(n_1173),
.A2(n_529),
.B(n_524),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1011),
.A2(n_1127),
.B1(n_1138),
.B2(n_1024),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1120),
.B(n_719),
.Y(n_1310)
);

AND3x1_ASAP7_75t_L g1311 ( 
.A(n_1012),
.B(n_442),
.C(n_428),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1102),
.A2(n_780),
.B(n_758),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1120),
.B(n_719),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1102),
.A2(n_814),
.B(n_811),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1051),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1130),
.A2(n_814),
.B(n_811),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1072),
.B(n_719),
.Y(n_1317)
);

NOR2x1_ASAP7_75t_SL g1318 ( 
.A(n_1130),
.B(n_719),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1064),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1051),
.A2(n_444),
.A3(n_442),
.B(n_549),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1148),
.A2(n_616),
.B(n_615),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1179),
.B(n_737),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1130),
.A2(n_814),
.B(n_811),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1148),
.A2(n_631),
.B(n_615),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1059),
.A2(n_444),
.B(n_556),
.C(n_555),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1138),
.A2(n_737),
.B1(n_743),
.B2(n_429),
.Y(n_1326)
);

NAND2x1p5_ASAP7_75t_L g1327 ( 
.A(n_1050),
.B(n_737),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1003),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1179),
.B(n_737),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1130),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1026),
.A2(n_743),
.B1(n_425),
.B2(n_422),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1060),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1073),
.B(n_1056),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1026),
.B(n_529),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1003),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1148),
.A2(n_615),
.B(n_631),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1093),
.B(n_1107),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1152),
.A2(n_631),
.B(n_639),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1158),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1006),
.A2(n_539),
.A3(n_532),
.B(n_534),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1026),
.B(n_531),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1020),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1007),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1152),
.A2(n_639),
.B(n_642),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_SL g1345 ( 
.A(n_1150),
.B(n_365),
.C(n_364),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1050),
.A2(n_821),
.B(n_743),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1107),
.B(n_743),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1010),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1107),
.B(n_1167),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1038),
.A2(n_280),
.B1(n_558),
.B2(n_553),
.Y(n_1350)
);

NAND2x1_ASAP7_75t_L g1351 ( 
.A(n_1009),
.B(n_1071),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1044),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1167),
.B(n_743),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1066),
.Y(n_1354)
);

AOI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1013),
.A2(n_639),
.B(n_642),
.Y(n_1355)
);

AOI21xp33_ASAP7_75t_L g1356 ( 
.A1(n_1098),
.A2(n_346),
.B(n_345),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1152),
.A2(n_642),
.B(n_539),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1020),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1225),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1261),
.A2(n_1178),
.B(n_1161),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1343),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1252),
.A2(n_1077),
.B(n_1021),
.Y(n_1362)
);

AND2x6_ASAP7_75t_L g1363 ( 
.A(n_1223),
.B(n_1138),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1247),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1261),
.A2(n_1178),
.B(n_1161),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1204),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1268),
.A2(n_1189),
.B(n_1025),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1330),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1256),
.A2(n_1030),
.B(n_1016),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1257),
.A2(n_1121),
.B(n_1158),
.C(n_1174),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1204),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1303),
.A2(n_1110),
.B(n_1154),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1270),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1303),
.A2(n_1168),
.B(n_1039),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1276),
.Y(n_1375)
);

OAI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1301),
.A2(n_1180),
.B1(n_1174),
.B2(n_1069),
.C(n_1192),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1297),
.Y(n_1377)
);

OR2x6_ASAP7_75t_L g1378 ( 
.A(n_1231),
.B(n_1170),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1271),
.B(n_1086),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1297),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1268),
.A2(n_1189),
.B(n_1048),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1330),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1328),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1296),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1328),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1270),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1305),
.A2(n_1052),
.B(n_1034),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1203),
.A2(n_1083),
.B(n_1071),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1207),
.A2(n_1049),
.B1(n_1081),
.B2(n_1169),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1333),
.B(n_1068),
.Y(n_1390)
);

BUFx2_ASAP7_75t_SL g1391 ( 
.A(n_1352),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1211),
.A2(n_1049),
.B1(n_1081),
.B2(n_1169),
.Y(n_1392)
);

AND3x2_ASAP7_75t_L g1393 ( 
.A(n_1285),
.B(n_1170),
.C(n_1332),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1269),
.A2(n_1063),
.B(n_1061),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1225),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1300),
.B(n_1042),
.C(n_1092),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1269),
.A2(n_1070),
.B(n_1066),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1202),
.A2(n_1075),
.B(n_1078),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1315),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1208),
.A2(n_1046),
.B(n_1087),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1349),
.B(n_1092),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1208),
.A2(n_1046),
.B(n_1089),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1249),
.B(n_1186),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1278),
.Y(n_1404)
);

OAI222xp33_ASAP7_75t_L g1405 ( 
.A1(n_1250),
.A2(n_1122),
.B1(n_1092),
.B2(n_1186),
.C1(n_1086),
.C2(n_1103),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1275),
.A2(n_1085),
.B(n_1070),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1297),
.B(n_1138),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1195),
.B(n_1068),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1198),
.A2(n_1169),
.B1(n_1068),
.B2(n_1114),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1275),
.A2(n_1097),
.B(n_1085),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1295),
.A2(n_1112),
.B(n_1097),
.Y(n_1411)
);

NOR2x1_ASAP7_75t_SL g1412 ( 
.A(n_1297),
.B(n_1071),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_SL g1413 ( 
.A1(n_1262),
.A2(n_1159),
.B(n_1074),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1295),
.A2(n_1112),
.B(n_1111),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1199),
.A2(n_1038),
.B(n_1131),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1333),
.A2(n_1122),
.B1(n_1092),
.B2(n_1056),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1333),
.A2(n_1122),
.B1(n_1056),
.B2(n_1128),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1214),
.A2(n_1083),
.B(n_1009),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1278),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1232),
.A2(n_1201),
.B(n_1309),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1221),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1201),
.B(n_1043),
.Y(n_1422)
);

OR2x6_ASAP7_75t_L g1423 ( 
.A(n_1330),
.B(n_1122),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1286),
.A2(n_1128),
.B(n_1114),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1319),
.B(n_1118),
.Y(n_1425)
);

INVx4_ASAP7_75t_SL g1426 ( 
.A(n_1248),
.Y(n_1426)
);

NAND2xp33_ASAP7_75t_SL g1427 ( 
.A(n_1223),
.B(n_1150),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1237),
.A2(n_1128),
.B(n_1096),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1209),
.B(n_1083),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1287),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_SL g1431 ( 
.A1(n_1228),
.A2(n_1053),
.B(n_1088),
.C(n_1028),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1220),
.A2(n_1046),
.B(n_1043),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1246),
.A2(n_1028),
.B(n_1053),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1299),
.A2(n_1307),
.B1(n_1263),
.B2(n_1250),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1246),
.A2(n_1028),
.B(n_1053),
.Y(n_1435)
);

BUFx2_ASAP7_75t_R g1436 ( 
.A(n_1335),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1237),
.A2(n_1096),
.B(n_1094),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_SL g1438 ( 
.A(n_1283),
.B(n_1177),
.C(n_1156),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1357),
.A2(n_1088),
.B(n_1140),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1287),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1290),
.Y(n_1441)
);

CKINVDCx16_ASAP7_75t_R g1442 ( 
.A(n_1277),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1263),
.B(n_1177),
.Y(n_1443)
);

O2A1O1Ixp5_ASAP7_75t_L g1444 ( 
.A1(n_1227),
.A2(n_1043),
.B(n_1088),
.C(n_1009),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1290),
.Y(n_1445)
);

BUFx2_ASAP7_75t_R g1446 ( 
.A(n_1335),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1212),
.A2(n_1115),
.B1(n_1156),
.B2(n_1082),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1196),
.B(n_1084),
.Y(n_1448)
);

AOI22x1_ASAP7_75t_L g1449 ( 
.A1(n_1206),
.A2(n_1166),
.B1(n_1065),
.B2(n_1096),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_SL g1450 ( 
.A1(n_1241),
.A2(n_1140),
.B(n_1046),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1357),
.A2(n_1140),
.B(n_1046),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1321),
.A2(n_1140),
.B(n_1046),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1354),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1334),
.A2(n_1084),
.B1(n_1094),
.B2(n_1106),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1354),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1273),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1341),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1277),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1200),
.A2(n_1094),
.B(n_1100),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1222),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1240),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1352),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1358),
.A2(n_1108),
.B1(n_1082),
.B2(n_1145),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1196),
.B(n_1166),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1308),
.A2(n_1105),
.B(n_1100),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1321),
.A2(n_1140),
.B(n_532),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1282),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1209),
.B(n_1045),
.Y(n_1468)
);

AOI211x1_ASAP7_75t_L g1469 ( 
.A1(n_1337),
.A2(n_1356),
.B(n_1293),
.C(n_1213),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1324),
.A2(n_1140),
.B(n_531),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1308),
.A2(n_1100),
.B(n_1106),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1215),
.A2(n_1023),
.B(n_1010),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1253),
.B(n_1065),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1339),
.B(n_1045),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1253),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1351),
.B(n_1221),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1200),
.A2(n_1106),
.B(n_1105),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1336),
.A2(n_553),
.B(n_537),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1332),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1230),
.B(n_1065),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1240),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1340),
.Y(n_1482)
);

AOI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1355),
.A2(n_1105),
.B(n_537),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1226),
.B(n_1065),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1221),
.B(n_1045),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1342),
.B(n_1166),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1340),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1282),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1236),
.A2(n_1045),
.B1(n_1057),
.B2(n_1166),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1254),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1282),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1282),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1336),
.A2(n_561),
.B(n_538),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1338),
.A2(n_538),
.B(n_547),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1251),
.Y(n_1495)
);

AO31x2_ASAP7_75t_L g1496 ( 
.A1(n_1228),
.A2(n_1010),
.A3(n_1023),
.B(n_1033),
.Y(n_1496)
);

AO21x1_ASAP7_75t_L g1497 ( 
.A1(n_1229),
.A2(n_245),
.B(n_1023),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1345),
.A2(n_1306),
.B1(n_1193),
.B2(n_1311),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1210),
.B(n_1057),
.Y(n_1499)
);

AO21x1_ASAP7_75t_L g1500 ( 
.A1(n_1233),
.A2(n_1023),
.B(n_1033),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1350),
.B(n_1057),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1251),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1291),
.A2(n_1145),
.B1(n_1101),
.B2(n_441),
.C(n_440),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1210),
.A2(n_1057),
.B1(n_1036),
.B2(n_1033),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1264),
.B(n_1101),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1340),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1338),
.A2(n_1344),
.B(n_1194),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1340),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1320),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1320),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1350),
.B(n_1033),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1320),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1244),
.A2(n_1036),
.B(n_104),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1344),
.A2(n_1036),
.B(n_106),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1320),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1194),
.A2(n_1036),
.B(n_101),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1221),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1292),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1210),
.A2(n_342),
.B1(n_361),
.B2(n_362),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1260),
.A2(n_172),
.B(n_118),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1348),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_SL g1522 ( 
.A1(n_1218),
.A2(n_226),
.B(n_225),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1348),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1248),
.B(n_363),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1325),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1325),
.Y(n_1526)
);

CKINVDCx9p33_ASAP7_75t_R g1527 ( 
.A(n_1347),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1327),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1331),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1248),
.B(n_366),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1294),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1234),
.B(n_369),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1260),
.A2(n_171),
.B(n_130),
.Y(n_1533)
);

BUFx8_ASAP7_75t_SL g1534 ( 
.A(n_1304),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1294),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1242),
.A2(n_401),
.B1(n_377),
.B2(n_434),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1322),
.Y(n_1537)
);

AO31x2_ASAP7_75t_L g1538 ( 
.A1(n_1497),
.A2(n_1288),
.A3(n_1318),
.B(n_1353),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1386),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1457),
.B(n_1234),
.Y(n_1540)
);

NOR2x1_ASAP7_75t_SL g1541 ( 
.A(n_1378),
.B(n_1304),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1361),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1379),
.B(n_1248),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1529),
.A2(n_1243),
.B1(n_1259),
.B2(n_1245),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1366),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1529),
.A2(n_1258),
.B1(n_1329),
.B2(n_1267),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1375),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1403),
.A2(n_374),
.B1(n_378),
.B2(n_382),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1460),
.B(n_1317),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1456),
.B(n_1317),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1423),
.B(n_1238),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1460),
.B(n_1310),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1384),
.Y(n_1553)
);

OR2x2_ASAP7_75t_SL g1554 ( 
.A(n_1442),
.B(n_1304),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1408),
.A2(n_1279),
.B1(n_1313),
.B2(n_388),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1443),
.A2(n_1317),
.B1(n_404),
.B2(n_405),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1434),
.B(n_1304),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1498),
.A2(n_387),
.B1(n_394),
.B2(n_413),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1386),
.Y(n_1559)
);

INVxp33_ASAP7_75t_L g1560 ( 
.A(n_1448),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1385),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1486),
.B(n_1238),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1499),
.B(n_1197),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1496),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1519),
.A2(n_433),
.B1(n_418),
.B2(n_1219),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1496),
.Y(n_1566)
);

CKINVDCx11_ASAP7_75t_R g1567 ( 
.A(n_1461),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1425),
.A2(n_1326),
.B1(n_1238),
.B2(n_1327),
.Y(n_1568)
);

OAI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1376),
.A2(n_1298),
.B1(n_1272),
.B2(n_1265),
.C(n_1274),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1499),
.B(n_1197),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1399),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1377),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1464),
.B(n_1524),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1454),
.A2(n_1197),
.B1(n_1281),
.B2(n_1239),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1395),
.B(n_1197),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1531),
.A2(n_1239),
.B1(n_1289),
.B2(n_1255),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1419),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1524),
.B(n_1281),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1462),
.B(n_1281),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1479),
.B(n_1281),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1462),
.B(n_1224),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1521),
.B(n_1224),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_R g1583 ( 
.A(n_1393),
.B(n_1239),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1430),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1400),
.A2(n_1205),
.B(n_1302),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1389),
.A2(n_1346),
.B1(n_1280),
.B2(n_1284),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1377),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1479),
.B(n_1216),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1390),
.B(n_12),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1390),
.B(n_1292),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1383),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1392),
.A2(n_1216),
.B1(n_1217),
.B2(n_1235),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1390),
.B(n_14),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1396),
.A2(n_1217),
.B1(n_1235),
.B2(n_1280),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1383),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1371),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1417),
.A2(n_1280),
.B1(n_1266),
.B2(n_1314),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1532),
.A2(n_1323),
.B1(n_1316),
.B2(n_1312),
.C(n_20),
.Y(n_1598)
);

BUFx4_ASAP7_75t_R g1599 ( 
.A(n_1534),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1534),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1440),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_L g1602 ( 
.A(n_1469),
.B(n_14),
.C(n_15),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1537),
.B(n_15),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1364),
.B(n_17),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1423),
.B(n_99),
.Y(n_1605)
);

BUFx4f_ASAP7_75t_SL g1606 ( 
.A(n_1461),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1475),
.B(n_21),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1445),
.Y(n_1608)
);

OAI222xp33_ASAP7_75t_L g1609 ( 
.A1(n_1503),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.C1(n_31),
.C2(n_32),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1359),
.B(n_22),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1371),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1490),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1496),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1370),
.B(n_29),
.C(n_33),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1423),
.B(n_224),
.Y(n_1615)
);

BUFx12f_ASAP7_75t_L g1616 ( 
.A(n_1458),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1523),
.B(n_34),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1490),
.Y(n_1618)
);

NOR3xp33_ASAP7_75t_SL g1619 ( 
.A(n_1438),
.B(n_34),
.C(n_35),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1391),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1373),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1401),
.B(n_36),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1401),
.B(n_36),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1530),
.B(n_38),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1404),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1436),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1416),
.B(n_38),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1535),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_SL g1629 ( 
.A(n_1505),
.B(n_1385),
.C(n_1481),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1405),
.B(n_45),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1516),
.A2(n_222),
.B(n_221),
.Y(n_1631)
);

AO22x1_ASAP7_75t_SL g1632 ( 
.A1(n_1474),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_1632)
);

AO21x1_ASAP7_75t_L g1633 ( 
.A1(n_1422),
.A2(n_55),
.B(n_56),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1447),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1525),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1423),
.B(n_138),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_R g1637 ( 
.A(n_1415),
.B(n_218),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1404),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1441),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1441),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1453),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1473),
.B(n_60),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1536),
.B(n_64),
.Y(n_1643)
);

OAI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1526),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_1644)
);

CKINVDCx20_ASAP7_75t_R g1645 ( 
.A(n_1481),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1530),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1373),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1504),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1409),
.A2(n_79),
.B1(n_80),
.B2(n_85),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1455),
.Y(n_1650)
);

O2A1O1Ixp5_ASAP7_75t_L g1651 ( 
.A1(n_1497),
.A2(n_1422),
.B(n_1500),
.C(n_1432),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1474),
.B(n_85),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1501),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1474),
.B(n_158),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1458),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_SL g1656 ( 
.A1(n_1484),
.A2(n_87),
.B(n_90),
.C(n_91),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1467),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_SL g1658 ( 
.A(n_1377),
.B(n_90),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1509),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1527),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1517),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1467),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1488),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1510),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1480),
.B(n_92),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1517),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1512),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1459),
.A2(n_1477),
.B1(n_1511),
.B2(n_1378),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1515),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1377),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1482),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1446),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1488),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1377),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1463),
.B(n_93),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1378),
.B(n_168),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1427),
.Y(n_1677)
);

INVx8_ASAP7_75t_L g1678 ( 
.A(n_1517),
.Y(n_1678)
);

AO32x1_ASAP7_75t_L g1679 ( 
.A1(n_1487),
.A2(n_1506),
.A3(n_1508),
.B1(n_1491),
.B2(n_1492),
.Y(n_1679)
);

NAND2x1_ASAP7_75t_L g1680 ( 
.A(n_1421),
.B(n_821),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1407),
.B(n_93),
.Y(n_1681)
);

CKINVDCx16_ASAP7_75t_R g1682 ( 
.A(n_1427),
.Y(n_1682)
);

OAI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1378),
.A2(n_97),
.B1(n_142),
.B2(n_144),
.Y(n_1683)
);

INVx6_ASAP7_75t_L g1684 ( 
.A(n_1380),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1420),
.A2(n_97),
.B1(n_147),
.B2(n_149),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1489),
.A2(n_821),
.B1(n_785),
.B2(n_163),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1388),
.A2(n_785),
.B(n_154),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1380),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1420),
.B(n_153),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1491),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1413),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.C(n_194),
.Y(n_1691)
);

CKINVDCx8_ASAP7_75t_R g1692 ( 
.A(n_1380),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1363),
.A2(n_204),
.B1(n_206),
.B2(n_209),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1420),
.B(n_1368),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1368),
.B(n_785),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1492),
.Y(n_1696)
);

O2A1O1Ixp33_ASAP7_75t_SL g1697 ( 
.A1(n_1402),
.A2(n_785),
.B(n_1472),
.C(n_1418),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1407),
.B(n_1368),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1382),
.B(n_1426),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1380),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1449),
.A2(n_1468),
.B1(n_1485),
.B2(n_1429),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1413),
.A2(n_1513),
.B1(n_1362),
.B2(n_1522),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1382),
.B(n_1426),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1382),
.B(n_1426),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1369),
.B(n_1468),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1513),
.A2(n_1362),
.B1(n_1522),
.B2(n_1398),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1513),
.B(n_1431),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1380),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1421),
.B(n_1528),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1485),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1421),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1415),
.B(n_1471),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1517),
.A2(n_1468),
.B1(n_1387),
.B2(n_1429),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1429),
.A2(n_1517),
.B1(n_1528),
.B2(n_1476),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1363),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1363),
.B(n_1528),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1412),
.B(n_1363),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_SL g1718 ( 
.A(n_1369),
.B(n_1500),
.C(n_1450),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1476),
.A2(n_1428),
.B1(n_1437),
.B2(n_1483),
.Y(n_1719)
);

BUFx2_ASAP7_75t_SL g1720 ( 
.A(n_1363),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1363),
.A2(n_1398),
.B1(n_1471),
.B2(n_1465),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1476),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1465),
.B(n_1471),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1630),
.A2(n_1398),
.B1(n_1450),
.B2(n_1465),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1657),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1563),
.B(n_1516),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1558),
.A2(n_1431),
.B1(n_1444),
.B2(n_1495),
.C(n_1502),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1542),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1630),
.A2(n_1533),
.B1(n_1520),
.B2(n_1451),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1558),
.A2(n_1502),
.B1(n_1495),
.B2(n_1518),
.C(n_1496),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1570),
.B(n_1496),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1646),
.A2(n_1428),
.B1(n_1437),
.B2(n_1372),
.Y(n_1732)
);

AOI222xp33_ASAP7_75t_L g1733 ( 
.A1(n_1609),
.A2(n_1494),
.B1(n_1493),
.B2(n_1478),
.C1(n_1518),
.C2(n_1394),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1573),
.B(n_1622),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1646),
.A2(n_1428),
.B1(n_1437),
.B2(n_1372),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_SL g1736 ( 
.A1(n_1614),
.A2(n_1533),
.B1(n_1520),
.B2(n_1451),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1634),
.A2(n_1372),
.B1(n_1374),
.B2(n_1394),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1660),
.A2(n_1548),
.B1(n_1560),
.B2(n_1556),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1619),
.A2(n_1424),
.B(n_1494),
.C(n_1493),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1548),
.A2(n_1483),
.B1(n_1374),
.B2(n_1514),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1598),
.A2(n_1452),
.B(n_1439),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1567),
.Y(n_1742)
);

OAI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1634),
.A2(n_1374),
.B(n_1478),
.C(n_1414),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1635),
.A2(n_1367),
.B1(n_1381),
.B2(n_1360),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1649),
.A2(n_1514),
.B1(n_1470),
.B2(n_1466),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1629),
.A2(n_1433),
.B1(n_1435),
.B2(n_1367),
.Y(n_1746)
);

AO31x2_ASAP7_75t_L g1747 ( 
.A1(n_1719),
.A2(n_1507),
.A3(n_1414),
.B(n_1411),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1627),
.A2(n_1470),
.B1(n_1466),
.B2(n_1435),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1618),
.B(n_1433),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1635),
.A2(n_1381),
.B1(n_1411),
.B2(n_1360),
.C(n_1365),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1602),
.A2(n_1365),
.B1(n_1507),
.B2(n_1406),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1560),
.A2(n_1397),
.B1(n_1406),
.B2(n_1410),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1585),
.A2(n_1397),
.B(n_1410),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1628),
.A2(n_1619),
.B1(n_1643),
.B2(n_1685),
.C(n_1565),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1561),
.A2(n_1645),
.B1(n_1682),
.B2(n_1677),
.Y(n_1755)
);

OAI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1644),
.A2(n_1675),
.B1(n_1624),
.B2(n_1653),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1628),
.A2(n_1644),
.B1(n_1685),
.B2(n_1633),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1623),
.B(n_1543),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1676),
.A2(n_1648),
.B1(n_1615),
.B2(n_1605),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1642),
.B(n_1578),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1683),
.A2(n_1691),
.B1(n_1544),
.B2(n_1668),
.Y(n_1761)
);

AOI222xp33_ASAP7_75t_L g1762 ( 
.A1(n_1658),
.A2(n_1683),
.B1(n_1565),
.B2(n_1540),
.C1(n_1668),
.C2(n_1610),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1589),
.B(n_1593),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1720),
.B(n_1705),
.Y(n_1764)
);

BUFx12f_ASAP7_75t_L g1765 ( 
.A(n_1567),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1605),
.A2(n_1636),
.B1(n_1557),
.B2(n_1615),
.Y(n_1766)
);

AOI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1656),
.A2(n_1555),
.B1(n_1604),
.B2(n_1546),
.C(n_1607),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1605),
.A2(n_1636),
.B1(n_1606),
.B2(n_1681),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1562),
.B(n_1552),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1612),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1656),
.A2(n_1555),
.B1(n_1603),
.B2(n_1569),
.C(n_1550),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1547),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1553),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_SL g1774 ( 
.A1(n_1636),
.A2(n_1606),
.B1(n_1541),
.B2(n_1689),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1652),
.B(n_1549),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1693),
.A2(n_1702),
.B(n_1626),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1549),
.A2(n_1665),
.B1(n_1654),
.B2(n_1581),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1702),
.A2(n_1620),
.B1(n_1706),
.B2(n_1568),
.C(n_1687),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1620),
.A2(n_1554),
.B1(n_1618),
.B2(n_1692),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1654),
.A2(n_1581),
.B1(n_1616),
.B2(n_1617),
.Y(n_1780)
);

AOI21xp33_ASAP7_75t_SL g1781 ( 
.A1(n_1655),
.A2(n_1595),
.B(n_1591),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1632),
.A2(n_1706),
.B1(n_1721),
.B2(n_1707),
.C(n_1592),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1718),
.B(n_1637),
.C(n_1651),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1539),
.A2(n_1559),
.B1(n_1600),
.B2(n_1621),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1559),
.Y(n_1785)
);

INVx4_ASAP7_75t_L g1786 ( 
.A(n_1599),
.Y(n_1786)
);

AO221x2_ASAP7_75t_L g1787 ( 
.A1(n_1713),
.A2(n_1701),
.B1(n_1586),
.B2(n_1714),
.C(n_1574),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1590),
.A2(n_1551),
.B1(n_1647),
.B2(n_1600),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_SL g1789 ( 
.A1(n_1672),
.A2(n_1571),
.B1(n_1579),
.B2(n_1715),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1575),
.A2(n_1551),
.B1(n_1716),
.B2(n_1698),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1577),
.A2(n_1584),
.B1(n_1601),
.B2(n_1608),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1580),
.A2(n_1705),
.B1(n_1684),
.B2(n_1694),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1582),
.A2(n_1686),
.B1(n_1639),
.B2(n_1625),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1651),
.A2(n_1707),
.B(n_1718),
.C(n_1631),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1588),
.B(n_1650),
.Y(n_1795)
);

OAI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1637),
.A2(n_1583),
.B1(n_1705),
.B2(n_1722),
.Y(n_1796)
);

OAI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1594),
.A2(n_1597),
.B1(n_1583),
.B2(n_1576),
.C(n_1697),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1576),
.A2(n_1596),
.B1(n_1545),
.B2(n_1641),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1723),
.B(n_1722),
.C(n_1671),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1659),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1664),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1596),
.A2(n_1638),
.B1(n_1611),
.B2(n_1640),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1667),
.B(n_1669),
.Y(n_1803)
);

BUFx4f_ASAP7_75t_L g1804 ( 
.A(n_1678),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1684),
.A2(n_1700),
.B1(n_1710),
.B2(n_1708),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1709),
.B(n_1674),
.Y(n_1806)
);

OAI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1572),
.A2(n_1708),
.B1(n_1688),
.B2(n_1587),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1599),
.B(n_1674),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1662),
.B(n_1690),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1717),
.B(n_1699),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1712),
.A2(n_1717),
.B1(n_1670),
.B2(n_1678),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1661),
.B(n_1666),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1711),
.A2(n_1695),
.B(n_1704),
.Y(n_1813)
);

INVxp33_ASAP7_75t_L g1814 ( 
.A(n_1661),
.Y(n_1814)
);

AOI222xp33_ASAP7_75t_L g1815 ( 
.A1(n_1703),
.A2(n_1564),
.B1(n_1566),
.B2(n_1613),
.C1(n_1673),
.C2(n_1663),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1666),
.A2(n_1680),
.B1(n_1696),
.B2(n_1538),
.C(n_1678),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1666),
.A2(n_682),
.B1(n_608),
.B2(n_629),
.C(n_897),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1679),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1538),
.A2(n_1529),
.B1(n_1403),
.B2(n_1630),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1538),
.A2(n_1529),
.B1(n_897),
.B2(n_1403),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1679),
.Y(n_1821)
);

CKINVDCx11_ASAP7_75t_R g1822 ( 
.A(n_1538),
.Y(n_1822)
);

BUFx12f_ASAP7_75t_L g1823 ( 
.A(n_1679),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1660),
.A2(n_1529),
.B1(n_897),
.B2(n_1403),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1542),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1644),
.A2(n_643),
.B1(n_1529),
.B2(n_1630),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1618),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_SL g1829 ( 
.A(n_1720),
.B(n_1701),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1542),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1832)
);

AO21x2_ASAP7_75t_L g1833 ( 
.A1(n_1585),
.A2(n_1432),
.B(n_1450),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1558),
.A2(n_682),
.B1(n_608),
.B2(n_629),
.C(n_897),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1560),
.B(n_447),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1836)
);

BUFx4f_ASAP7_75t_L g1837 ( 
.A(n_1616),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1676),
.A2(n_1615),
.B(n_1605),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1644),
.A2(n_643),
.B1(n_1529),
.B2(n_1630),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1612),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1841)
);

A2O1A1Ixp33_ASAP7_75t_L g1842 ( 
.A1(n_1630),
.A2(n_897),
.B(n_839),
.C(n_700),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1644),
.A2(n_643),
.B1(n_1529),
.B2(n_1630),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1573),
.B(n_1622),
.Y(n_1845)
);

AO31x2_ASAP7_75t_L g1846 ( 
.A1(n_1719),
.A2(n_1497),
.A3(n_1707),
.B(n_1500),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1619),
.B(n_897),
.C(n_700),
.Y(n_1847)
);

CKINVDCx16_ASAP7_75t_R g1848 ( 
.A(n_1561),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1561),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1573),
.B(n_1622),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1573),
.B(n_1623),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1558),
.A2(n_897),
.B1(n_1529),
.B2(n_980),
.Y(n_1852)
);

A2O1A1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1630),
.A2(n_897),
.B(n_839),
.C(n_700),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1558),
.A2(n_897),
.B1(n_1529),
.B2(n_980),
.Y(n_1854)
);

AOI222xp33_ASAP7_75t_L g1855 ( 
.A1(n_1609),
.A2(n_1257),
.B1(n_682),
.B2(n_1403),
.C1(n_608),
.C2(n_643),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1697),
.A2(n_1422),
.B(n_1432),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1573),
.B(n_1623),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1859)
);

BUFx8_ASAP7_75t_SL g1860 ( 
.A(n_1561),
.Y(n_1860)
);

INVx11_ASAP7_75t_L g1861 ( 
.A(n_1616),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1548),
.A2(n_897),
.B1(n_700),
.B2(n_839),
.C(n_682),
.Y(n_1863)
);

OAI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1644),
.A2(n_643),
.B1(n_1529),
.B2(n_1630),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1660),
.A2(n_1529),
.B1(n_897),
.B2(n_1403),
.Y(n_1865)
);

OAI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1644),
.A2(n_643),
.B1(n_1529),
.B2(n_1630),
.Y(n_1866)
);

OAI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1644),
.A2(n_643),
.B1(n_1529),
.B2(n_1630),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_SL g1868 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_643),
.B2(n_897),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_SL g1869 ( 
.A1(n_1634),
.A2(n_1403),
.B1(n_1529),
.B2(n_897),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1614),
.A2(n_897),
.B(n_700),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1660),
.A2(n_1529),
.B1(n_897),
.B2(n_1403),
.Y(n_1872)
);

OAI211xp5_ASAP7_75t_SL g1873 ( 
.A1(n_1619),
.A2(n_682),
.B(n_1164),
.C(n_1062),
.Y(n_1873)
);

OAI21xp33_ASAP7_75t_L g1874 ( 
.A1(n_1548),
.A2(n_897),
.B(n_700),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1618),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1660),
.A2(n_1529),
.B1(n_897),
.B2(n_1403),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1630),
.A2(n_1529),
.B1(n_1403),
.B2(n_608),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1874),
.A2(n_1869),
.B1(n_1863),
.B2(n_1834),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1821),
.B(n_1846),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1800),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1818),
.B(n_1846),
.Y(n_1881)
);

NAND2x1_ASAP7_75t_L g1882 ( 
.A(n_1838),
.B(n_1764),
.Y(n_1882)
);

INVx2_ASAP7_75t_SL g1883 ( 
.A(n_1749),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1846),
.B(n_1833),
.Y(n_1884)
);

AO31x2_ASAP7_75t_L g1885 ( 
.A1(n_1794),
.A2(n_1752),
.A3(n_1740),
.B(n_1856),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1846),
.B(n_1833),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1725),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1801),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1747),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1758),
.B(n_1769),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1731),
.B(n_1787),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1747),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1787),
.B(n_1747),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1747),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1803),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1795),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1731),
.B(n_1787),
.Y(n_1897)
);

NAND2x1_ASAP7_75t_L g1898 ( 
.A(n_1783),
.B(n_1746),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1726),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1825),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1820),
.B(n_1842),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1830),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1799),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1809),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1724),
.B(n_1753),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1724),
.B(n_1753),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1810),
.B(n_1829),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1810),
.B(n_1741),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1728),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1819),
.B(n_1772),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1819),
.B(n_1773),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1822),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1792),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1823),
.B(n_1815),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1855),
.A2(n_1826),
.B1(n_1839),
.B2(n_1844),
.Y(n_1915)
);

INVxp67_ASAP7_75t_L g1916 ( 
.A(n_1785),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1791),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1750),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1732),
.B(n_1735),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1797),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1732),
.B(n_1735),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1791),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1816),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1748),
.B(n_1730),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1790),
.Y(n_1925)
);

BUFx3_ASAP7_75t_L g1926 ( 
.A(n_1875),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1729),
.B(n_1798),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1798),
.B(n_1744),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1806),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1812),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1778),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1813),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1811),
.B(n_1760),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1751),
.B(n_1737),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1737),
.B(n_1851),
.Y(n_1935)
);

OR2x6_ASAP7_75t_L g1936 ( 
.A(n_1743),
.B(n_1805),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1826),
.A2(n_1867),
.B1(n_1839),
.B2(n_1844),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1857),
.B(n_1727),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1770),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1802),
.B(n_1734),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1845),
.B(n_1850),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1796),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1733),
.B(n_1775),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1840),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1828),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1782),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1739),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1736),
.B(n_1745),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1761),
.B(n_1788),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1807),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1763),
.B(n_1757),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1757),
.B(n_1793),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1793),
.B(n_1789),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1784),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1766),
.B(n_1786),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1779),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1777),
.B(n_1774),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1786),
.B(n_1768),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1756),
.B(n_1776),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1771),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1814),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1853),
.B(n_1852),
.Y(n_1962)
);

OR2x6_ASAP7_75t_SL g1963 ( 
.A(n_1847),
.B(n_1742),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1756),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1762),
.B(n_1759),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1891),
.B(n_1780),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1939),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1891),
.B(n_1808),
.Y(n_1968)
);

NAND3xp33_ASAP7_75t_L g1969 ( 
.A(n_1878),
.B(n_1871),
.C(n_1831),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1891),
.B(n_1868),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1890),
.B(n_1767),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_R g1972 ( 
.A(n_1960),
.B(n_1849),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1897),
.B(n_1848),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1878),
.A2(n_1854),
.B(n_1877),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1880),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1881),
.B(n_1755),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1897),
.B(n_1835),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1962),
.A2(n_1901),
.B1(n_1864),
.B2(n_1866),
.C(n_1867),
.Y(n_1978)
);

AOI31xp33_ASAP7_75t_L g1979 ( 
.A1(n_1946),
.A2(n_1843),
.A3(n_1870),
.B(n_1862),
.Y(n_1979)
);

OA21x2_ASAP7_75t_L g1980 ( 
.A1(n_1889),
.A2(n_1754),
.B(n_1817),
.Y(n_1980)
);

OAI211xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1937),
.A2(n_1877),
.B(n_1858),
.C(n_1859),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1909),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1945),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1897),
.B(n_1899),
.Y(n_1984)
);

OAI31xp33_ASAP7_75t_L g1985 ( 
.A1(n_1962),
.A2(n_1864),
.A3(n_1866),
.B(n_1870),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1881),
.B(n_1893),
.Y(n_1986)
);

OAI211xp5_ASAP7_75t_L g1987 ( 
.A1(n_1901),
.A2(n_1841),
.B(n_1843),
.C(n_1862),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1915),
.A2(n_1937),
.B1(n_1946),
.B2(n_1831),
.Y(n_1988)
);

OAI221xp5_ASAP7_75t_SL g1989 ( 
.A1(n_1915),
.A2(n_1841),
.B1(n_1859),
.B2(n_1858),
.C(n_1836),
.Y(n_1989)
);

AOI21x1_ASAP7_75t_L g1990 ( 
.A1(n_1898),
.A2(n_1738),
.B(n_1876),
.Y(n_1990)
);

NAND4xp25_ASAP7_75t_L g1991 ( 
.A(n_1960),
.B(n_1836),
.C(n_1832),
.D(n_1827),
.Y(n_1991)
);

OA21x2_ASAP7_75t_L g1992 ( 
.A1(n_1889),
.A2(n_1892),
.B(n_1884),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1899),
.B(n_1832),
.Y(n_1993)
);

OAI21xp33_ASAP7_75t_SL g1994 ( 
.A1(n_1953),
.A2(n_1965),
.B(n_1959),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1880),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1888),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1881),
.B(n_1893),
.Y(n_1997)
);

CKINVDCx9p33_ASAP7_75t_R g1998 ( 
.A(n_1890),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1888),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1900),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1907),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1965),
.A2(n_1872),
.B1(n_1865),
.B2(n_1824),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1899),
.B(n_1935),
.Y(n_2003)
);

OAI21x1_ASAP7_75t_L g2004 ( 
.A1(n_1894),
.A2(n_1827),
.B(n_1804),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1907),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1945),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1899),
.B(n_1765),
.Y(n_2007)
);

AOI33xp33_ASAP7_75t_L g2008 ( 
.A1(n_1965),
.A2(n_1873),
.A3(n_1860),
.B1(n_1781),
.B2(n_1861),
.B3(n_1837),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1926),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_R g2010 ( 
.A(n_1929),
.B(n_1837),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_1898),
.B(n_1804),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1931),
.A2(n_1952),
.B1(n_1959),
.B2(n_1920),
.Y(n_2012)
);

AO21x2_ASAP7_75t_L g2013 ( 
.A1(n_1889),
.A2(n_1892),
.B(n_1947),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1939),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1887),
.Y(n_2015)
);

AOI32xp33_ASAP7_75t_L g2016 ( 
.A1(n_1952),
.A2(n_1931),
.A3(n_1920),
.B1(n_1959),
.B2(n_1964),
.Y(n_2016)
);

OAI33xp33_ASAP7_75t_L g2017 ( 
.A1(n_1964),
.A2(n_1947),
.A3(n_1922),
.B1(n_1917),
.B2(n_1893),
.B3(n_1910),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1963),
.B(n_1941),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1945),
.Y(n_2019)
);

OAI211xp5_ASAP7_75t_SL g2020 ( 
.A1(n_1931),
.A2(n_1920),
.B(n_1916),
.C(n_1917),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1931),
.A2(n_1952),
.B1(n_1920),
.B2(n_1957),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1899),
.B(n_1935),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1963),
.A2(n_1953),
.B1(n_1956),
.B2(n_1949),
.Y(n_2023)
);

OAI221xp5_ASAP7_75t_L g2024 ( 
.A1(n_1882),
.A2(n_1936),
.B1(n_1903),
.B2(n_1948),
.C(n_1932),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1935),
.B(n_1883),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1900),
.Y(n_2026)
);

AOI222xp33_ASAP7_75t_L g2027 ( 
.A1(n_1949),
.A2(n_1924),
.B1(n_1921),
.B2(n_1919),
.C1(n_1928),
.C2(n_1938),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_1945),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1902),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1940),
.B(n_1896),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1957),
.A2(n_1955),
.B1(n_1924),
.B2(n_1949),
.Y(n_2031)
);

OR2x6_ASAP7_75t_L g2032 ( 
.A(n_1882),
.B(n_1936),
.Y(n_2032)
);

NAND4xp25_ASAP7_75t_SL g2033 ( 
.A(n_1924),
.B(n_1948),
.C(n_1953),
.D(n_1934),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1902),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_1914),
.A2(n_1927),
.B1(n_1948),
.B2(n_1903),
.C(n_1934),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1955),
.B(n_1958),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1883),
.B(n_1904),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_1936),
.A2(n_1932),
.B1(n_1956),
.B2(n_1910),
.C(n_1911),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1957),
.A2(n_1955),
.B1(n_1958),
.B2(n_1938),
.Y(n_2039)
);

OAI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_1963),
.A2(n_1936),
.B1(n_1956),
.B2(n_1942),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1975),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1975),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2030),
.B(n_1879),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2015),
.B(n_1879),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1995),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_1992),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1986),
.B(n_1886),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2003),
.B(n_1905),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1995),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1967),
.B(n_1879),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2003),
.B(n_1905),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1986),
.B(n_1886),
.Y(n_2052)
);

NAND2xp33_ASAP7_75t_SL g2053 ( 
.A(n_1972),
.B(n_1912),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2022),
.B(n_1906),
.Y(n_2054)
);

AND2x4_ASAP7_75t_SL g2055 ( 
.A(n_2032),
.B(n_1907),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2025),
.B(n_1906),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_2013),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_2009),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2025),
.B(n_1906),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_2009),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1984),
.B(n_2001),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1992),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_2007),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1984),
.B(n_1908),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2014),
.B(n_1896),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1996),
.B(n_1895),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1992),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1996),
.Y(n_2068)
);

AND2x2_ASAP7_75t_SL g2069 ( 
.A(n_1980),
.B(n_1912),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_1997),
.B(n_1886),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1999),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_2013),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1999),
.B(n_1895),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2000),
.B(n_1918),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1992),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2000),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2013),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2026),
.Y(n_2078)
);

BUFx8_ASAP7_75t_L g2079 ( 
.A(n_1987),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2026),
.B(n_1918),
.Y(n_2080)
);

NOR3xp33_ASAP7_75t_SL g2081 ( 
.A(n_1969),
.B(n_1911),
.C(n_1950),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_1976),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1971),
.B(n_1941),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2001),
.B(n_1908),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_L g2085 ( 
.A(n_1978),
.B(n_1938),
.C(n_1922),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2005),
.B(n_1908),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2029),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2005),
.B(n_1908),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2029),
.B(n_2034),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2037),
.B(n_1976),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2034),
.B(n_1918),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_1969),
.A2(n_1955),
.B1(n_1934),
.B2(n_1927),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1982),
.B(n_1918),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1973),
.B(n_1930),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_2083),
.B(n_2007),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_2085),
.B(n_1977),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2041),
.Y(n_2097)
);

INVxp67_ASAP7_75t_SL g2098 ( 
.A(n_2074),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2041),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2042),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_L g2101 ( 
.A(n_2085),
.B(n_1977),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2082),
.B(n_2035),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2042),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2082),
.B(n_1885),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2063),
.B(n_2018),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2090),
.B(n_1885),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2065),
.B(n_1993),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2090),
.B(n_1885),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2045),
.Y(n_2109)
);

NAND2x1p5_ASAP7_75t_L g2110 ( 
.A(n_2069),
.B(n_2011),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2056),
.B(n_1973),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2065),
.B(n_2092),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2047),
.B(n_1885),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2045),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2049),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2056),
.B(n_1968),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2049),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2068),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2047),
.B(n_1885),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2068),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2071),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2071),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2076),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2056),
.B(n_1968),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2046),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2059),
.B(n_2032),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2052),
.B(n_1885),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_2046),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2076),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2078),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2078),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2052),
.B(n_1885),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_2058),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2046),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2046),
.Y(n_2135)
);

NAND2x1p5_ASAP7_75t_L g2136 ( 
.A(n_2069),
.B(n_2011),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_SL g2137 ( 
.A(n_2069),
.B(n_2024),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2074),
.B(n_1993),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2059),
.B(n_2061),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2087),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2087),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2059),
.B(n_2032),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2089),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_2080),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2089),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2066),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2066),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2061),
.B(n_2032),
.Y(n_2148)
);

NOR2x1_ASAP7_75t_L g2149 ( 
.A(n_2063),
.B(n_2020),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2080),
.B(n_1944),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2139),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2104),
.B(n_2070),
.Y(n_2152)
);

NAND2xp33_ASAP7_75t_R g2153 ( 
.A(n_2102),
.B(n_2081),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2104),
.B(n_2070),
.Y(n_2154)
);

CKINVDCx16_ASAP7_75t_R g2155 ( 
.A(n_2137),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2106),
.B(n_2091),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2103),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2096),
.B(n_2027),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2103),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2101),
.B(n_2112),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2139),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2109),
.Y(n_2162)
);

AND2x4_ASAP7_75t_SL g2163 ( 
.A(n_2148),
.B(n_2081),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2126),
.B(n_2064),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2109),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2126),
.B(n_2142),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2142),
.B(n_2064),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2148),
.B(n_2061),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2149),
.B(n_1994),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_2111),
.B(n_2055),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2114),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2125),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_SL g2173 ( 
.A(n_2110),
.B(n_1985),
.C(n_2023),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_2146),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2111),
.B(n_2116),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2114),
.Y(n_2176)
);

INVxp67_ASAP7_75t_L g2177 ( 
.A(n_2105),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2150),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2107),
.B(n_1994),
.Y(n_2179)
);

NAND4xp25_ASAP7_75t_L g2180 ( 
.A(n_2106),
.B(n_1985),
.C(n_2002),
.D(n_1974),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_2133),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2117),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2138),
.B(n_1970),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_SL g2184 ( 
.A(n_2110),
.B(n_2038),
.Y(n_2184)
);

INVx4_ASAP7_75t_L g2185 ( 
.A(n_2133),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2117),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2095),
.B(n_1970),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2116),
.B(n_2048),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2098),
.B(n_2031),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2108),
.B(n_2091),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2118),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2110),
.B(n_2063),
.Y(n_2192)
);

INVx2_ASAP7_75t_SL g2193 ( 
.A(n_2136),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2108),
.B(n_2050),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2124),
.B(n_2016),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2118),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2124),
.B(n_2048),
.Y(n_2197)
);

AOI22xp33_ASAP7_75t_L g2198 ( 
.A1(n_2136),
.A2(n_2079),
.B1(n_1981),
.B2(n_2033),
.Y(n_2198)
);

NOR2x1_ASAP7_75t_L g2199 ( 
.A(n_2097),
.B(n_2040),
.Y(n_2199)
);

NAND3xp33_ASAP7_75t_SL g2200 ( 
.A(n_2136),
.B(n_2016),
.C(n_2053),
.Y(n_2200)
);

NOR4xp25_ASAP7_75t_SL g2201 ( 
.A(n_2123),
.B(n_2010),
.C(n_1998),
.D(n_2036),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2125),
.Y(n_2202)
);

OR2x6_ASAP7_75t_L g2203 ( 
.A(n_2113),
.B(n_1936),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2144),
.B(n_2048),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2147),
.B(n_2043),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2181),
.B(n_2185),
.Y(n_2206)
);

OAI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_2155),
.A2(n_1990),
.B1(n_1979),
.B2(n_1980),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2166),
.B(n_2084),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2162),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2162),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2166),
.B(n_2084),
.Y(n_2211)
);

OAI22xp33_ASAP7_75t_L g2212 ( 
.A1(n_2184),
.A2(n_1990),
.B1(n_1980),
.B2(n_1912),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2170),
.Y(n_2213)
);

OAI21xp33_ASAP7_75t_L g2214 ( 
.A1(n_2169),
.A2(n_2160),
.B(n_2180),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2189),
.B(n_2113),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2173),
.A2(n_2079),
.B1(n_1991),
.B2(n_1980),
.Y(n_2216)
);

AOI211xp5_ASAP7_75t_L g2217 ( 
.A1(n_2169),
.A2(n_1989),
.B(n_1988),
.C(n_2127),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2165),
.Y(n_2218)
);

AOI32xp33_ASAP7_75t_L g2219 ( 
.A1(n_2163),
.A2(n_2021),
.A3(n_1966),
.B1(n_1914),
.B2(n_2012),
.Y(n_2219)
);

OAI322xp33_ASAP7_75t_L g2220 ( 
.A1(n_2153),
.A2(n_2158),
.A3(n_2002),
.B1(n_2177),
.B2(n_2119),
.C1(n_2127),
.C2(n_2132),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2174),
.B(n_2143),
.Y(n_2221)
);

AOI32xp33_ASAP7_75t_L g2222 ( 
.A1(n_2163),
.A2(n_1966),
.A3(n_1914),
.B1(n_2039),
.B2(n_1927),
.Y(n_2222)
);

AOI21xp33_ASAP7_75t_L g2223 ( 
.A1(n_2199),
.A2(n_2079),
.B(n_2119),
.Y(n_2223)
);

AND2x4_ASAP7_75t_L g2224 ( 
.A(n_2181),
.B(n_2055),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2165),
.Y(n_2225)
);

INVxp67_ASAP7_75t_L g2226 ( 
.A(n_2200),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2157),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2159),
.Y(n_2228)
);

INVx1_ASAP7_75t_SL g2229 ( 
.A(n_2185),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2187),
.B(n_2079),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2185),
.B(n_2143),
.Y(n_2231)
);

NOR2xp67_ASAP7_75t_L g2232 ( 
.A(n_2193),
.B(n_2145),
.Y(n_2232)
);

OAI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_2195),
.A2(n_1912),
.B1(n_1936),
.B2(n_1913),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2198),
.A2(n_2201),
.B1(n_2179),
.B2(n_1912),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2193),
.Y(n_2235)
);

OR2x6_ASAP7_75t_L g2236 ( 
.A(n_2192),
.B(n_2170),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2183),
.B(n_2145),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2178),
.B(n_2051),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2175),
.B(n_2051),
.Y(n_2239)
);

AOI32xp33_ASAP7_75t_L g2240 ( 
.A1(n_2168),
.A2(n_2055),
.A3(n_2132),
.B1(n_2086),
.B2(n_2088),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2170),
.B(n_1944),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2168),
.B(n_2086),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2171),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2175),
.Y(n_2244)
);

INVxp67_ASAP7_75t_L g2245 ( 
.A(n_2203),
.Y(n_2245)
);

AOI211xp5_ASAP7_75t_L g2246 ( 
.A1(n_2176),
.A2(n_2017),
.B(n_1921),
.C(n_1919),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_2203),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_L g2248 ( 
.A(n_2164),
.B(n_1941),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2209),
.Y(n_2249)
);

AOI31xp33_ASAP7_75t_L g2250 ( 
.A1(n_2226),
.A2(n_2161),
.A3(n_2151),
.B(n_1958),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2210),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2218),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2214),
.A2(n_1958),
.B(n_1955),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2225),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2217),
.B(n_2151),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2206),
.Y(n_2256)
);

OR2x2_ASAP7_75t_L g2257 ( 
.A(n_2244),
.B(n_2161),
.Y(n_2257)
);

O2A1O1Ixp33_ASAP7_75t_L g2258 ( 
.A1(n_2234),
.A2(n_2203),
.B(n_2182),
.C(n_2186),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2227),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2228),
.Y(n_2260)
);

INVxp67_ASAP7_75t_L g2261 ( 
.A(n_2206),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2243),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2229),
.B(n_2216),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2231),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2221),
.Y(n_2265)
);

OAI21xp33_ASAP7_75t_L g2266 ( 
.A1(n_2219),
.A2(n_2203),
.B(n_2194),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2215),
.B(n_2191),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2221),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2229),
.Y(n_2269)
);

OAI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2234),
.A2(n_2196),
.B(n_2004),
.Y(n_2270)
);

OAI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2246),
.A2(n_1912),
.B1(n_2164),
.B2(n_2167),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2235),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2235),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2220),
.A2(n_2205),
.B(n_2093),
.Y(n_2274)
);

NOR4xp75_ASAP7_75t_L g2275 ( 
.A(n_2230),
.B(n_2204),
.C(n_2197),
.D(n_2188),
.Y(n_2275)
);

OAI21xp5_ASAP7_75t_SL g2276 ( 
.A1(n_2222),
.A2(n_1958),
.B(n_1951),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_SL g2277 ( 
.A1(n_2207),
.A2(n_1912),
.B1(n_1913),
.B2(n_1925),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2224),
.B(n_2167),
.Y(n_2278)
);

OR2x6_ASAP7_75t_L g2279 ( 
.A(n_2269),
.B(n_2236),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2278),
.B(n_2236),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2249),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2278),
.B(n_2236),
.Y(n_2282)
);

XOR2x2_ASAP7_75t_L g2283 ( 
.A(n_2275),
.B(n_2263),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2251),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2261),
.B(n_2241),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2256),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2277),
.A2(n_2212),
.B1(n_2233),
.B2(n_2213),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2252),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2254),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_2256),
.Y(n_2290)
);

NAND2xp33_ASAP7_75t_R g2291 ( 
.A(n_2270),
.B(n_2224),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2272),
.B(n_2273),
.Y(n_2292)
);

NOR2xp67_ASAP7_75t_L g2293 ( 
.A(n_2261),
.B(n_2232),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2259),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2260),
.Y(n_2295)
);

INVxp67_ASAP7_75t_SL g2296 ( 
.A(n_2258),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2262),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2257),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2255),
.B(n_2264),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2257),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2267),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2267),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2286),
.Y(n_2303)
);

NOR4xp25_ASAP7_75t_L g2304 ( 
.A(n_2299),
.B(n_2266),
.C(n_2265),
.D(n_2268),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_SL g2305 ( 
.A(n_2280),
.B(n_2223),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2290),
.B(n_2253),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_2293),
.B(n_2277),
.Y(n_2307)
);

OAI221xp5_ASAP7_75t_L g2308 ( 
.A1(n_2296),
.A2(n_2283),
.B1(n_2276),
.B2(n_2291),
.C(n_2287),
.Y(n_2308)
);

INVx1_ASAP7_75t_SL g2309 ( 
.A(n_2280),
.Y(n_2309)
);

NAND4xp25_ASAP7_75t_SL g2310 ( 
.A(n_2282),
.B(n_2274),
.C(n_2223),
.D(n_2240),
.Y(n_2310)
);

NAND4xp25_ASAP7_75t_L g2311 ( 
.A(n_2285),
.B(n_2271),
.C(n_2245),
.D(n_2247),
.Y(n_2311)
);

OAI221xp5_ASAP7_75t_L g2312 ( 
.A1(n_2283),
.A2(n_2250),
.B1(n_2237),
.B2(n_2238),
.C(n_2239),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2290),
.Y(n_2313)
);

AOI21xp33_ASAP7_75t_SL g2314 ( 
.A1(n_2292),
.A2(n_2211),
.B(n_2208),
.Y(n_2314)
);

NOR3xp33_ASAP7_75t_L g2315 ( 
.A(n_2292),
.B(n_2008),
.C(n_2172),
.Y(n_2315)
);

NOR3xp33_ASAP7_75t_SL g2316 ( 
.A(n_2291),
.B(n_2248),
.C(n_2050),
.Y(n_2316)
);

OAI211xp5_ASAP7_75t_SL g2317 ( 
.A1(n_2294),
.A2(n_2172),
.B(n_2202),
.C(n_2194),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2303),
.Y(n_2318)
);

AOI21xp33_ASAP7_75t_L g2319 ( 
.A1(n_2308),
.A2(n_2279),
.B(n_2298),
.Y(n_2319)
);

OAI211xp5_ASAP7_75t_L g2320 ( 
.A1(n_2304),
.A2(n_2286),
.B(n_2282),
.C(n_2300),
.Y(n_2320)
);

OAI221xp5_ASAP7_75t_SL g2321 ( 
.A1(n_2312),
.A2(n_2279),
.B1(n_2301),
.B2(n_2302),
.C(n_2295),
.Y(n_2321)
);

AO22x2_ASAP7_75t_L g2322 ( 
.A1(n_2309),
.A2(n_2289),
.B1(n_2288),
.B2(n_2284),
.Y(n_2322)
);

NAND4xp25_ASAP7_75t_L g2323 ( 
.A(n_2305),
.B(n_2297),
.C(n_2281),
.D(n_2279),
.Y(n_2323)
);

OAI321xp33_ASAP7_75t_L g2324 ( 
.A1(n_2307),
.A2(n_2279),
.A3(n_2152),
.B1(n_2154),
.B2(n_2242),
.C(n_2190),
.Y(n_2324)
);

NAND3xp33_ASAP7_75t_SL g2325 ( 
.A(n_2316),
.B(n_2154),
.C(n_2152),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2313),
.B(n_2188),
.Y(n_2326)
);

OAI211xp5_ASAP7_75t_L g2327 ( 
.A1(n_2311),
.A2(n_2202),
.B(n_2190),
.C(n_2156),
.Y(n_2327)
);

AOI221xp5_ASAP7_75t_L g2328 ( 
.A1(n_2310),
.A2(n_2204),
.B1(n_2057),
.B2(n_2072),
.C(n_2134),
.Y(n_2328)
);

NOR4xp75_ASAP7_75t_L g2329 ( 
.A(n_2306),
.B(n_2128),
.C(n_2197),
.D(n_2044),
.Y(n_2329)
);

AOI222xp33_ASAP7_75t_L g2330 ( 
.A1(n_2317),
.A2(n_2072),
.B1(n_2057),
.B2(n_1951),
.C1(n_1921),
.C2(n_1919),
.Y(n_2330)
);

BUFx2_ASAP7_75t_L g2331 ( 
.A(n_2322),
.Y(n_2331)
);

AOI221xp5_ASAP7_75t_L g2332 ( 
.A1(n_2321),
.A2(n_2315),
.B1(n_2314),
.B2(n_2317),
.C(n_2128),
.Y(n_2332)
);

OAI21xp33_ASAP7_75t_SL g2333 ( 
.A1(n_2323),
.A2(n_2156),
.B(n_2128),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2326),
.B(n_2094),
.Y(n_2334)
);

NOR2x1p5_ASAP7_75t_L g2335 ( 
.A(n_2318),
.B(n_2058),
.Y(n_2335)
);

INVx1_ASAP7_75t_SL g2336 ( 
.A(n_2319),
.Y(n_2336)
);

OAI32xp33_ASAP7_75t_L g2337 ( 
.A1(n_2324),
.A2(n_2135),
.A3(n_2134),
.B1(n_2062),
.B2(n_2067),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2320),
.Y(n_2338)
);

NAND2xp33_ASAP7_75t_R g2339 ( 
.A(n_2329),
.B(n_1907),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_2328),
.Y(n_2340)
);

AOI222xp33_ASAP7_75t_L g2341 ( 
.A1(n_2325),
.A2(n_1951),
.B1(n_2135),
.B2(n_2067),
.C1(n_2075),
.C2(n_2062),
.Y(n_2341)
);

NAND4xp75_ASAP7_75t_L g2342 ( 
.A(n_2338),
.B(n_2327),
.C(n_2330),
.D(n_2088),
.Y(n_2342)
);

AOI221xp5_ASAP7_75t_L g2343 ( 
.A1(n_2331),
.A2(n_1916),
.B1(n_2067),
.B2(n_2062),
.C(n_2075),
.Y(n_2343)
);

NAND2xp33_ASAP7_75t_R g2344 ( 
.A(n_2334),
.B(n_1907),
.Y(n_2344)
);

OA21x2_ASAP7_75t_L g2345 ( 
.A1(n_2336),
.A2(n_2075),
.B(n_2123),
.Y(n_2345)
);

OAI211xp5_ASAP7_75t_SL g2346 ( 
.A1(n_2336),
.A2(n_2093),
.B(n_2044),
.C(n_1961),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2340),
.B(n_2332),
.Y(n_2347)
);

NOR4xp75_ASAP7_75t_SL g2348 ( 
.A(n_2333),
.B(n_2043),
.C(n_2073),
.D(n_2060),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2335),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_SL g2350 ( 
.A(n_2341),
.B(n_2028),
.C(n_1983),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2342),
.A2(n_2347),
.B1(n_2350),
.B2(n_2339),
.Y(n_2351)
);

HB1xp67_ASAP7_75t_L g2352 ( 
.A(n_2345),
.Y(n_2352)
);

NAND5xp2_ASAP7_75t_L g2353 ( 
.A(n_2349),
.B(n_2337),
.C(n_1942),
.D(n_1943),
.E(n_1933),
.Y(n_2353)
);

NOR5xp2_ASAP7_75t_L g2354 ( 
.A(n_2346),
.B(n_2141),
.C(n_2140),
.D(n_2131),
.E(n_2130),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2345),
.B(n_2099),
.Y(n_2355)
);

NAND3xp33_ASAP7_75t_SL g2356 ( 
.A(n_2343),
.B(n_1956),
.C(n_2019),
.Y(n_2356)
);

NOR2x1_ASAP7_75t_L g2357 ( 
.A(n_2348),
.B(n_2058),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2352),
.Y(n_2358)
);

NAND4xp25_ASAP7_75t_L g2359 ( 
.A(n_2351),
.B(n_2344),
.C(n_2060),
.D(n_1943),
.Y(n_2359)
);

NAND4xp25_ASAP7_75t_SL g2360 ( 
.A(n_2357),
.B(n_2094),
.C(n_2006),
.D(n_1923),
.Y(n_2360)
);

NAND3xp33_ASAP7_75t_L g2361 ( 
.A(n_2355),
.B(n_2060),
.C(n_1912),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2358),
.Y(n_2362)
);

INVxp67_ASAP7_75t_L g2363 ( 
.A(n_2359),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2362),
.B(n_2363),
.Y(n_2364)
);

BUFx2_ASAP7_75t_L g2365 ( 
.A(n_2364),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_R g2366 ( 
.A1(n_2364),
.A2(n_2360),
.B1(n_2361),
.B2(n_2356),
.Y(n_2366)
);

AOI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2365),
.A2(n_2353),
.B1(n_2354),
.B2(n_2129),
.Y(n_2367)
);

OAI21xp5_ASAP7_75t_SL g2368 ( 
.A1(n_2366),
.A2(n_1954),
.B(n_2121),
.Y(n_2368)
);

AOI21x1_ASAP7_75t_L g2369 ( 
.A1(n_2368),
.A2(n_2120),
.B(n_2115),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2367),
.Y(n_2370)
);

AOI222xp33_ASAP7_75t_L g2371 ( 
.A1(n_2370),
.A2(n_2122),
.B1(n_2100),
.B2(n_2077),
.C1(n_2051),
.C2(n_2054),
.Y(n_2371)
);

OAI221xp5_ASAP7_75t_R g2372 ( 
.A1(n_2371),
.A2(n_2369),
.B1(n_2077),
.B2(n_2004),
.C(n_2073),
.Y(n_2372)
);

AOI211xp5_ASAP7_75t_L g2373 ( 
.A1(n_2372),
.A2(n_1954),
.B(n_2077),
.C(n_1925),
.Y(n_2373)
);


endmodule