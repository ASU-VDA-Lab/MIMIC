module fake_netlist_5_255_n_770 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_770);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_770;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_629;
wire n_590;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_699;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_647;
wire n_710;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_38),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_79),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_22),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_47),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_46),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_21),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_61),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_122),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_2),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_33),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_111),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_5),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_10),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_48),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_37),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_35),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_90),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_50),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_80),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_42),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_68),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_4),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_149),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_27),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_59),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_23),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_137),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_118),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_70),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_85),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_108),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_18),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_40),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_100),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_153),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_0),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

CKINVDCx6p67_ASAP7_75t_R g215 ( 
.A(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_0),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_24),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_1),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_2),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_3),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_174),
.Y(n_223)
);

AOI22x1_ASAP7_75t_SL g224 ( 
.A1(n_177),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_161),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_156),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_178),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

CKINVDCx6p67_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_25),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_26),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_6),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_9),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_157),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_156),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_165),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_180),
.A2(n_11),
.B(n_12),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_189),
.A2(n_13),
.B(n_14),
.Y(n_251)
);

BUFx8_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_176),
.B(n_187),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_157),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_210),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_192),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

BUFx6f_ASAP7_75t_SL g261 ( 
.A(n_218),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_196),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_158),
.C(n_162),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_202),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_236),
.B(n_210),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_158),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_236),
.B(n_162),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_221),
.B(n_185),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_223),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_214),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_214),
.B(n_207),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_214),
.B(n_219),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_242),
.B(n_185),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_209),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_208),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_231),
.B(n_208),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_223),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_28),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_216),
.B(n_168),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_240),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_269),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_256),
.A2(n_235),
.B1(n_215),
.B2(n_241),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_217),
.Y(n_307)
);

O2A1O1Ixp5_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_238),
.B(n_222),
.C(n_248),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_217),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_217),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_256),
.A2(n_238),
.B1(n_250),
.B2(n_212),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_226),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_260),
.B(n_217),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_267),
.B(n_246),
.C(n_230),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_267),
.A2(n_238),
.B1(n_250),
.B2(n_212),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_215),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_226),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_260),
.B(n_217),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_241),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_279),
.B(n_225),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_265),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_296),
.B(n_225),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_264),
.B(n_248),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_235),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_250),
.B1(n_212),
.B2(n_251),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_227),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_276),
.B(n_225),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_259),
.B(n_244),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_290),
.A2(n_261),
.B1(n_302),
.B2(n_260),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_258),
.B(n_225),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_297),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

NOR2x1p5_ASAP7_75t_L g339 ( 
.A(n_262),
.B(n_232),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_240),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_259),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_263),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_274),
.B(n_225),
.Y(n_345)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_261),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_274),
.B(n_172),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_263),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_286),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_268),
.B(n_240),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_278),
.B(n_173),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_272),
.B(n_182),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_278),
.B(n_184),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_268),
.B(n_240),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_270),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_293),
.A2(n_237),
.B1(n_239),
.B2(n_186),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_261),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_271),
.B(n_240),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_275),
.B(n_234),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_272),
.B(n_188),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_278),
.B(n_194),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_275),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_272),
.B(n_195),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_302),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_282),
.B(n_252),
.Y(n_368)
);

O2A1O1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_305),
.A2(n_324),
.B(n_320),
.C(n_358),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_308),
.A2(n_251),
.B(n_272),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_228),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_228),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_272),
.B(n_277),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_322),
.A2(n_337),
.B(n_319),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_312),
.A2(n_277),
.B(n_280),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_314),
.A2(n_280),
.B(n_291),
.Y(n_378)
);

AO32x1_ASAP7_75t_L g379 ( 
.A1(n_323),
.A2(n_298),
.A3(n_292),
.B1(n_291),
.B2(n_234),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_294),
.Y(n_380)
);

BUFx4f_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_332),
.B(n_294),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_345),
.A2(n_292),
.B(n_298),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_335),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_283),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_313),
.B(n_283),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_330),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_313),
.A2(n_318),
.B1(n_306),
.B2(n_347),
.Y(n_388)
);

AOI21x1_ASAP7_75t_L g389 ( 
.A1(n_351),
.A2(n_289),
.B(n_288),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_318),
.B(n_327),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_284),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_304),
.A2(n_340),
.B(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_284),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_355),
.A2(n_361),
.B(n_309),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_352),
.A2(n_289),
.B(n_288),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_333),
.B(n_285),
.Y(n_397)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_355),
.A2(n_285),
.B(n_213),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_354),
.A2(n_213),
.B(n_252),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_361),
.A2(n_252),
.B(n_87),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_307),
.A2(n_86),
.B(n_155),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_367),
.B(n_224),
.Y(n_402)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_315),
.B(n_224),
.C(n_84),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_367),
.B(n_13),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_309),
.A2(n_89),
.B(n_152),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_339),
.A2(n_83),
.B1(n_147),
.B2(n_146),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_321),
.B(n_15),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_311),
.A2(n_82),
.B(n_145),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_338),
.B(n_341),
.Y(n_409)
);

NAND2x1p5_ASAP7_75t_L g410 ( 
.A(n_342),
.B(n_29),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_346),
.Y(n_411)
);

O2A1O1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_362),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_368),
.B(n_16),
.Y(n_413)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_362),
.B(n_17),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_311),
.A2(n_93),
.B(n_144),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_367),
.B(n_19),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_343),
.A2(n_91),
.B1(n_143),
.B2(n_30),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_31),
.Y(n_420)
);

O2A1O1Ixp5_ASAP7_75t_L g421 ( 
.A1(n_353),
.A2(n_94),
.B(n_142),
.C(n_32),
.Y(n_421)
);

OAI21x1_ASAP7_75t_L g422 ( 
.A1(n_356),
.A2(n_81),
.B(n_141),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_346),
.A2(n_78),
.B1(n_140),
.B2(n_34),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_367),
.A2(n_95),
.B1(n_138),
.B2(n_36),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_334),
.A2(n_77),
.B(n_134),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_363),
.A2(n_76),
.B(n_133),
.Y(n_426)
);

OR2x6_ASAP7_75t_L g427 ( 
.A(n_360),
.B(n_19),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_342),
.B(n_359),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_360),
.A2(n_96),
.B1(n_39),
.B2(n_41),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_357),
.A2(n_365),
.B(n_364),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_366),
.A2(n_97),
.B(n_43),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_359),
.A2(n_98),
.B(n_44),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_359),
.A2(n_99),
.B(n_45),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_367),
.B(n_20),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_342),
.Y(n_436)
);

AO21x1_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_20),
.B(n_49),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_385),
.A2(n_51),
.B(n_52),
.Y(n_438)
);

AOI211x1_ASAP7_75t_L g439 ( 
.A1(n_392),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_375),
.B(n_56),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_392),
.A2(n_57),
.B(n_58),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_389),
.A2(n_154),
.B(n_62),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_374),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_394),
.A2(n_65),
.B(n_67),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_377),
.A2(n_71),
.B(n_72),
.Y(n_446)
);

AOI221xp5_ASAP7_75t_SL g447 ( 
.A1(n_369),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.C(n_101),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_390),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_370),
.A2(n_105),
.B(n_106),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_376),
.A2(n_107),
.B(n_110),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_378),
.A2(n_112),
.B(n_113),
.Y(n_451)
);

AO31x2_ASAP7_75t_L g452 ( 
.A1(n_388),
.A2(n_114),
.A3(n_115),
.B(n_116),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_413),
.B(n_117),
.Y(n_453)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_386),
.A2(n_398),
.B(n_396),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_436),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_372),
.B(n_120),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_428),
.A2(n_382),
.B(n_380),
.Y(n_457)
);

BUFx12f_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

BUFx12f_ASAP7_75t_L g459 ( 
.A(n_427),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_371),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_460)
);

AOI221x1_ASAP7_75t_L g461 ( 
.A1(n_400),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.C(n_132),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_427),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_373),
.A2(n_383),
.B(n_422),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_407),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

BUFx12f_ASAP7_75t_L g467 ( 
.A(n_434),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_399),
.B(n_424),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_430),
.A2(n_391),
.B(n_420),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_395),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_409),
.A2(n_430),
.B(n_431),
.C(n_402),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_415),
.B(n_417),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_404),
.A2(n_418),
.B(n_387),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_414),
.B(n_384),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_410),
.B(n_406),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_403),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_421),
.A2(n_426),
.B(n_412),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_411),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_381),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_403),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_432),
.A2(n_433),
.B(n_425),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_423),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_429),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_419),
.A2(n_401),
.B1(n_405),
.B2(n_408),
.Y(n_486)
);

OA22x2_ASAP7_75t_L g487 ( 
.A1(n_379),
.A2(n_306),
.B1(n_256),
.B2(n_267),
.Y(n_487)
);

BUFx4f_ASAP7_75t_L g488 ( 
.A(n_416),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_379),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_389),
.A2(n_394),
.B(n_392),
.Y(n_490)
);

AOI222xp33_ASAP7_75t_L g491 ( 
.A1(n_474),
.A2(n_482),
.B1(n_485),
.B2(n_462),
.C1(n_456),
.C2(n_471),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_446),
.A2(n_441),
.B1(n_484),
.B2(n_437),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_446),
.A2(n_484),
.B1(n_487),
.B2(n_460),
.Y(n_493)
);

O2A1O1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_476),
.A2(n_475),
.B(n_453),
.C(n_466),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_442),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_481),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_463),
.A2(n_454),
.B(n_483),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_440),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_470),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_490),
.A2(n_457),
.B(n_469),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

AO21x2_ASAP7_75t_L g505 ( 
.A1(n_477),
.A2(n_473),
.B(n_445),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_478),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_455),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_458),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_464),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_481),
.Y(n_510)
);

AO32x2_ASAP7_75t_L g511 ( 
.A1(n_486),
.A2(n_448),
.A3(n_489),
.B1(n_447),
.B2(n_439),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_449),
.A2(n_443),
.B(n_451),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_464),
.Y(n_513)
);

AOI221x1_ASAP7_75t_L g514 ( 
.A1(n_477),
.A2(n_445),
.B1(n_479),
.B2(n_438),
.C(n_450),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_468),
.A2(n_461),
.B(n_444),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_444),
.Y(n_516)
);

OAI221xp5_ASAP7_75t_L g517 ( 
.A1(n_447),
.A2(n_488),
.B1(n_439),
.B2(n_459),
.C(n_452),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_488),
.B(n_452),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_452),
.A2(n_228),
.B1(n_371),
.B2(n_414),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_472),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_472),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_472),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_482),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_478),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_454),
.A2(n_469),
.B(n_457),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_442),
.B(n_374),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_472),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_482),
.A2(n_315),
.B1(n_414),
.B2(n_403),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_463),
.A2(n_389),
.B(n_454),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_463),
.A2(n_389),
.B(n_454),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_480),
.B(n_481),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_471),
.B(n_371),
.C(n_305),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_529),
.Y(n_536)
);

AND2x4_ASAP7_75t_SL g537 ( 
.A(n_501),
.B(n_529),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_513),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_513),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_535),
.A2(n_492),
.B1(n_531),
.B2(n_493),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_503),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_531),
.B(n_523),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_520),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_529),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_521),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_522),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_530),
.Y(n_547)
);

AO21x1_ASAP7_75t_SL g548 ( 
.A1(n_492),
.A2(n_493),
.B(n_518),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_495),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_532),
.A2(n_533),
.B(n_512),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_509),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

OAI21xp33_ASAP7_75t_SL g553 ( 
.A1(n_515),
.A2(n_491),
.B(n_509),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_500),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_528),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_496),
.B(n_499),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_496),
.B(n_499),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_534),
.B(n_501),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_504),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_507),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_529),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_516),
.A2(n_519),
.B1(n_494),
.B2(n_517),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_526),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_510),
.B(n_534),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

BUFx2_ASAP7_75t_SL g567 ( 
.A(n_508),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_498),
.A2(n_502),
.B(n_514),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_511),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_510),
.B(n_505),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_519),
.B(n_516),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_511),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_525),
.B(n_506),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_505),
.A2(n_535),
.B1(n_315),
.B2(n_531),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_511),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_497),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_551),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_549),
.B(n_497),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_551),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_542),
.B(n_497),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_542),
.B(n_545),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_564),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_564),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_541),
.B(n_546),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_543),
.B(n_546),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_559),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_570),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_559),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_539),
.B(n_559),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_543),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_545),
.B(n_574),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_559),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_568),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_547),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_570),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_575),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_565),
.B(n_555),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_538),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_558),
.B(n_561),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_560),
.B(n_554),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_558),
.B(n_561),
.Y(n_603)
);

INVx2_ASAP7_75t_R g604 ( 
.A(n_566),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_554),
.B(n_548),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_556),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_552),
.B(n_556),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_552),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_548),
.B(n_540),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_571),
.B(n_563),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_569),
.B(n_572),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_553),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_567),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_553),
.B(n_562),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_570),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_557),
.B(n_576),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_570),
.A2(n_576),
.B1(n_567),
.B2(n_573),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_536),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_544),
.B(n_536),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_583),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_613),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_609),
.B(n_570),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_583),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_599),
.B(n_570),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_584),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_595),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_588),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_568),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_606),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_570),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_595),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_597),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_609),
.B(n_550),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_588),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_598),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_610),
.B(n_544),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_582),
.B(n_544),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_588),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_608),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_597),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_582),
.B(n_544),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_604),
.B(n_612),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_612),
.B(n_537),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_577),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_577),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_604),
.B(n_537),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_616),
.B(n_603),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_601),
.B(n_586),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_587),
.B(n_589),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_604),
.B(n_581),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_586),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_579),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_607),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_634),
.B(n_614),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_648),
.B(n_592),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_650),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_625),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_624),
.B(n_617),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_625),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_620),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_643),
.B(n_594),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_634),
.B(n_614),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_651),
.B(n_605),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_643),
.B(n_594),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_654),
.B(n_592),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_640),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_628),
.B(n_615),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_628),
.B(n_615),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_649),
.B(n_606),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_651),
.B(n_605),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_652),
.B(n_578),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_638),
.B(n_602),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_621),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_628),
.B(n_615),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_650),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_629),
.B(n_594),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_631),
.B(n_593),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_638),
.B(n_611),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_620),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_642),
.B(n_611),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_642),
.B(n_602),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_623),
.Y(n_683)
);

AND2x4_ASAP7_75t_SL g684 ( 
.A(n_650),
.B(n_596),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_658),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_666),
.B(n_630),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_662),
.B(n_629),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_660),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_662),
.B(n_637),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_665),
.B(n_637),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_661),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_683),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_665),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_680),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_680),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_677),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_655),
.B(n_622),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_677),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_655),
.B(n_622),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_657),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_657),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_679),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_663),
.B(n_644),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_663),
.B(n_627),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_664),
.B(n_671),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_687),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_700),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_686),
.B(n_667),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_705),
.B(n_664),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_685),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_689),
.B(n_671),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_705),
.B(n_656),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_688),
.Y(n_713)
);

OAI32xp33_ASAP7_75t_L g714 ( 
.A1(n_704),
.A2(n_672),
.A3(n_670),
.B1(n_674),
.B2(n_682),
.Y(n_714)
);

OAI32xp33_ASAP7_75t_L g715 ( 
.A1(n_704),
.A2(n_673),
.A3(n_659),
.B1(n_647),
.B2(n_678),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_689),
.B(n_676),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_691),
.B(n_659),
.C(n_591),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_692),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_690),
.B(n_681),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_708),
.B(n_697),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_710),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_707),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_717),
.A2(n_706),
.B1(n_669),
.B2(n_668),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_713),
.Y(n_724)
);

AOI221xp5_ASAP7_75t_L g725 ( 
.A1(n_715),
.A2(n_702),
.B1(n_697),
.B2(n_699),
.C(n_703),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_723),
.A2(n_717),
.B(n_714),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_725),
.A2(n_596),
.B1(n_588),
.B2(n_675),
.Y(n_727)
);

OAI221xp5_ASAP7_75t_L g728 ( 
.A1(n_720),
.A2(n_724),
.B1(n_721),
.B2(n_722),
.C(n_718),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_725),
.B(n_707),
.C(n_712),
.Y(n_729)
);

AOI222xp33_ASAP7_75t_L g730 ( 
.A1(n_725),
.A2(n_719),
.B1(n_709),
.B2(n_699),
.C1(n_703),
.C2(n_693),
.Y(n_730)
);

AOI32xp33_ASAP7_75t_L g731 ( 
.A1(n_725),
.A2(n_701),
.A3(n_700),
.B1(n_698),
.B2(n_696),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_726),
.B(n_731),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_729),
.B(n_711),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_728),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_727),
.A2(n_716),
.B(n_695),
.Y(n_735)
);

NOR2x1_ASAP7_75t_L g736 ( 
.A(n_732),
.B(n_701),
.Y(n_736)
);

OAI211xp5_ASAP7_75t_L g737 ( 
.A1(n_734),
.A2(n_730),
.B(n_701),
.C(n_700),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_733),
.B(n_694),
.Y(n_738)
);

NOR2x1_ASAP7_75t_L g739 ( 
.A(n_736),
.B(n_735),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_738),
.B(n_693),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_737),
.B(n_591),
.C(n_618),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_736),
.B(n_585),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_698),
.Y(n_743)
);

XNOR2xp5_ASAP7_75t_L g744 ( 
.A(n_741),
.B(n_684),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_740),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_742),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_739),
.B(n_580),
.C(n_690),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_740),
.Y(n_748)
);

AOI211xp5_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_687),
.B(n_644),
.C(n_588),
.Y(n_749)
);

AND3x1_ASAP7_75t_L g750 ( 
.A(n_747),
.B(n_696),
.C(n_635),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_745),
.B(n_679),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_743),
.Y(n_752)
);

OAI22x1_ASAP7_75t_L g753 ( 
.A1(n_748),
.A2(n_639),
.B1(n_619),
.B2(n_668),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_746),
.B(n_681),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_751),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_SL g756 ( 
.A1(n_752),
.A2(n_744),
.B1(n_647),
.B2(n_635),
.C(n_615),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_754),
.B(n_639),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_749),
.A2(n_619),
.B(n_590),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_757),
.A2(n_753),
.B(n_750),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_755),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_756),
.A2(n_639),
.B1(n_684),
.B2(n_641),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_758),
.A2(n_639),
.B1(n_626),
.B2(n_633),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_760),
.A2(n_619),
.B(n_580),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_762),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_759),
.B(n_632),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_765),
.A2(n_761),
.B(n_619),
.Y(n_766)
);

OAI322xp33_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_600),
.A3(n_630),
.B1(n_653),
.B2(n_646),
.C1(n_645),
.C2(n_636),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_766),
.A2(n_763),
.B(n_767),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_768),
.B(n_587),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_600),
.B(n_639),
.Y(n_770)
);


endmodule