module real_jpeg_5064_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_1),
.Y(n_108)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_1),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_2),
.A2(n_42),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_42),
.B1(n_112),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_2),
.A2(n_42),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_145),
.C(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_2),
.B(n_244),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_2),
.A2(n_251),
.B(n_253),
.C(n_254),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_2),
.B(n_264),
.C(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_2),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_2),
.B(n_210),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_2),
.B(n_21),
.Y(n_290)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_4),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_5),
.Y(n_370)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_6),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_46),
.B1(n_50),
.B2(n_53),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_38),
.B1(n_53),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_7),
.A2(n_53),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_7),
.A2(n_53),
.B1(n_71),
.B2(n_183),
.Y(n_182)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_10),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_80),
.B1(n_84),
.B2(n_87),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_87),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_11),
.A2(n_87),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_11),
.A2(n_87),
.B1(n_158),
.B2(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_365),
.B(n_367),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_361),
.Y(n_14)
);

AO21x1_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_133),
.B(n_360),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_17),
.B(n_128),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_116),
.C(n_127),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_18),
.A2(n_19),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_44),
.C(n_88),
.Y(n_19)
);

XNOR2x1_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_20),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_20),
.B(n_198),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_20),
.A2(n_175),
.B1(n_176),
.B2(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_20),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_20),
.A2(n_217),
.B1(n_247),
.B2(n_257),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_20),
.B(n_167),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_20),
.A2(n_217),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_20),
.A2(n_175),
.B(n_213),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_20),
.A2(n_217),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_20),
.A2(n_217),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_31),
.B(n_40),
.Y(n_20)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_21),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_27),
.Y(n_144)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_32)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_33),
.Y(n_130)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_42),
.A2(n_68),
.B(n_71),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_44),
.A2(n_88),
.B1(n_89),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_44),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_54),
.B1(n_67),
.B2(n_79),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_45),
.A2(n_54),
.B1(n_67),
.B2(n_142),
.Y(n_338)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_67),
.B(n_79),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AO21x2_ASAP7_75t_SL g141 ( 
.A1(n_55),
.A2(n_67),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_67),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_56)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_57),
.Y(n_252)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_67),
.Y(n_244)
);

OA22x2_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_76),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_86),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_88),
.A2(n_89),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_89),
.B(n_217),
.C(n_338),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_110),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_90),
.B(n_99),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_90),
.A2(n_99),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_90),
.Y(n_208)
);

NAND2x1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_99),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_98),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_94),
.Y(n_265)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_99),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_109),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_100),
.B(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g266 ( 
.A(n_113),
.Y(n_266)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_116),
.B(n_127),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_126),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_129),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g363 ( 
.A1(n_118),
.A2(n_126),
.B(n_129),
.Y(n_363)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_128),
.B(n_363),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_128),
.B(n_363),
.Y(n_364)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_354),
.B(n_359),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_332),
.B(n_351),
.Y(n_134)
);

OAI211xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_237),
.B(n_326),
.C(n_331),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_219),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_137),
.A2(n_219),
.B(n_327),
.C(n_330),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_201),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_138),
.B(n_201),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_174),
.C(n_186),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_139),
.B(n_174),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_146),
.B1(n_172),
.B2(n_173),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_140),
.B(n_187),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_140),
.A2(n_172),
.B1(n_226),
.B2(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_141),
.B(n_207),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_141),
.A2(n_200),
.B(n_217),
.C(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_141),
.A2(n_167),
.B1(n_198),
.B2(n_223),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_141),
.A2(n_198),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_146),
.A2(n_197),
.B(n_199),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_167),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_147),
.A2(n_167),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_147),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_154),
.B1(n_160),
.B2(n_164),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_152),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_154),
.B1(n_189),
.B2(n_195),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_167),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_167),
.A2(n_223),
.B1(n_243),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_167),
.A2(n_223),
.B1(n_261),
.B2(n_262),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_167),
.A2(n_223),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_167),
.A2(n_198),
.B(n_249),
.C(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_167),
.B(n_198),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_167),
.A2(n_188),
.B1(n_223),
.B2(n_317),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_185),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_179),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_190),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_207)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_197),
.B(n_199),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_188),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_198),
.A2(n_206),
.B(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_198),
.B(n_234),
.C(n_289),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AND3x1_ASAP7_75t_L g319 ( 
.A(n_200),
.B(n_296),
.C(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_218),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_205),
.B(n_212),
.C(n_218),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

FAx1_ASAP7_75t_L g334 ( 
.A(n_211),
.B(n_335),
.CI(n_340),
.CON(n_334),
.SN(n_334)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_217),
.B(n_346),
.C(n_350),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_235),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_220),
.B(n_235),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.C(n_225),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_221),
.B(n_222),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_243),
.C(n_245),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_223),
.B(n_286),
.C(n_293),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_225),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_227),
.A2(n_228),
.B1(n_234),
.B2(n_245),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_234),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_234),
.A2(n_245),
.B1(n_250),
.B2(n_256),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_234),
.A2(n_245),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_250),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_308),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_298),
.B(n_307),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_284),
.B(n_297),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_258),
.B(n_283),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_245),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_257),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_270),
.B(n_282),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_267),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_294),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_321),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_311),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_318),
.C(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_328),
.B(n_329),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_342),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_341),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_334),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_341),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_343),
.Y(n_353)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_342),
.A2(n_352),
.B(n_353),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_350),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_358),
.Y(n_359)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

INVx8_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_366),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

BUFx12f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);


endmodule