module fake_jpeg_7431_n_234 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_23),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_27),
.B1(n_26),
.B2(n_20),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_29),
.B1(n_14),
.B2(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_55),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_14),
.B1(n_26),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_15),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_24),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_61),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_57),
.B1(n_25),
.B2(n_17),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_37),
.C(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_69),
.B1(n_58),
.B2(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_48),
.B1(n_43),
.B2(n_49),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_14),
.B1(n_17),
.B2(n_25),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_39),
.C(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_39),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_15),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_57),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_56),
.B1(n_49),
.B2(n_53),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_84),
.B1(n_76),
.B2(n_74),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_91),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_56),
.B1(n_49),
.B2(n_48),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_88),
.B1(n_96),
.B2(n_21),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_54),
.B1(n_48),
.B2(n_32),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_32),
.B1(n_78),
.B2(n_45),
.Y(n_118)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_94),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_101),
.B(n_21),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_72),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_112),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_71),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_38),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_70),
.B1(n_68),
.B2(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_59),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_68),
.B1(n_72),
.B2(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_64),
.B1(n_62),
.B2(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_10),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_12),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_89),
.A3(n_83),
.B1(n_97),
.B2(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_83),
.A3(n_85),
.B1(n_22),
.B2(n_17),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_0),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_143),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_108),
.B1(n_99),
.B2(n_82),
.Y(n_161)
);

CKINVDCx12_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_110),
.B(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_12),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_132),
.C(n_138),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_107),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_152),
.C(n_153),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_133),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_149),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_22),
.B(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_115),
.B1(n_114),
.B2(n_118),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_157),
.B1(n_126),
.B2(n_127),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_117),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_117),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_86),
.C(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_162),
.B1(n_136),
.B2(n_137),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_108),
.B1(n_105),
.B2(n_119),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_132),
.B1(n_129),
.B2(n_139),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_168),
.B1(n_162),
.B2(n_159),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_135),
.B1(n_139),
.B2(n_141),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_175),
.B(n_179),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_124),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_178),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_146),
.B1(n_156),
.B2(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_125),
.B1(n_127),
.B2(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_9),
.B(n_2),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_152),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_171),
.B(n_163),
.C(n_165),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_153),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_154),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_178),
.C(n_164),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_196),
.C(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_175),
.C(n_148),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_179),
.B1(n_174),
.B2(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_86),
.C(n_100),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_93),
.C(n_22),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_203),
.C(n_38),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_38),
.C(n_45),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_198),
.B(n_180),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_205),
.B(n_8),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_201),
.A2(n_189),
.B(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_189),
.B(n_2),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_212),
.C(n_13),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_7),
.B(n_3),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_4),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_210),
.B(n_6),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_216),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_207),
.C(n_205),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_221),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_9),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_215),
.B(n_5),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_227),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_9),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_11),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_226),
.C(n_221),
.Y(n_231)
);

AO21x2_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_225),
.B(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_13),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_1),
.Y(n_234)
);


endmodule