module fake_netlist_6_1886_n_2299 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2299);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2299;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_2292;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_92),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_90),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_47),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_91),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_99),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_177),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_42),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_45),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_47),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_116),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_19),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_137),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_185),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_30),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_193),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_141),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_26),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_43),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_103),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_129),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_115),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_88),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_48),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_166),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_89),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_71),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_10),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVxp33_ASAP7_75t_SL g258 ( 
.A(n_39),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_64),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_168),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_148),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_61),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_100),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_164),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_178),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_126),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_145),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_188),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_49),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_45),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_139),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_21),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_73),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_201),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_86),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_63),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_103),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_58),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_128),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_218),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_170),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_61),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_197),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_25),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_77),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_102),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_202),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_114),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_40),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_39),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_13),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_87),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_58),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_144),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_41),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_120),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_86),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_112),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_135),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_198),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_181),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_186),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_189),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_53),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_123),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_206),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_92),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_85),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_169),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_77),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_40),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_173),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_105),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_63),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_134),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_102),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_119),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_207),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_184),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_80),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_110),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_1),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_36),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_111),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_90),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_64),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_122),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_194),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_105),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_55),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_104),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_133),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_132),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_195),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_21),
.Y(n_341)
);

BUFx8_ASAP7_75t_SL g342 ( 
.A(n_7),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_143),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_159),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_78),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_131),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_138),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_200),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_97),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_149),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_22),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_117),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_17),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_179),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_66),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_88),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_203),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_217),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_70),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_11),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_82),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_6),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_150),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_204),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_209),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_42),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_196),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_84),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_43),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_162),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_153),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_174),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_16),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_7),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_30),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_100),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_38),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_54),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_65),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_154),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_0),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_37),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_67),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_32),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_44),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_124),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_53),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_95),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_29),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_83),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_38),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_46),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_57),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_213),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_140),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_55),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_71),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_11),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_15),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_31),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_158),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_49),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_17),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_212),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_205),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_2),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_14),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_51),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_36),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_15),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_35),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_37),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_94),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_81),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_96),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_83),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_97),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_3),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_51),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_74),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_107),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_214),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_0),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_32),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_6),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_121),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_76),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_125),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_163),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_73),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_84),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_220),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_228),
.B(n_2),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_342),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_230),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_266),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_320),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_320),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_320),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_320),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_233),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_269),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_225),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_236),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_262),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_320),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_310),
.B(n_3),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_262),
.B(n_4),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_311),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_320),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_407),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_407),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_407),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_239),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_338),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_240),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_243),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_356),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_333),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_244),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_248),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_428),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_333),
.B(n_4),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_301),
.B(n_5),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_414),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_301),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_347),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_405),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_250),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_348),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_428),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_253),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_261),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_414),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_265),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_425),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_310),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_267),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_242),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_425),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_425),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_277),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_425),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_425),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_270),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_273),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_225),
.A2(n_8),
.B(n_9),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_276),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_229),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_229),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_229),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_281),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_282),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_242),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_245),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_245),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_285),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_245),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_290),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_288),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_241),
.B(n_8),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_292),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_251),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_304),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_306),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_308),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_309),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_251),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_321),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_241),
.B(n_9),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_325),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_330),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_251),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_278),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_278),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_278),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_341),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_334),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_343),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_221),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_341),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_344),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_341),
.Y(n_531)
);

BUFx2_ASAP7_75t_SL g532 ( 
.A(n_241),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_221),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_346),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_258),
.B(n_10),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_357),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_358),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_249),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_242),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_228),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_219),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_364),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_465),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_437),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_225),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_465),
.Y(n_553)
);

AND3x1_ASAP7_75t_L g554 ( 
.A(n_448),
.B(n_402),
.C(n_360),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_432),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_360),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_435),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_436),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_439),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_532),
.B(n_373),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_440),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_475),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_440),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_441),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_446),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_444),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_446),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_465),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_442),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_539),
.B(n_283),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_450),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_477),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_542),
.Y(n_576)
);

NAND2x1_ASAP7_75t_L g577 ( 
.A(n_443),
.B(n_428),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_477),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_449),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_477),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_455),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_532),
.B(n_360),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_457),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_471),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_458),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_509),
.B(n_402),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_477),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_477),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_472),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_473),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_459),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_463),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_485),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_451),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_471),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_464),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_474),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_447),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_443),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_451),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_486),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_478),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_518),
.B(n_402),
.Y(n_604)
);

INVx6_ASAP7_75t_L g605 ( 
.A(n_433),
.Y(n_605)
);

BUFx8_ASAP7_75t_L g606 ( 
.A(n_468),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_468),
.B(n_428),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_493),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_496),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_460),
.B(n_354),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_495),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_452),
.B(n_283),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_500),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_453),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_453),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_454),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_505),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_454),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_443),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_480),
.B(n_365),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_456),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_483),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_456),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_461),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_495),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_494),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_433),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_466),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_510),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_541),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_R g633 ( 
.A(n_512),
.B(n_370),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_555),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_604),
.B(n_514),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_573),
.B(n_498),
.Y(n_636)
);

BUFx6f_ASAP7_75t_SL g637 ( 
.A(n_573),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_605),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_605),
.B(n_536),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_604),
.B(n_515),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_560),
.B(n_520),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_564),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_595),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_595),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_560),
.A2(n_462),
.B1(n_507),
.B2(n_501),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_586),
.B(n_527),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_600),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_595),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_621),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_605),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_586),
.B(n_530),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_550),
.B(n_535),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_612),
.B(n_283),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_633),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_550),
.B(n_573),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_607),
.Y(n_656)
);

BUFx6f_ASAP7_75t_SL g657 ( 
.A(n_573),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_546),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_616),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_550),
.B(n_537),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_616),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_613),
.B(n_498),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_R g663 ( 
.A(n_562),
.B(n_434),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_605),
.B(n_538),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_546),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_633),
.B(n_543),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_564),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_616),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_605),
.B(n_467),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_582),
.B(n_445),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_600),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_558),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_557),
.B(n_513),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_622),
.Y(n_674)
);

INVxp33_ASAP7_75t_L g675 ( 
.A(n_584),
.Y(n_675)
);

INVx4_ASAP7_75t_SL g676 ( 
.A(n_607),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_547),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_584),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_553),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_613),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_566),
.B(n_517),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_568),
.B(n_581),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_622),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_547),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_607),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_553),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_607),
.B(n_466),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_SL g688 ( 
.A1(n_611),
.A2(n_490),
.B1(n_508),
.B2(n_502),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_607),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_607),
.B(n_582),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_551),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_613),
.B(n_503),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_607),
.A2(n_443),
.B1(n_234),
.B2(n_254),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_585),
.B(n_519),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_554),
.B(n_503),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_552),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_599),
.B(n_497),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_591),
.B(n_487),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_592),
.B(n_526),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_607),
.B(n_469),
.Y(n_703)
);

AND2x6_ASAP7_75t_L g704 ( 
.A(n_612),
.B(n_318),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_597),
.B(n_487),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_559),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_599),
.A2(n_540),
.B1(n_502),
.B2(n_271),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_596),
.B(n_594),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_598),
.B(n_540),
.Y(n_709)
);

NAND2x1p5_ASAP7_75t_L g710 ( 
.A(n_612),
.B(n_249),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_602),
.B(n_354),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_612),
.B(n_318),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_576),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_612),
.A2(n_234),
.B1(n_254),
.B2(n_232),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_632),
.B(n_497),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_608),
.B(n_610),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_554),
.A2(n_339),
.B1(n_318),
.B2(n_246),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_572),
.Y(n_718)
);

AO22x2_ASAP7_75t_L g719 ( 
.A1(n_594),
.A2(n_339),
.B1(n_246),
.B2(n_271),
.Y(n_719)
);

INVx5_ASAP7_75t_L g720 ( 
.A(n_612),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_559),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_SL g722 ( 
.A1(n_606),
.A2(n_272),
.B1(n_326),
.B2(n_231),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_553),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_561),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_561),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_624),
.Y(n_726)
);

AO22x2_ASAP7_75t_L g727 ( 
.A1(n_556),
.A2(n_339),
.B1(n_419),
.B2(n_387),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_556),
.B(n_469),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_626),
.B(n_499),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_632),
.B(n_499),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_553),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_553),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_631),
.B(n_354),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_575),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_614),
.B(n_222),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_628),
.B(n_504),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_563),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_565),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_618),
.B(n_354),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_628),
.B(n_223),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_596),
.Y(n_742)
);

AND2x6_ASAP7_75t_L g743 ( 
.A(n_626),
.B(n_428),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_576),
.A2(n_419),
.B1(n_423),
.B2(n_387),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_600),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_562),
.B(n_257),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_626),
.A2(n_226),
.B1(n_227),
.B2(n_224),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_565),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_567),
.B(n_504),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_624),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_575),
.Y(n_751)
);

INVx4_ASAP7_75t_SL g752 ( 
.A(n_626),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_606),
.B(n_363),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_567),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_569),
.B(n_470),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_569),
.B(n_470),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_571),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_626),
.B(n_506),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_624),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_571),
.B(n_574),
.Y(n_760)
);

AND2x6_ASAP7_75t_L g761 ( 
.A(n_626),
.B(n_428),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_574),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_606),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_606),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_601),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_601),
.B(n_476),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_579),
.Y(n_767)
);

AO21x2_ASAP7_75t_L g768 ( 
.A1(n_609),
.A2(n_259),
.B(n_257),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_609),
.B(n_476),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_615),
.B(n_506),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_615),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_583),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_617),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_587),
.Y(n_774)
);

INVx6_ASAP7_75t_L g775 ( 
.A(n_549),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_617),
.B(n_237),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_544),
.B(n_259),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_619),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_619),
.B(n_625),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_625),
.Y(n_780)
);

AND2x6_ASAP7_75t_L g781 ( 
.A(n_544),
.B(n_268),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_629),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_575),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_589),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_629),
.Y(n_785)
);

AND2x6_ASAP7_75t_L g786 ( 
.A(n_544),
.B(n_268),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_630),
.B(n_238),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_729),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_635),
.B(n_603),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_729),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_646),
.A2(n_394),
.B1(n_395),
.B2(n_371),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_651),
.B(n_630),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_637),
.A2(n_422),
.B1(n_426),
.B2(n_401),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_670),
.B(n_511),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_655),
.B(n_620),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_729),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_758),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_758),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_670),
.B(n_511),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_680),
.A2(n_300),
.B1(n_302),
.B2(n_286),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_680),
.B(n_620),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_758),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_640),
.B(n_620),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_697),
.A2(n_300),
.B1(n_302),
.B2(n_286),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_652),
.B(n_623),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_637),
.A2(n_429),
.B1(n_307),
.B2(n_312),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_660),
.B(n_620),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_708),
.B(n_423),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_697),
.A2(n_307),
.B1(n_312),
.B2(n_305),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_664),
.B(n_549),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_720),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_636),
.B(n_549),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_636),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_636),
.B(n_549),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_654),
.B(n_746),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_706),
.B(n_587),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_649),
.B(n_479),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_658),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_699),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_658),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_706),
.B(n_587),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_757),
.B(n_587),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_SL g823 ( 
.A1(n_688),
.A2(n_381),
.B1(n_382),
.B2(n_355),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_697),
.A2(n_315),
.B1(n_323),
.B2(n_305),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_763),
.B(n_315),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_765),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_735),
.B(n_627),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_757),
.B(n_588),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_765),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_699),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_665),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_690),
.A2(n_324),
.B1(n_327),
.B2(n_323),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_762),
.B(n_588),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_654),
.B(n_363),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_641),
.B(n_590),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_675),
.B(n_247),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_762),
.B(n_588),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_715),
.B(n_516),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_638),
.B(n_588),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_771),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_771),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_638),
.B(n_545),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_780),
.Y(n_843)
);

AO22x1_ASAP7_75t_L g844 ( 
.A1(n_653),
.A2(n_327),
.B1(n_340),
.B2(n_324),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_637),
.A2(n_350),
.B1(n_352),
.B2(n_340),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_746),
.B(n_649),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_650),
.B(n_545),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_650),
.B(n_545),
.Y(n_848)
);

NOR2x1p5_ASAP7_75t_L g849 ( 
.A(n_708),
.B(n_232),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_728),
.B(n_548),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_710),
.B(n_548),
.Y(n_851)
);

AND3x1_ASAP7_75t_L g852 ( 
.A(n_645),
.B(n_289),
.C(n_284),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_720),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_L g854 ( 
.A(n_736),
.B(n_284),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_665),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_742),
.B(n_255),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_713),
.B(n_289),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_715),
.B(n_516),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_714),
.A2(n_350),
.B1(n_367),
.B2(n_352),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_657),
.A2(n_372),
.B1(n_380),
.B2(n_367),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_657),
.A2(n_380),
.B1(n_386),
.B2(n_372),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_684),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_713),
.B(n_293),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_741),
.B(n_666),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_677),
.A2(n_386),
.B(n_404),
.C(n_577),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_L g866 ( 
.A(n_720),
.B(n_235),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_684),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_711),
.B(n_256),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_710),
.B(n_548),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_710),
.B(n_662),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_730),
.B(n_521),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_736),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_662),
.B(n_570),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_691),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_662),
.B(n_570),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_707),
.B(n_363),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_691),
.Y(n_877)
);

BUFx8_ASAP7_75t_L g878 ( 
.A(n_764),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_692),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_693),
.Y(n_880)
);

AND2x6_ASAP7_75t_SL g881 ( 
.A(n_705),
.B(n_293),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_678),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_L g883 ( 
.A(n_747),
.B(n_263),
.C(n_260),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_724),
.A2(n_778),
.B(n_725),
.C(n_760),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_774),
.A2(n_577),
.B(n_404),
.C(n_570),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_780),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_693),
.B(n_575),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_693),
.B(n_575),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_692),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_698),
.B(n_575),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_733),
.B(n_264),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_720),
.A2(n_580),
.B(n_578),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_657),
.A2(n_390),
.B1(n_415),
.B2(n_363),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_672),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_698),
.B(n_578),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_701),
.B(n_578),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_642),
.B(n_297),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_L g898 ( 
.A(n_730),
.B(n_787),
.C(n_776),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_669),
.A2(n_235),
.B1(n_479),
.B2(n_481),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_722),
.B(n_275),
.C(n_274),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_701),
.B(n_721),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_721),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_737),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_653),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_737),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_738),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_739),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_739),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_682),
.B(n_279),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_709),
.B(n_481),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_748),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_653),
.A2(n_235),
.B1(n_393),
.B2(n_398),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_748),
.B(n_578),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_754),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_754),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_773),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_773),
.B(n_578),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_782),
.B(n_578),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_763),
.B(n_280),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_782),
.B(n_580),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_SL g921 ( 
.A1(n_764),
.A2(n_242),
.B1(n_252),
.B2(n_412),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_785),
.B(n_580),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_785),
.B(n_580),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_639),
.B(n_521),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_667),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_669),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_643),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_740),
.B(n_287),
.Y(n_928)
);

AO22x1_ASAP7_75t_L g929 ( 
.A1(n_653),
.A2(n_388),
.B1(n_297),
.B2(n_298),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_653),
.A2(n_235),
.B1(n_388),
.B2(n_398),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_749),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_720),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_643),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_644),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_639),
.B(n_291),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_669),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_743),
.B(n_580),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_743),
.B(n_580),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_743),
.B(n_761),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_749),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_770),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_770),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_743),
.B(n_593),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_653),
.A2(n_235),
.B1(n_298),
.B2(n_303),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_669),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_672),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_639),
.B(n_303),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_743),
.B(n_761),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_743),
.B(n_761),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_685),
.B(n_294),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_644),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_L g952 ( 
.A(n_761),
.B(n_235),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_761),
.B(n_593),
.Y(n_953)
);

OAI22xp33_ASAP7_75t_L g954 ( 
.A1(n_639),
.A2(n_753),
.B1(n_744),
.B2(n_779),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_648),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_685),
.B(n_600),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_717),
.A2(n_235),
.B1(n_482),
.B2(n_484),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_685),
.B(n_295),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_761),
.B(n_593),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_794),
.B(n_717),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_794),
.B(n_717),
.Y(n_961)
);

BUFx2_ASAP7_75t_SL g962 ( 
.A(n_904),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_925),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_792),
.B(n_752),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_894),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_788),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_894),
.Y(n_967)
);

BUFx12f_ASAP7_75t_L g968 ( 
.A(n_878),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_889),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_788),
.Y(n_970)
);

NAND2xp33_ASAP7_75t_SL g971 ( 
.A(n_815),
.B(n_716),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_799),
.B(n_752),
.Y(n_972)
);

OR2x4_ASAP7_75t_L g973 ( 
.A(n_808),
.B(n_864),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_889),
.Y(n_974)
);

AO22x1_ASAP7_75t_L g975 ( 
.A1(n_926),
.A2(n_712),
.B1(n_704),
.B2(n_777),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_924),
.A2(n_717),
.B1(n_712),
.B2(n_704),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_811),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_799),
.B(n_727),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_796),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_882),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_818),
.B(n_752),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_924),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_790),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_818),
.B(n_752),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_790),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_811),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_926),
.B(n_676),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_797),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_789),
.B(n_673),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_897),
.Y(n_991)
);

INVx3_ASAP7_75t_SL g992 ( 
.A(n_946),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_R g993 ( 
.A(n_946),
.B(n_634),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_820),
.B(n_704),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_820),
.B(n_704),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_902),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_797),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_936),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_831),
.B(n_855),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_902),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_936),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_905),
.Y(n_1002)
);

AND3x1_ASAP7_75t_SL g1003 ( 
.A(n_849),
.B(n_329),
.C(n_322),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_798),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_798),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_945),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_872),
.B(n_727),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_831),
.B(n_704),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_880),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_880),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_905),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_906),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_802),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_802),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_855),
.B(n_704),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_R g1016 ( 
.A(n_827),
.B(n_634),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_826),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_945),
.B(n_676),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_880),
.A2(n_712),
.B1(n_768),
.B2(n_727),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_906),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_811),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_878),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_907),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_947),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_862),
.B(n_867),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_805),
.B(n_681),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_904),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_878),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_826),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_881),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_898),
.A2(n_712),
.B1(n_696),
.B2(n_702),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_SL g1032 ( 
.A(n_846),
.B(n_663),
.C(n_718),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_947),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_872),
.B(n_772),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_862),
.B(n_712),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_854),
.Y(n_1036)
);

AO22x1_ASAP7_75t_L g1037 ( 
.A1(n_900),
.A2(n_712),
.B1(n_781),
.B2(n_777),
.Y(n_1037)
);

INVx3_ASAP7_75t_SL g1038 ( 
.A(n_823),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_897),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_931),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_829),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_811),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_829),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_811),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_840),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_838),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_867),
.B(n_874),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_907),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_904),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_870),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_939),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_874),
.B(n_768),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_813),
.A2(n_768),
.B1(n_727),
.B2(n_719),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_931),
.B(n_719),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_L g1055 ( 
.A(n_948),
.B(n_656),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_840),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_877),
.B(n_679),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_841),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_940),
.B(n_676),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_893),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_877),
.B(n_679),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_940),
.B(n_676),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_841),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_SL g1064 ( 
.A(n_876),
.B(n_767),
.C(n_718),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_819),
.B(n_767),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_911),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_835),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_954),
.A2(n_813),
.B1(n_935),
.B2(n_830),
.Y(n_1068)
);

INVxp33_ASAP7_75t_L g1069 ( 
.A(n_836),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_879),
.B(n_679),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_879),
.B(n_686),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_819),
.B(n_685),
.Y(n_1072)
);

BUFx12f_ASAP7_75t_L g1073 ( 
.A(n_849),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_949),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_903),
.B(n_686),
.Y(n_1075)
);

INVxp67_ASAP7_75t_SL g1076 ( 
.A(n_887),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_911),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_941),
.B(n_784),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_843),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_852),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_SL g1081 ( 
.A(n_834),
.B(n_299),
.C(n_296),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_916),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_808),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_830),
.B(n_700),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_909),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_854),
.Y(n_1086)
);

NOR2x1p5_ASAP7_75t_L g1087 ( 
.A(n_857),
.B(n_313),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_838),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_916),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_853),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_903),
.B(n_686),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_R g1092 ( 
.A(n_941),
.B(n_772),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_857),
.B(n_772),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_SL g1094 ( 
.A(n_825),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_843),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_886),
.Y(n_1096)
);

AND3x2_ASAP7_75t_SL g1097 ( 
.A(n_957),
.B(n_719),
.C(n_886),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_853),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_927),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_908),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_858),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_910),
.B(n_817),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_942),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_SL g1104 ( 
.A(n_868),
.B(n_316),
.C(n_314),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_942),
.B(n_685),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_807),
.A2(n_687),
.B1(n_703),
.B2(n_689),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_SL g1107 ( 
.A(n_891),
.B(n_319),
.C(n_317),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_928),
.B(n_331),
.C(n_328),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_832),
.A2(n_719),
.B1(n_786),
.B2(n_781),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_858),
.B(n_656),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_927),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_933),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_871),
.B(n_648),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_863),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_853),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_795),
.A2(n_689),
.B(n_656),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_825),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_914),
.B(n_723),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_914),
.B(n_915),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_933),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_915),
.B(n_723),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_932),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_871),
.B(n_884),
.Y(n_1123)
);

AND2x6_ASAP7_75t_SL g1124 ( 
.A(n_856),
.B(n_322),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_934),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_919),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_934),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_951),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_863),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_R g1130 ( 
.A(n_866),
.B(n_772),
.Y(n_1130)
);

AND2x4_ASAP7_75t_SL g1131 ( 
.A(n_825),
.B(n_252),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_901),
.B(n_723),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_825),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_951),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_801),
.B(n_732),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_803),
.B(n_732),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_800),
.A2(n_786),
.B1(n_777),
.B2(n_781),
.Y(n_1137)
);

NOR3xp33_ASAP7_75t_SL g1138 ( 
.A(n_883),
.B(n_345),
.C(n_335),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_816),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_899),
.A2(n_656),
.B1(n_689),
.B2(n_775),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_932),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_955),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_873),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_804),
.B(n_732),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_SL g1146 ( 
.A(n_865),
.B(n_351),
.C(n_349),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_875),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_888),
.Y(n_1148)
);

AND2x6_ASAP7_75t_SL g1149 ( 
.A(n_821),
.B(n_329),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_809),
.B(n_353),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_991),
.A2(n_921),
.B(n_791),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1052),
.A2(n_810),
.A3(n_850),
.B(n_890),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_SL g1153 ( 
.A(n_962),
.B(n_851),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1031),
.B(n_806),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1019),
.A2(n_885),
.B(n_895),
.Y(n_1155)
);

NAND2x1_ASAP7_75t_L g1156 ( 
.A(n_1044),
.B(n_734),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1049),
.A2(n_869),
.B(n_814),
.Y(n_1157)
);

AOI211x1_ASAP7_75t_L g1158 ( 
.A1(n_1054),
.A2(n_929),
.B(n_844),
.C(n_828),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_983),
.B(n_822),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_972),
.A2(n_812),
.B(n_896),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1026),
.B(n_793),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1046),
.B(n_824),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_990),
.B(n_860),
.C(n_845),
.Y(n_1163)
);

AO22x2_ASAP7_75t_L g1164 ( 
.A1(n_1007),
.A2(n_336),
.B1(n_337),
.B2(n_332),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_999),
.A2(n_917),
.A3(n_918),
.B(n_913),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1068),
.A2(n_861),
.B(n_833),
.C(n_837),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1123),
.A2(n_859),
.B1(n_839),
.B2(n_842),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_981),
.A2(n_922),
.B(n_920),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_971),
.A2(n_958),
.B1(n_950),
.B2(n_866),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1049),
.A2(n_848),
.B(n_847),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1046),
.B(n_929),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1101),
.B(n_912),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1069),
.B(n_923),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_969),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1136),
.A2(n_756),
.B(n_755),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_985),
.A2(n_892),
.B(n_937),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1076),
.A2(n_943),
.B(n_938),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_964),
.A2(n_959),
.B(n_953),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1101),
.B(n_844),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1039),
.B(n_930),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1147),
.A2(n_952),
.B(n_944),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_994),
.A2(n_783),
.B(n_734),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1067),
.A2(n_952),
.B1(n_775),
.B2(n_734),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_1090),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_966),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_SL g1186 ( 
.A(n_962),
.B(n_731),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_995),
.A2(n_783),
.B(n_661),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1116),
.A2(n_956),
.B(n_751),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1088),
.B(n_766),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_963),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_984),
.Y(n_1191)
);

AOI221x1_ASAP7_75t_L g1192 ( 
.A1(n_978),
.A2(n_769),
.B1(n_683),
.B2(n_759),
.C(n_750),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_1025),
.A2(n_661),
.B(n_659),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1147),
.A2(n_695),
.B(n_668),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_960),
.B(n_659),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_963),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1008),
.A2(n_783),
.B(n_674),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1040),
.B(n_668),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1033),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_974),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1015),
.A2(n_683),
.B(n_674),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1040),
.B(n_694),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_960),
.B(n_694),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1035),
.A2(n_750),
.B(n_726),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1144),
.A2(n_759),
.B(n_726),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1090),
.A2(n_956),
.B(n_751),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_974),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_996),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_993),
.Y(n_1209)
);

OAI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1114),
.A2(n_362),
.B(n_359),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_983),
.B(n_731),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1144),
.A2(n_523),
.B(n_522),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_961),
.B(n_522),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_996),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1000),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1144),
.A2(n_524),
.B(n_523),
.Y(n_1216)
);

BUFx12f_ASAP7_75t_L g1217 ( 
.A(n_968),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_1110),
.A2(n_361),
.B(n_332),
.C(n_336),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1000),
.Y(n_1219)
);

BUFx10_ASAP7_75t_L g1220 ( 
.A(n_965),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1103),
.B(n_775),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1123),
.A2(n_1148),
.B(n_976),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1103),
.B(n_775),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_965),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1047),
.A2(n_525),
.B(n_524),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1123),
.A2(n_786),
.B(n_781),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1119),
.A2(n_529),
.B(n_525),
.Y(n_1227)
);

AOI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1057),
.A2(n_484),
.B(n_482),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1100),
.A2(n_391),
.A3(n_337),
.B(n_361),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1002),
.Y(n_1230)
);

NOR2xp67_ASAP7_75t_L g1231 ( 
.A(n_1107),
.B(n_967),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1061),
.A2(n_1071),
.B(n_1070),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1148),
.A2(n_781),
.B(n_777),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_961),
.B(n_529),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_973),
.A2(n_731),
.B1(n_751),
.B2(n_417),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1084),
.B(n_731),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1113),
.B(n_777),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_977),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1113),
.B(n_531),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_SL g1240 ( 
.A1(n_1053),
.A2(n_377),
.B(n_368),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1145),
.A2(n_781),
.B(n_777),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1129),
.B(n_786),
.Y(n_1242)
);

BUFx4_ASAP7_75t_SL g1243 ( 
.A(n_1022),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_970),
.B(n_786),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1106),
.A2(n_786),
.B(n_489),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1078),
.B(n_731),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1002),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_970),
.B(n_366),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_967),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1009),
.A2(n_751),
.B(n_593),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1090),
.A2(n_671),
.B(n_647),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1090),
.A2(n_671),
.B(n_647),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1075),
.A2(n_533),
.B(n_531),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1060),
.A2(n_412),
.B1(n_252),
.B2(n_374),
.Y(n_1254)
);

NOR2x1_ASAP7_75t_SL g1255 ( 
.A(n_1009),
.B(n_368),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1098),
.A2(n_671),
.B(n_647),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1059),
.B(n_1062),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1078),
.B(n_369),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_979),
.B(n_375),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_979),
.B(n_376),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1098),
.A2(n_745),
.B(n_593),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1098),
.A2(n_745),
.B(n_593),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1091),
.A2(n_488),
.B(n_489),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1083),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_982),
.B(n_379),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1083),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1011),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1098),
.A2(n_1122),
.B(n_1115),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1011),
.A2(n_416),
.A3(n_378),
.B(n_384),
.Y(n_1269)
);

AOI211x1_ASAP7_75t_L g1270 ( 
.A1(n_1054),
.A2(n_378),
.B(n_416),
.C(n_384),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1098),
.A2(n_745),
.B(n_600),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1132),
.A2(n_492),
.B(n_491),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1118),
.A2(n_1077),
.B(n_1020),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_973),
.B(n_383),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1078),
.B(n_1039),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_980),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1082),
.A2(n_492),
.B(n_491),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_992),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1012),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1082),
.A2(n_431),
.B(n_393),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1059),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1122),
.A2(n_600),
.B(n_431),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1122),
.A2(n_600),
.B(n_377),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_992),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1122),
.A2(n_391),
.B(n_109),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_968),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1082),
.A2(n_235),
.B(n_216),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_978),
.B(n_252),
.Y(n_1288)
);

AOI21x1_ASAP7_75t_L g1289 ( 
.A1(n_975),
.A2(n_235),
.B(n_113),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1132),
.A2(n_430),
.B(n_427),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1033),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_982),
.B(n_385),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1132),
.A2(n_421),
.B(n_420),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1089),
.A2(n_235),
.B(n_215),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_973),
.B(n_389),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1009),
.A2(n_210),
.B(n_208),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1122),
.A2(n_187),
.B(n_127),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1007),
.B(n_374),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1024),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_SL g1300 ( 
.A1(n_1012),
.A2(n_192),
.B(n_190),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_989),
.B(n_392),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_989),
.B(n_396),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_997),
.A2(n_418),
.B(n_413),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_980),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1020),
.A2(n_183),
.B(n_182),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1089),
.A2(n_175),
.B(n_167),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1115),
.A2(n_165),
.B(n_130),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1089),
.A2(n_161),
.B(n_160),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1022),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_997),
.B(n_397),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1023),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1161),
.B(n_1067),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1185),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_SL g1314 ( 
.A1(n_1222),
.A2(n_984),
.B(n_1094),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1205),
.A2(n_1048),
.B(n_1023),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1174),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1205),
.A2(n_1066),
.B(n_1048),
.Y(n_1317)
);

INVx8_ASAP7_75t_L g1318 ( 
.A(n_1184),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1212),
.A2(n_1066),
.B(n_1096),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1196),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1196),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1195),
.B(n_1203),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1212),
.A2(n_1096),
.B(n_1029),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1163),
.A2(n_1036),
.B1(n_1086),
.B2(n_1060),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1154),
.A2(n_1080),
.B1(n_1038),
.B2(n_1085),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1304),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1288),
.B(n_1001),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1151),
.A2(n_1093),
.B(n_1080),
.C(n_1032),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1216),
.A2(n_1029),
.B(n_1017),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1192),
.A2(n_1041),
.B(n_1017),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1174),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1216),
.A2(n_1043),
.B(n_1041),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1274),
.A2(n_1038),
.B1(n_1085),
.B2(n_1087),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1201),
.A2(n_1197),
.B(n_1187),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1257),
.B(n_1001),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1166),
.A2(n_1102),
.B(n_1135),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1299),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1250),
.A2(n_1142),
.B(n_1115),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1214),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1214),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1295),
.A2(n_1150),
.B1(n_1117),
.B2(n_1126),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1192),
.A2(n_1045),
.B(n_1043),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1257),
.B(n_1281),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1288),
.B(n_1006),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1291),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1275),
.A2(n_1150),
.B1(n_1117),
.B2(n_1126),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1200),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1201),
.A2(n_1056),
.B(n_1045),
.Y(n_1348)
);

BUFx4f_ASAP7_75t_SL g1349 ( 
.A(n_1217),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1215),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1181),
.A2(n_1135),
.B(n_1005),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1215),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1187),
.A2(n_1058),
.B(n_1056),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1257),
.B(n_1006),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1219),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1219),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1254),
.A2(n_1016),
.B1(n_1064),
.B2(n_1030),
.C(n_1104),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1230),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1225),
.A2(n_1227),
.B(n_1253),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1173),
.A2(n_1093),
.B(n_1108),
.C(n_1081),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1197),
.A2(n_1063),
.B(n_1058),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1182),
.A2(n_1079),
.B(n_1063),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1230),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1225),
.A2(n_1095),
.B(n_1079),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1182),
.A2(n_1095),
.B(n_1120),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1281),
.B(n_1004),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1281),
.B(n_1004),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1159),
.A2(n_1073),
.B1(n_1094),
.B2(n_1050),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1213),
.B(n_1005),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_SL g1370 ( 
.A1(n_1300),
.A2(n_1014),
.B(n_1013),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1195),
.B(n_1013),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1278),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1258),
.A2(n_1138),
.B(n_1034),
.C(n_1014),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1203),
.B(n_1121),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1209),
.A2(n_1133),
.B1(n_1073),
.B2(n_1030),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1168),
.A2(n_1125),
.B(n_1127),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1237),
.A2(n_1135),
.B(n_986),
.Y(n_1377)
);

AOI221xp5_ASAP7_75t_L g1378 ( 
.A1(n_1240),
.A2(n_1065),
.B1(n_403),
.B2(n_406),
.C(n_399),
.Y(n_1378)
);

AOI21xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1224),
.A2(n_1133),
.B(n_1034),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1267),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1200),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1207),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1207),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1224),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1309),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_SL g1386 ( 
.A(n_1303),
.B(n_1092),
.C(n_1249),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1264),
.A2(n_1131),
.B1(n_1094),
.B2(n_1028),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1168),
.A2(n_1120),
.B(n_1125),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1227),
.A2(n_1120),
.B(n_1125),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1267),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1189),
.B(n_1050),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1176),
.A2(n_1128),
.B(n_1127),
.Y(n_1392)
);

BUFx4f_ASAP7_75t_L g1393 ( 
.A(n_1180),
.Y(n_1393)
);

BUFx5_ASAP7_75t_L g1394 ( 
.A(n_1279),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1276),
.B(n_1291),
.Y(n_1395)
);

NAND2x1p5_ASAP7_75t_L g1396 ( 
.A(n_1184),
.B(n_1050),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1176),
.A2(n_1128),
.B(n_1127),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1199),
.B(n_1131),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1167),
.A2(n_986),
.B(n_1109),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_SL g1400 ( 
.A1(n_1179),
.A2(n_1072),
.B(n_1143),
.C(n_1111),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1277),
.A2(n_1128),
.B(n_1099),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1169),
.A2(n_998),
.B(n_1146),
.C(n_1139),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1279),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1159),
.B(n_984),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1245),
.A2(n_1134),
.B(n_1143),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1311),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1208),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1159),
.B(n_1059),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1153),
.A2(n_1134),
.A3(n_1111),
.B(n_1141),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1311),
.Y(n_1410)
);

BUFx4f_ASAP7_75t_SL g1411 ( 
.A(n_1217),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1190),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_SL g1413 ( 
.A1(n_1300),
.A2(n_1099),
.B(n_1112),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1277),
.A2(n_1112),
.B(n_1141),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1188),
.A2(n_1027),
.B(n_1010),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1213),
.B(n_1121),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1272),
.A2(n_986),
.B(n_1010),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1184),
.B(n_1062),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1231),
.A2(n_1209),
.B1(n_1249),
.B2(n_1190),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1162),
.A2(n_998),
.B(n_1139),
.C(n_1010),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1208),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1234),
.B(n_1050),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1184),
.B(n_1062),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1298),
.A2(n_1050),
.B1(n_1034),
.B2(n_998),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1247),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1253),
.A2(n_1027),
.B(n_1137),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1290),
.A2(n_1140),
.B(n_1121),
.C(n_1105),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1264),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1247),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1298),
.A2(n_1210),
.B1(n_1180),
.B2(n_1293),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1239),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1239),
.B(n_1130),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1232),
.A2(n_1027),
.B(n_1055),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1232),
.A2(n_975),
.B(n_1097),
.Y(n_1434)
);

BUFx4_ASAP7_75t_SL g1435 ( 
.A(n_1278),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1287),
.A2(n_1097),
.B(n_1105),
.Y(n_1436)
);

AOI32xp33_ASAP7_75t_L g1437 ( 
.A1(n_1164),
.A2(n_400),
.A3(n_408),
.B1(n_411),
.B2(n_409),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1273),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1184),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1266),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1273),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1234),
.B(n_1034),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1287),
.A2(n_1097),
.B(n_1105),
.Y(n_1443)
);

NAND2x1p5_ASAP7_75t_L g1444 ( 
.A(n_1238),
.B(n_1051),
.Y(n_1444)
);

AO32x2_ASAP7_75t_L g1445 ( 
.A1(n_1235),
.A2(n_1003),
.A3(n_1044),
.B1(n_1142),
.B2(n_1037),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1309),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1294),
.A2(n_1037),
.B(n_1074),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1238),
.B(n_988),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1285),
.A2(n_1074),
.B(n_1051),
.C(n_988),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1273),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1294),
.A2(n_1074),
.B(n_1051),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1273),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1280),
.A2(n_1074),
.B(n_1051),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1193),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1160),
.A2(n_988),
.B(n_1018),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1280),
.A2(n_1051),
.B(n_1074),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1228),
.A2(n_1018),
.B(n_1044),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1193),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1269),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1193),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1269),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_SL g1462 ( 
.A1(n_1305),
.A2(n_1296),
.B(n_1153),
.Y(n_1462)
);

AOI21xp33_ASAP7_75t_L g1463 ( 
.A1(n_1248),
.A2(n_1018),
.B(n_1028),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1193),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1259),
.A2(n_410),
.B1(n_987),
.B2(n_1042),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1269),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1269),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1171),
.A2(n_374),
.B1(n_412),
.B2(n_1042),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1238),
.B(n_977),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1226),
.A2(n_1149),
.B(n_1124),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1170),
.A2(n_1042),
.B(n_1021),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1269),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1156),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_SL g1474 ( 
.A1(n_1211),
.A2(n_1042),
.B(n_1021),
.C(n_987),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1260),
.B(n_1042),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1165),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1306),
.A2(n_1021),
.B(n_987),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1306),
.A2(n_1021),
.B(n_987),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1177),
.A2(n_1021),
.B(n_987),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1268),
.B(n_977),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_SL g1481 ( 
.A1(n_1236),
.A2(n_977),
.B(n_157),
.C(n_156),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1198),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1308),
.A2(n_977),
.B(n_14),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1308),
.B(n_151),
.Y(n_1484)
);

AOI222xp33_ASAP7_75t_L g1485 ( 
.A1(n_1312),
.A2(n_374),
.B1(n_412),
.B2(n_1240),
.C1(n_1164),
.C2(n_1310),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1343),
.B(n_1284),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1470),
.A2(n_1393),
.B1(n_1164),
.B2(n_1385),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1343),
.B(n_1284),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_SL g1489 ( 
.A(n_1385),
.B(n_1220),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1393),
.B(n_1220),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1393),
.B(n_1220),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1313),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1338),
.A2(n_1186),
.B(n_1157),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1313),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1325),
.B(n_1266),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_SL g1496 ( 
.A(n_1384),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1419),
.A2(n_1265),
.B1(n_1302),
.B2(n_1301),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1369),
.A2(n_1191),
.B1(n_1164),
.B2(n_1270),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1439),
.B(n_1246),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1372),
.Y(n_1500)
);

OR2x6_ASAP7_75t_L g1501 ( 
.A(n_1314),
.B(n_1296),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1432),
.A2(n_1327),
.B1(n_1344),
.B2(n_1386),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1333),
.A2(n_1292),
.B1(n_1286),
.B2(n_1242),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1374),
.B(n_1171),
.Y(n_1504)
);

AOI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1437),
.A2(n_1218),
.B1(n_1158),
.B2(n_1305),
.C(n_1172),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1318),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1322),
.B(n_1152),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1318),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_SL g1509 ( 
.A(n_1384),
.B(n_1286),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1372),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1435),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1322),
.B(n_1172),
.Y(n_1512)
);

NAND2x1_ASAP7_75t_L g1513 ( 
.A(n_1439),
.B(n_1314),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1320),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1345),
.B(n_1229),
.Y(n_1515)
);

OAI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1341),
.A2(n_1183),
.B1(n_1307),
.B2(n_1297),
.C(n_1241),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1357),
.A2(n_1202),
.B1(n_1178),
.B2(n_1244),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1420),
.A2(n_1204),
.B(n_1233),
.Y(n_1518)
);

INVxp33_ASAP7_75t_L g1519 ( 
.A(n_1395),
.Y(n_1519)
);

CKINVDCx14_ASAP7_75t_R g1520 ( 
.A(n_1446),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1320),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1446),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1428),
.A2(n_1255),
.B1(n_1186),
.B2(n_1221),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_SL g1524 ( 
.A1(n_1373),
.A2(n_1370),
.B(n_1462),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1343),
.B(n_1255),
.Y(n_1525)
);

OAI211xp5_ASAP7_75t_L g1526 ( 
.A1(n_1378),
.A2(n_1283),
.B(n_1282),
.C(n_1194),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1482),
.B(n_1152),
.Y(n_1527)
);

AOI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1430),
.A2(n_1175),
.B(n_1155),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1347),
.Y(n_1529)
);

CKINVDCx11_ASAP7_75t_R g1530 ( 
.A(n_1428),
.Y(n_1530)
);

CKINVDCx6p67_ASAP7_75t_R g1531 ( 
.A(n_1440),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1324),
.A2(n_1223),
.B1(n_1155),
.B2(n_1175),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1318),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1374),
.B(n_1229),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1442),
.A2(n_1155),
.B1(n_1175),
.B2(n_1156),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1363),
.Y(n_1536)
);

INVx8_ASAP7_75t_L g1537 ( 
.A(n_1318),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1369),
.A2(n_1155),
.B1(n_1206),
.B2(n_1289),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1316),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1346),
.A2(n_1175),
.B1(n_1243),
.B2(n_1262),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1335),
.B(n_1229),
.Y(n_1541)
);

CKINVDCx8_ASAP7_75t_R g1542 ( 
.A(n_1440),
.Y(n_1542)
);

BUFx4f_ASAP7_75t_L g1543 ( 
.A(n_1335),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1442),
.A2(n_1261),
.B1(n_1271),
.B2(n_1252),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1347),
.Y(n_1545)
);

AND2x6_ASAP7_75t_L g1546 ( 
.A(n_1431),
.B(n_1404),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1331),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1381),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1463),
.A2(n_1256),
.B1(n_1251),
.B2(n_1229),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1321),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1349),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1416),
.A2(n_1229),
.B1(n_1165),
.B2(n_1152),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1412),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1479),
.A2(n_1152),
.B(n_1165),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1411),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1416),
.B(n_1165),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_R g1557 ( 
.A(n_1335),
.B(n_118),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1391),
.B(n_1152),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1431),
.A2(n_1165),
.B1(n_1289),
.B2(n_1228),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1408),
.A2(n_1263),
.B1(n_16),
.B2(n_18),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1336),
.A2(n_1263),
.B(n_146),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1408),
.A2(n_12),
.B1(n_18),
.B2(n_19),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1321),
.B(n_12),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1331),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1326),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_L g1566 ( 
.A(n_1360),
.B(n_20),
.C(n_22),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1354),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1337),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1398),
.Y(n_1569)
);

AO221x2_ASAP7_75t_L g1570 ( 
.A1(n_1375),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1354),
.B(n_23),
.Y(n_1571)
);

INVx6_ASAP7_75t_L g1572 ( 
.A(n_1354),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1399),
.A2(n_142),
.B(n_27),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1408),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_1574)
);

AND2x6_ASAP7_75t_L g1575 ( 
.A(n_1404),
.B(n_28),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1422),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1404),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_SL g1578 ( 
.A(n_1480),
.B(n_1439),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1422),
.A2(n_34),
.B1(n_44),
.B2(n_46),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1387),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1328),
.B(n_1424),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1371),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1381),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1468),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.C(n_56),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1418),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1482),
.B(n_56),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1448),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1339),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1371),
.B(n_59),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1475),
.B(n_59),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1449),
.A2(n_60),
.B(n_62),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1402),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.C(n_66),
.Y(n_1592)
);

INVx4_ASAP7_75t_SL g1593 ( 
.A(n_1469),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1368),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1594)
);

OR2x6_ASAP7_75t_L g1595 ( 
.A(n_1480),
.B(n_68),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1351),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1418),
.B(n_72),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1370),
.A2(n_108),
.B1(n_75),
.B2(n_76),
.Y(n_1598)
);

CKINVDCx11_ASAP7_75t_R g1599 ( 
.A(n_1418),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1366),
.Y(n_1600)
);

OAI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1465),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.C(n_79),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1483),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1366),
.B(n_82),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1340),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1379),
.A2(n_85),
.B1(n_87),
.B2(n_89),
.C(n_91),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1405),
.A2(n_108),
.B(n_94),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1382),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1340),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1350),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1334),
.A2(n_98),
.B(n_99),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1334),
.A2(n_98),
.B(n_101),
.Y(n_1611)
);

OR2x6_ASAP7_75t_SL g1612 ( 
.A(n_1350),
.B(n_101),
.Y(n_1612)
);

OAI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1480),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1352),
.B(n_106),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1352),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1421),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1366),
.A2(n_1367),
.B1(n_1455),
.B2(n_1377),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1448),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1355),
.A2(n_1403),
.B1(n_1380),
.B2(n_1358),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1367),
.B(n_1356),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1427),
.A2(n_1400),
.B(n_1481),
.C(n_1413),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1358),
.A2(n_1410),
.B1(n_1390),
.B2(n_1406),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1423),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1423),
.Y(n_1625)
);

INVxp33_ASAP7_75t_L g1626 ( 
.A(n_1367),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1405),
.A2(n_1417),
.B(n_1480),
.Y(n_1627)
);

OAI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1484),
.A2(n_1380),
.B1(n_1406),
.B2(n_1403),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1423),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1390),
.B(n_1410),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1421),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1448),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1434),
.A2(n_1353),
.B(n_1361),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1425),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1425),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1396),
.A2(n_1476),
.B1(n_1429),
.B2(n_1466),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1396),
.A2(n_1476),
.B1(n_1429),
.B2(n_1466),
.Y(n_1637)
);

OAI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1444),
.A2(n_1396),
.B1(n_1484),
.B2(n_1436),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1469),
.Y(n_1639)
);

AO31x2_ASAP7_75t_L g1640 ( 
.A1(n_1472),
.A2(n_1459),
.A3(n_1467),
.B(n_1461),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1382),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1383),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_SL g1643 ( 
.A1(n_1473),
.A2(n_1461),
.B(n_1459),
.C(n_1467),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1383),
.B(n_1407),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1407),
.Y(n_1645)
);

OAI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1444),
.A2(n_1484),
.B1(n_1443),
.B2(n_1436),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1436),
.A2(n_1443),
.B1(n_1444),
.B2(n_1472),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1394),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1462),
.A2(n_1443),
.B1(n_1436),
.B2(n_1455),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1394),
.B(n_1469),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1455),
.A2(n_1443),
.B1(n_1394),
.B2(n_1413),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1409),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1330),
.A2(n_1342),
.B1(n_1438),
.B2(n_1441),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1445),
.B(n_1394),
.Y(n_1654)
);

OR2x6_ASAP7_75t_L g1655 ( 
.A(n_1453),
.B(n_1456),
.Y(n_1655)
);

OR2x6_ASAP7_75t_L g1656 ( 
.A(n_1453),
.B(n_1456),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1330),
.A2(n_1342),
.B1(n_1438),
.B2(n_1441),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_SL g1658 ( 
.A1(n_1483),
.A2(n_1394),
.B1(n_1405),
.B2(n_1434),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1353),
.A2(n_1361),
.B(n_1348),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1474),
.A2(n_1452),
.B1(n_1450),
.B2(n_1460),
.C(n_1458),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1473),
.B(n_1471),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1394),
.A2(n_1473),
.B1(n_1483),
.B2(n_1478),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1394),
.B(n_1452),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1483),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1570),
.A2(n_1394),
.B1(n_1342),
.B2(n_1330),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1512),
.B(n_1450),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1504),
.B(n_1409),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1503),
.A2(n_1478),
.B1(n_1477),
.B2(n_1342),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1492),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1502),
.B(n_1409),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1639),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1616),
.A2(n_1478),
.B1(n_1477),
.B2(n_1330),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1573),
.A2(n_1451),
.B(n_1447),
.C(n_1471),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1515),
.B(n_1409),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1570),
.A2(n_1364),
.B1(n_1464),
.B2(n_1454),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1573),
.A2(n_1451),
.B(n_1447),
.C(n_1415),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_SL g1677 ( 
.A(n_1581),
.B(n_1464),
.Y(n_1677)
);

OAI211xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1605),
.A2(n_1454),
.B(n_1460),
.C(n_1458),
.Y(n_1678)
);

AO22x1_ASAP7_75t_L g1679 ( 
.A1(n_1575),
.A2(n_1445),
.B1(n_1409),
.B2(n_1478),
.Y(n_1679)
);

AOI222xp33_ASAP7_75t_L g1680 ( 
.A1(n_1584),
.A2(n_1329),
.B1(n_1332),
.B2(n_1426),
.C1(n_1348),
.C2(n_1445),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1485),
.A2(n_1364),
.B1(n_1457),
.B2(n_1329),
.Y(n_1681)
);

BUFx12f_ASAP7_75t_L g1682 ( 
.A(n_1555),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1494),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1510),
.Y(n_1684)
);

OAI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1557),
.A2(n_1592),
.B1(n_1601),
.B2(n_1595),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1534),
.B(n_1445),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1497),
.A2(n_1477),
.B1(n_1457),
.B2(n_1364),
.Y(n_1687)
);

AOI21xp33_ASAP7_75t_L g1688 ( 
.A1(n_1485),
.A2(n_1457),
.B(n_1477),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1571),
.B(n_1445),
.Y(n_1689)
);

OAI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1595),
.A2(n_1364),
.B1(n_1359),
.B2(n_1332),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1487),
.A2(n_1359),
.B1(n_1426),
.B2(n_1323),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1593),
.B(n_1362),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1495),
.A2(n_1415),
.B1(n_1362),
.B2(n_1392),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1640),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1566),
.A2(n_1433),
.B1(n_1389),
.B2(n_1392),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1540),
.A2(n_1397),
.B1(n_1323),
.B2(n_1359),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1567),
.B(n_1365),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1596),
.A2(n_1359),
.B1(n_1433),
.B2(n_1388),
.C(n_1376),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1659),
.A2(n_1388),
.B(n_1376),
.Y(n_1699)
);

OAI211xp5_ASAP7_75t_L g1700 ( 
.A1(n_1562),
.A2(n_1397),
.B(n_1365),
.C(n_1389),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1613),
.A2(n_1319),
.B1(n_1317),
.B2(n_1315),
.C(n_1414),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1591),
.A2(n_1561),
.B(n_1516),
.C(n_1622),
.Y(n_1702)
);

AO31x2_ASAP7_75t_L g1703 ( 
.A1(n_1538),
.A2(n_1401),
.A3(n_1319),
.B(n_1317),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1519),
.B(n_1568),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1574),
.A2(n_1315),
.B1(n_1401),
.B2(n_1414),
.C(n_1577),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1663),
.Y(n_1706)
);

AOI21xp33_ASAP7_75t_L g1707 ( 
.A1(n_1526),
.A2(n_1517),
.B(n_1561),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1553),
.B(n_1586),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1582),
.A2(n_1602),
.B1(n_1576),
.B2(n_1579),
.Y(n_1709)
);

AOI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1513),
.A2(n_1538),
.B(n_1606),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1599),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1507),
.B(n_1556),
.Y(n_1712)
);

BUFx12f_ASAP7_75t_L g1713 ( 
.A(n_1522),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1582),
.A2(n_1579),
.B1(n_1576),
.B2(n_1609),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1580),
.A2(n_1542),
.B1(n_1595),
.B2(n_1531),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1621),
.B(n_1541),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1565),
.A2(n_1543),
.B1(n_1569),
.B2(n_1496),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1507),
.B(n_1590),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_SL g1720 ( 
.A1(n_1575),
.A2(n_1594),
.B1(n_1489),
.B2(n_1609),
.Y(n_1720)
);

OR2x6_ASAP7_75t_L g1721 ( 
.A(n_1501),
.B(n_1524),
.Y(n_1721)
);

BUFx4f_ASAP7_75t_SL g1722 ( 
.A(n_1551),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1575),
.A2(n_1594),
.B1(n_1563),
.B2(n_1541),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1489),
.A2(n_1491),
.B1(n_1490),
.B2(n_1509),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1575),
.A2(n_1509),
.B1(n_1597),
.B2(n_1546),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1505),
.A2(n_1598),
.B1(n_1560),
.B2(n_1528),
.C(n_1589),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1586),
.A2(n_1597),
.B1(n_1530),
.B2(n_1520),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1614),
.A2(n_1498),
.B1(n_1572),
.B2(n_1603),
.Y(n_1728)
);

NAND4xp25_ASAP7_75t_L g1729 ( 
.A(n_1552),
.B(n_1536),
.C(n_1558),
.D(n_1527),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1498),
.A2(n_1572),
.B1(n_1543),
.B2(n_1486),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1523),
.A2(n_1510),
.B1(n_1521),
.B2(n_1617),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1486),
.A2(n_1488),
.B1(n_1532),
.B2(n_1528),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1514),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1539),
.Y(n_1735)
);

AOI222xp33_ASAP7_75t_L g1736 ( 
.A1(n_1612),
.A2(n_1488),
.B1(n_1518),
.B2(n_1626),
.C1(n_1525),
.C2(n_1587),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1550),
.A2(n_1527),
.B1(n_1500),
.B2(n_1632),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1627),
.A2(n_1554),
.B(n_1518),
.Y(n_1738)
);

OAI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1500),
.A2(n_1619),
.B1(n_1618),
.B2(n_1501),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1525),
.A2(n_1500),
.B1(n_1585),
.B2(n_1499),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1546),
.A2(n_1624),
.B1(n_1625),
.B2(n_1639),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1585),
.A2(n_1499),
.B1(n_1651),
.B2(n_1629),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1547),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1629),
.A2(n_1501),
.B1(n_1625),
.B2(n_1624),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1639),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1546),
.A2(n_1631),
.B1(n_1635),
.B2(n_1634),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1578),
.A2(n_1638),
.B(n_1650),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1546),
.A2(n_1628),
.B1(n_1654),
.B2(n_1610),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1636),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1537),
.B(n_1637),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1564),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1549),
.A2(n_1544),
.B(n_1559),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1649),
.A2(n_1664),
.B(n_1658),
.C(n_1511),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1619),
.A2(n_1535),
.B1(n_1588),
.B2(n_1615),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1646),
.A2(n_1662),
.B(n_1643),
.Y(n_1755)
);

AOI222xp33_ASAP7_75t_L g1756 ( 
.A1(n_1604),
.A2(n_1608),
.B1(n_1620),
.B2(n_1623),
.C1(n_1630),
.C2(n_1641),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1648),
.A2(n_1636),
.B1(n_1637),
.B2(n_1647),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1611),
.A2(n_1642),
.B1(n_1645),
.B2(n_1529),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1537),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1545),
.B(n_1548),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1633),
.A2(n_1660),
.B(n_1661),
.C(n_1537),
.Y(n_1761)
);

AOI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1647),
.A2(n_1652),
.B1(n_1653),
.B2(n_1657),
.C(n_1633),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1583),
.A2(n_1607),
.B1(n_1644),
.B2(n_1533),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1506),
.B(n_1508),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1653),
.B(n_1657),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1508),
.A2(n_1533),
.B1(n_1661),
.B2(n_1659),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1655),
.A2(n_1656),
.B1(n_990),
.B2(n_1312),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1655),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1655),
.A2(n_1570),
.B1(n_1485),
.B2(n_1161),
.Y(n_1769)
);

BUFx4f_ASAP7_75t_SL g1770 ( 
.A(n_1656),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1656),
.B(n_1026),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1659),
.A2(n_1633),
.B(n_1554),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1570),
.A2(n_1485),
.B1(n_1161),
.B2(n_1592),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1566),
.B(n_1386),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_SL g1775 ( 
.A1(n_1570),
.A2(n_990),
.B1(n_1026),
.B2(n_1592),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1570),
.A2(n_1485),
.B1(n_1161),
.B2(n_1592),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1503),
.A2(n_990),
.B1(n_1312),
.B2(n_1026),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1503),
.A2(n_990),
.B1(n_1312),
.B2(n_1026),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1570),
.A2(n_1485),
.B1(n_1161),
.B2(n_1592),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1504),
.B(n_1534),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_SL g1781 ( 
.A1(n_1570),
.A2(n_990),
.B1(n_1026),
.B2(n_1592),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1504),
.B(n_1534),
.Y(n_1782)
);

AOI222xp33_ASAP7_75t_L g1783 ( 
.A1(n_1573),
.A2(n_876),
.B1(n_1161),
.B2(n_990),
.C1(n_1026),
.C2(n_1584),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1503),
.A2(n_990),
.B1(n_1312),
.B2(n_1026),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1570),
.A2(n_1161),
.B1(n_990),
.B2(n_1026),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1510),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1515),
.B(n_1534),
.Y(n_1787)
);

AOI222xp33_ASAP7_75t_L g1788 ( 
.A1(n_1573),
.A2(n_876),
.B1(n_1161),
.B2(n_990),
.C1(n_1026),
.C2(n_1584),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1504),
.B(n_1534),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1570),
.A2(n_990),
.B1(n_1026),
.B2(n_1592),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1570),
.A2(n_1161),
.B1(n_990),
.B2(n_1026),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1592),
.A2(n_990),
.B1(n_1026),
.B2(n_1254),
.C(n_722),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1503),
.A2(n_990),
.B1(n_1312),
.B2(n_1026),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1573),
.A2(n_1026),
.B1(n_990),
.B2(n_864),
.C(n_1254),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1503),
.A2(n_990),
.B1(n_1312),
.B2(n_1026),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1510),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1512),
.B(n_1026),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1570),
.A2(n_1485),
.B1(n_1161),
.B2(n_1592),
.Y(n_1798)
);

AND2x4_ASAP7_75t_SL g1799 ( 
.A(n_1500),
.B(n_1220),
.Y(n_1799)
);

INVxp33_ASAP7_75t_SL g1800 ( 
.A(n_1522),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1515),
.B(n_1534),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1599),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1570),
.A2(n_1161),
.B1(n_990),
.B2(n_1026),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1570),
.A2(n_1161),
.B1(n_990),
.B2(n_1026),
.Y(n_1804)
);

INVx4_ASAP7_75t_L g1805 ( 
.A(n_1500),
.Y(n_1805)
);

OAI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1557),
.A2(n_1592),
.B1(n_1601),
.B2(n_1573),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1493),
.A2(n_1338),
.B(n_1314),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1570),
.A2(n_1485),
.B1(n_1161),
.B2(n_1592),
.Y(n_1809)
);

OAI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1557),
.A2(n_1592),
.B1(n_1601),
.B2(n_1573),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1503),
.A2(n_990),
.B1(n_1026),
.B2(n_789),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1573),
.A2(n_1026),
.B1(n_990),
.B2(n_864),
.C(n_1254),
.Y(n_1812)
);

OAI21xp33_ASAP7_75t_L g1813 ( 
.A1(n_1573),
.A2(n_990),
.B(n_1026),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1570),
.A2(n_1485),
.B1(n_1161),
.B2(n_1592),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_L g1815 ( 
.A(n_1566),
.B(n_1026),
.C(n_990),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1573),
.A2(n_1026),
.B(n_990),
.C(n_1161),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1592),
.A2(n_536),
.B1(n_1026),
.B2(n_990),
.C(n_707),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1492),
.Y(n_1818)
);

AOI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1592),
.A2(n_536),
.B1(n_1026),
.B2(n_990),
.C(n_707),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1694),
.Y(n_1820)
);

OAI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1816),
.A2(n_1815),
.B(n_1812),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1794),
.A2(n_1813),
.B(n_1811),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1686),
.B(n_1712),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1706),
.B(n_1719),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1703),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1689),
.B(n_1787),
.Y(n_1826)
);

AOI33xp33_ASAP7_75t_L g1827 ( 
.A1(n_1785),
.A2(n_1804),
.A3(n_1791),
.B1(n_1803),
.B2(n_1773),
.B3(n_1809),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1692),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1801),
.B(n_1780),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1703),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1782),
.B(n_1789),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1749),
.B(n_1667),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1768),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1699),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1770),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1735),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1703),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1773),
.A2(n_1779),
.B1(n_1776),
.B2(n_1814),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1749),
.B(n_1765),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1734),
.Y(n_1840)
);

AOI21x1_ASAP7_75t_L g1841 ( 
.A1(n_1679),
.A2(n_1771),
.B(n_1755),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1743),
.B(n_1751),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1669),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1704),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1684),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1721),
.B(n_1750),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1721),
.B(n_1750),
.Y(n_1847)
);

INVx3_ASAP7_75t_SL g1848 ( 
.A(n_1799),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_1683),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1708),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1770),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1800),
.B(n_1777),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1721),
.B(n_1750),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1818),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1674),
.B(n_1717),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1757),
.B(n_1762),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1738),
.B(n_1729),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1754),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1703),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1772),
.Y(n_1860)
);

OR2x6_ASAP7_75t_L g1861 ( 
.A(n_1808),
.B(n_1747),
.Y(n_1861)
);

BUFx12f_ASAP7_75t_L g1862 ( 
.A(n_1713),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1697),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1666),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1670),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1665),
.B(n_1675),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1772),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1690),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1690),
.Y(n_1869)
);

AOI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1776),
.A2(n_1809),
.B1(n_1798),
.B2(n_1814),
.C(n_1779),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1665),
.B(n_1675),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1702),
.A2(n_1788),
.B(n_1783),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1672),
.B(n_1772),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1761),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1798),
.A2(n_1795),
.B1(n_1784),
.B2(n_1793),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1760),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1775),
.A2(n_1790),
.B1(n_1781),
.B2(n_1709),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1687),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1668),
.B(n_1767),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1710),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1733),
.B(n_1748),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1733),
.B(n_1752),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1693),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1698),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1696),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1766),
.B(n_1673),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1691),
.B(n_1677),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1756),
.B(n_1797),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1744),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1705),
.Y(n_1890)
);

INVx5_ASAP7_75t_L g1891 ( 
.A(n_1714),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1676),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1681),
.B(n_1766),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1681),
.B(n_1736),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1786),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1688),
.B(n_1746),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1746),
.B(n_1728),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1728),
.B(n_1731),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1709),
.A2(n_1769),
.B1(n_1792),
.B2(n_1715),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1731),
.B(n_1769),
.Y(n_1900)
);

AOI33xp33_ASAP7_75t_L g1901 ( 
.A1(n_1817),
.A2(n_1819),
.A3(n_1715),
.B1(n_1810),
.B2(n_1806),
.B3(n_1720),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1732),
.B(n_1737),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1758),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1758),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1739),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1739),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1730),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1737),
.B(n_1742),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1680),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1701),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1707),
.B(n_1774),
.Y(n_1911)
);

OAI211xp5_ASAP7_75t_L g1912 ( 
.A1(n_1778),
.A2(n_1726),
.B(n_1723),
.C(n_1753),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1805),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1868),
.B(n_1700),
.Y(n_1914)
);

AOI33xp33_ASAP7_75t_L g1915 ( 
.A1(n_1838),
.A2(n_1810),
.A3(n_1806),
.B1(n_1685),
.B2(n_1727),
.B3(n_1725),
.Y(n_1915)
);

AO21x2_ASAP7_75t_L g1916 ( 
.A1(n_1880),
.A2(n_1830),
.B(n_1825),
.Y(n_1916)
);

OAI33xp33_ASAP7_75t_L g1917 ( 
.A1(n_1877),
.A2(n_1685),
.A3(n_1716),
.B1(n_1678),
.B2(n_1718),
.B3(n_1740),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1877),
.A2(n_1727),
.B1(n_1763),
.B2(n_1796),
.C(n_1724),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1872),
.A2(n_1763),
.B1(n_1802),
.B2(n_1711),
.C(n_1671),
.Y(n_1919)
);

AOI31xp33_ASAP7_75t_L g1920 ( 
.A1(n_1872),
.A2(n_1741),
.A3(n_1764),
.B(n_1807),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1850),
.Y(n_1921)
);

OAI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1821),
.A2(n_1711),
.B1(n_1802),
.B2(n_1671),
.C(n_1805),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1836),
.Y(n_1923)
);

OAI211xp5_ASAP7_75t_L g1924 ( 
.A1(n_1875),
.A2(n_1870),
.B(n_1821),
.C(n_1912),
.Y(n_1924)
);

OAI322xp33_ASAP7_75t_L g1925 ( 
.A1(n_1875),
.A2(n_1711),
.A3(n_1802),
.B1(n_1745),
.B2(n_1759),
.C1(n_1722),
.C2(n_1695),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1824),
.B(n_1807),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1828),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1868),
.B(n_1711),
.Y(n_1928)
);

INVx4_ASAP7_75t_L g1929 ( 
.A(n_1848),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1824),
.B(n_1745),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1870),
.A2(n_1802),
.B1(n_1745),
.B2(n_1722),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1862),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1891),
.Y(n_1933)
);

OAI211xp5_ASAP7_75t_L g1934 ( 
.A1(n_1822),
.A2(n_1682),
.B(n_1745),
.C(n_1911),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1822),
.A2(n_1899),
.B1(n_1874),
.B2(n_1911),
.C(n_1857),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1862),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1899),
.A2(n_1874),
.B1(n_1856),
.B2(n_1882),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1823),
.B(n_1826),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1882),
.A2(n_1856),
.B1(n_1881),
.B2(n_1894),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1828),
.Y(n_1940)
);

INVxp67_ASAP7_75t_L g1941 ( 
.A(n_1864),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1823),
.B(n_1826),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1881),
.A2(n_1894),
.B1(n_1900),
.B2(n_1909),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1843),
.Y(n_1944)
);

BUFx12f_ASAP7_75t_L g1945 ( 
.A(n_1862),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1854),
.Y(n_1946)
);

OAI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1857),
.A2(n_1888),
.B1(n_1909),
.B2(n_1852),
.C(n_1861),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1832),
.B(n_1839),
.Y(n_1948)
);

OAI211xp5_ASAP7_75t_L g1949 ( 
.A1(n_1910),
.A2(n_1888),
.B(n_1883),
.C(n_1885),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1829),
.B(n_1855),
.Y(n_1950)
);

AOI32xp33_ASAP7_75t_L g1951 ( 
.A1(n_1900),
.A2(n_1866),
.A3(n_1871),
.B1(n_1897),
.B2(n_1898),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1902),
.A2(n_1906),
.B1(n_1908),
.B2(n_1898),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1849),
.Y(n_1953)
);

AOI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1910),
.A2(n_1883),
.B1(n_1885),
.B2(n_1878),
.C(n_1858),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1833),
.Y(n_1955)
);

OR2x6_ASAP7_75t_L g1956 ( 
.A(n_1861),
.B(n_1846),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1902),
.A2(n_1906),
.B1(n_1908),
.B2(n_1897),
.Y(n_1957)
);

OR2x6_ASAP7_75t_L g1958 ( 
.A(n_1861),
.B(n_1846),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1876),
.Y(n_1959)
);

BUFx3_ASAP7_75t_L g1960 ( 
.A(n_1848),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1845),
.A2(n_1895),
.B1(n_1840),
.B2(n_1905),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1869),
.B(n_1878),
.Y(n_1962)
);

AOI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1866),
.A2(n_1871),
.B1(n_1890),
.B2(n_1893),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1820),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1832),
.B(n_1839),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1833),
.Y(n_1966)
);

OR2x6_ASAP7_75t_L g1967 ( 
.A(n_1861),
.B(n_1846),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1844),
.B(n_1848),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1863),
.B(n_1855),
.Y(n_1969)
);

NAND4xp25_ASAP7_75t_L g1970 ( 
.A(n_1901),
.B(n_1827),
.C(n_1869),
.D(n_1858),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1829),
.B(n_1876),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1891),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1890),
.A2(n_1893),
.B1(n_1886),
.B2(n_1905),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1863),
.Y(n_1974)
);

INVx5_ASAP7_75t_SL g1975 ( 
.A(n_1861),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1879),
.A2(n_1890),
.B1(n_1886),
.B2(n_1851),
.Y(n_1976)
);

AOI31xp33_ASAP7_75t_SL g1977 ( 
.A1(n_1879),
.A2(n_1887),
.A3(n_1884),
.B(n_1889),
.Y(n_1977)
);

INVxp67_ASAP7_75t_L g1978 ( 
.A(n_1842),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1849),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1896),
.A2(n_1886),
.B1(n_1853),
.B2(n_1847),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1884),
.A2(n_1896),
.B(n_1892),
.Y(n_1981)
);

NOR2x2_ASAP7_75t_L g1982 ( 
.A(n_1907),
.B(n_1889),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1886),
.A2(n_1851),
.B1(n_1835),
.B2(n_1887),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1916),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1923),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1916),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1923),
.Y(n_1987)
);

INVxp33_ASAP7_75t_L g1988 ( 
.A(n_1935),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1964),
.Y(n_1989)
);

AND4x1_ASAP7_75t_L g1990 ( 
.A(n_1915),
.B(n_1892),
.C(n_1873),
.D(n_1904),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1964),
.Y(n_1991)
);

INVxp67_ASAP7_75t_SL g1992 ( 
.A(n_1962),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1933),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1933),
.B(n_1834),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1938),
.B(n_1860),
.Y(n_1995)
);

AND2x4_ASAP7_75t_SL g1996 ( 
.A(n_1956),
.B(n_1853),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1962),
.B(n_1865),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1956),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1942),
.B(n_1867),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1956),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1969),
.B(n_1837),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1956),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1969),
.B(n_1837),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1944),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1946),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1947),
.B(n_1831),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1959),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1958),
.B(n_1859),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1927),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1955),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1982),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1927),
.Y(n_2012)
);

AND2x4_ASAP7_75t_SL g2013 ( 
.A(n_1958),
.B(n_1853),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1940),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1982),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1958),
.B(n_1967),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1914),
.B(n_1837),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1951),
.B(n_1891),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1914),
.B(n_1859),
.Y(n_2019)
);

NAND2x1p5_ASAP7_75t_L g2020 ( 
.A(n_1972),
.B(n_1891),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1940),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1953),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1979),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1978),
.Y(n_2024)
);

INVx4_ASAP7_75t_L g2025 ( 
.A(n_1958),
.Y(n_2025)
);

NOR2x1_ASAP7_75t_L g2026 ( 
.A(n_1977),
.B(n_1820),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1967),
.B(n_1825),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1967),
.B(n_1825),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1972),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1967),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1991),
.Y(n_2031)
);

INVxp67_ASAP7_75t_SL g2032 ( 
.A(n_2026),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2006),
.B(n_1921),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1996),
.B(n_1980),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_2026),
.B(n_1981),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2004),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_2011),
.B(n_2015),
.Y(n_2037)
);

A2O1A1Ixp33_ASAP7_75t_L g2038 ( 
.A1(n_1988),
.A2(n_1924),
.B(n_1915),
.C(n_1937),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1991),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2004),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2011),
.B(n_1948),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1985),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2006),
.B(n_1941),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_1997),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_2011),
.B(n_1966),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1985),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1997),
.B(n_1963),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_2011),
.B(n_1950),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1997),
.B(n_1948),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1985),
.Y(n_2050)
);

OAI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1988),
.A2(n_1949),
.B(n_1939),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2007),
.B(n_1965),
.Y(n_2052)
);

NOR2x1p5_ASAP7_75t_L g2053 ( 
.A(n_2015),
.B(n_1945),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1987),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1987),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2007),
.B(n_1965),
.Y(n_2056)
);

NOR3xp33_ASAP7_75t_L g2057 ( 
.A(n_2018),
.B(n_1934),
.C(n_1917),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2007),
.B(n_1954),
.Y(n_2058)
);

INVx3_ASAP7_75t_L g2059 ( 
.A(n_2020),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1986),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2015),
.B(n_1975),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2024),
.B(n_1930),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_2010),
.Y(n_2063)
);

NOR2x1p5_ASAP7_75t_L g2064 ( 
.A(n_2015),
.B(n_1945),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2024),
.B(n_1926),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_2010),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1987),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2001),
.B(n_1975),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2001),
.B(n_1975),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1989),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2004),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2001),
.B(n_1975),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1989),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1989),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2024),
.B(n_1971),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_2017),
.B(n_1974),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2001),
.B(n_1828),
.Y(n_2077)
);

NAND2xp67_ASAP7_75t_L g2078 ( 
.A(n_2030),
.B(n_1932),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2005),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2005),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2005),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2017),
.B(n_1884),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2005),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2003),
.B(n_1828),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2058),
.B(n_2026),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2042),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_2035),
.A2(n_2018),
.B(n_1920),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_2053),
.B(n_2025),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2061),
.B(n_2016),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_2063),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2061),
.B(n_2016),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2042),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_2037),
.B(n_2017),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2037),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2041),
.B(n_2016),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2041),
.B(n_2064),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_2059),
.B(n_2025),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2047),
.B(n_1943),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_2051),
.B(n_1929),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2068),
.B(n_2016),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2048),
.B(n_2017),
.Y(n_2101)
);

NAND3xp33_ASAP7_75t_L g2102 ( 
.A(n_2038),
.B(n_1990),
.C(n_1970),
.Y(n_2102)
);

NOR4xp25_ASAP7_75t_SL g2103 ( 
.A(n_2032),
.B(n_1922),
.C(n_1992),
.D(n_1919),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_2033),
.B(n_1932),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2046),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_2043),
.B(n_1936),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2046),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2050),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2057),
.B(n_1992),
.Y(n_2109)
);

INVx1_ASAP7_75t_SL g2110 ( 
.A(n_2082),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2068),
.B(n_2030),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2050),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2065),
.B(n_1957),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2054),
.Y(n_2114)
);

BUFx2_ASAP7_75t_L g2115 ( 
.A(n_2066),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2054),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2075),
.B(n_1952),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2082),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2055),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2055),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2067),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2067),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2070),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_2059),
.B(n_2025),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2070),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2048),
.B(n_2019),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2069),
.B(n_2030),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2060),
.Y(n_2128)
);

INVx6_ASAP7_75t_L g2129 ( 
.A(n_2034),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2036),
.Y(n_2130)
);

OR2x4_ASAP7_75t_L g2131 ( 
.A(n_2045),
.B(n_1968),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2040),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2069),
.B(n_2030),
.Y(n_2133)
);

AOI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2102),
.A2(n_2034),
.B1(n_1931),
.B2(n_1976),
.Y(n_2134)
);

AOI21xp33_ASAP7_75t_L g2135 ( 
.A1(n_2102),
.A2(n_2078),
.B(n_1983),
.Y(n_2135)
);

AOI221xp5_ASAP7_75t_L g2136 ( 
.A1(n_2087),
.A2(n_2044),
.B1(n_1925),
.B2(n_1973),
.C(n_1961),
.Y(n_2136)
);

AOI221x1_ASAP7_75t_L g2137 ( 
.A1(n_2109),
.A2(n_1929),
.B1(n_2039),
.B2(n_2031),
.C(n_2022),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2099),
.A2(n_2034),
.B1(n_2025),
.B2(n_1998),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2093),
.Y(n_2139)
);

OAI21xp33_ASAP7_75t_L g2140 ( 
.A1(n_2085),
.A2(n_2098),
.B(n_2096),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_2103),
.A2(n_2131),
.B(n_2113),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2130),
.Y(n_2142)
);

OAI32xp33_ASAP7_75t_L g2143 ( 
.A1(n_2103),
.A2(n_1990),
.A3(n_2045),
.B1(n_1928),
.B2(n_2031),
.Y(n_2143)
);

AOI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_2115),
.A2(n_1918),
.B1(n_2062),
.B2(n_2059),
.C(n_2039),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2115),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2086),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2117),
.B(n_2078),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_2104),
.B(n_1936),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2094),
.B(n_2049),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2096),
.B(n_2072),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_2129),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2086),
.Y(n_2152)
);

INVx1_ASAP7_75t_SL g2153 ( 
.A(n_2088),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2093),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2095),
.Y(n_2155)
);

NOR2x1_ASAP7_75t_L g2156 ( 
.A(n_2088),
.B(n_1960),
.Y(n_2156)
);

O2A1O1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_2090),
.A2(n_1928),
.B(n_1960),
.C(n_1990),
.Y(n_2157)
);

INVx3_ASAP7_75t_SL g2158 ( 
.A(n_2088),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2090),
.B(n_2052),
.Y(n_2159)
);

OAI31xp33_ASAP7_75t_L g2160 ( 
.A1(n_2088),
.A2(n_2002),
.A3(n_2000),
.B(n_1998),
.Y(n_2160)
);

OAI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2131),
.A2(n_2129),
.B1(n_2025),
.B2(n_2002),
.Y(n_2161)
);

AOI322xp5_ASAP7_75t_L g2162 ( 
.A1(n_2106),
.A2(n_2056),
.A3(n_2072),
.B1(n_2084),
.B2(n_2077),
.C1(n_1999),
.C2(n_1995),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2130),
.Y(n_2163)
);

O2A1O1Ixp33_ASAP7_75t_L g2164 ( 
.A1(n_2094),
.A2(n_2020),
.B(n_2000),
.C(n_1998),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_2131),
.B(n_1929),
.Y(n_2165)
);

INVxp67_ASAP7_75t_SL g2166 ( 
.A(n_2089),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2089),
.A2(n_2025),
.B1(n_1998),
.B2(n_2002),
.Y(n_2167)
);

AOI211xp5_ASAP7_75t_SL g2168 ( 
.A1(n_2091),
.A2(n_1835),
.B(n_1998),
.C(n_2002),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2095),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2107),
.Y(n_2170)
);

NAND2xp33_ASAP7_75t_L g2171 ( 
.A(n_2091),
.B(n_2020),
.Y(n_2171)
);

OAI22xp5_ASAP7_75t_L g2172 ( 
.A1(n_2129),
.A2(n_2025),
.B1(n_2002),
.B2(n_2000),
.Y(n_2172)
);

OAI21xp5_ASAP7_75t_SL g2173 ( 
.A1(n_2141),
.A2(n_2100),
.B(n_2133),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2145),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2140),
.B(n_2111),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2166),
.B(n_2110),
.Y(n_2176)
);

AOI222xp33_ASAP7_75t_L g2177 ( 
.A1(n_2143),
.A2(n_2118),
.B1(n_2100),
.B2(n_2111),
.C1(n_2133),
.C2(n_2127),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2136),
.B(n_2127),
.Y(n_2178)
);

AOI32xp33_ASAP7_75t_L g2179 ( 
.A1(n_2156),
.A2(n_2124),
.A3(n_2097),
.B1(n_2002),
.B2(n_2000),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2165),
.A2(n_2129),
.B1(n_2097),
.B2(n_2124),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2146),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2153),
.B(n_2132),
.Y(n_2182)
);

INVx2_ASAP7_75t_SL g2183 ( 
.A(n_2151),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_2135),
.A2(n_1903),
.B1(n_1904),
.B2(n_2124),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_SL g2185 ( 
.A1(n_2134),
.A2(n_2097),
.B(n_2124),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2146),
.Y(n_2186)
);

A2O1A1Ixp33_ASAP7_75t_L g2187 ( 
.A1(n_2143),
.A2(n_1998),
.B(n_2000),
.C(n_1851),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2159),
.B(n_2155),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2144),
.A2(n_2132),
.B1(n_2108),
.B2(n_2119),
.C(n_2125),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2138),
.A2(n_2000),
.B1(n_2020),
.B2(n_1996),
.Y(n_2190)
);

AOI322xp5_ASAP7_75t_L g2191 ( 
.A1(n_2161),
.A2(n_2147),
.A3(n_2150),
.B1(n_2155),
.B2(n_2169),
.C1(n_2151),
.C2(n_2148),
.Y(n_2191)
);

NOR2x1_ASAP7_75t_L g2192 ( 
.A(n_2157),
.B(n_2092),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_2150),
.B(n_2097),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2169),
.B(n_2101),
.Y(n_2194)
);

INVxp33_ASAP7_75t_L g2195 ( 
.A(n_2137),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2139),
.B(n_2101),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2158),
.Y(n_2197)
);

OAI221xp5_ASAP7_75t_L g2198 ( 
.A1(n_2160),
.A2(n_2126),
.B1(n_2020),
.B2(n_2125),
.C(n_2119),
.Y(n_2198)
);

OAI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_2137),
.A2(n_2116),
.B(n_2108),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2152),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2158),
.B(n_2077),
.Y(n_2201)
);

NAND2xp33_ASAP7_75t_SL g2202 ( 
.A(n_2172),
.B(n_2126),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2183),
.B(n_2168),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2181),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_2178),
.B(n_2167),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_2197),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_2179),
.B(n_2164),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2193),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2186),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2195),
.A2(n_2149),
.B1(n_2154),
.B2(n_2139),
.Y(n_2210)
);

INVx3_ASAP7_75t_SL g2211 ( 
.A(n_2174),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2189),
.B(n_2154),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2200),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2196),
.Y(n_2214)
);

AOI22x1_ASAP7_75t_L g2215 ( 
.A1(n_2177),
.A2(n_2142),
.B1(n_2163),
.B2(n_2170),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2189),
.B(n_2162),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_2193),
.Y(n_2217)
);

AOI222xp33_ASAP7_75t_L g2218 ( 
.A1(n_2195),
.A2(n_2171),
.B1(n_2152),
.B2(n_2170),
.C1(n_2116),
.C2(n_2120),
.Y(n_2218)
);

INVx1_ASAP7_75t_SL g2219 ( 
.A(n_2202),
.Y(n_2219)
);

NOR3xp33_ASAP7_75t_SL g2220 ( 
.A(n_2185),
.B(n_2105),
.C(n_2092),
.Y(n_2220)
);

INVxp67_ASAP7_75t_L g2221 ( 
.A(n_2175),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2173),
.B(n_2149),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2201),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2176),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2182),
.Y(n_2225)
);

OR2x2_ASAP7_75t_L g2226 ( 
.A(n_2188),
.B(n_2105),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2212),
.B(n_2184),
.Y(n_2227)
);

NOR2x1_ASAP7_75t_L g2228 ( 
.A(n_2224),
.B(n_2187),
.Y(n_2228)
);

NAND4xp25_ASAP7_75t_L g2229 ( 
.A(n_2205),
.B(n_2191),
.C(n_2180),
.D(n_2187),
.Y(n_2229)
);

NAND4xp75_ASAP7_75t_L g2230 ( 
.A(n_2216),
.B(n_2192),
.C(n_2199),
.D(n_2194),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2211),
.B(n_2184),
.Y(n_2231)
);

AOI211xp5_ASAP7_75t_L g2232 ( 
.A1(n_2219),
.A2(n_2190),
.B(n_2198),
.C(n_2171),
.Y(n_2232)
);

NOR3xp33_ASAP7_75t_L g2233 ( 
.A(n_2206),
.B(n_2221),
.C(n_2224),
.Y(n_2233)
);

NOR4xp25_ASAP7_75t_L g2234 ( 
.A(n_2210),
.B(n_2123),
.C(n_2122),
.D(n_2121),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2204),
.Y(n_2235)
);

NAND4xp75_ASAP7_75t_L g2236 ( 
.A(n_2220),
.B(n_2203),
.C(n_2207),
.D(n_2217),
.Y(n_2236)
);

AOI221x1_ASAP7_75t_L g2237 ( 
.A1(n_2204),
.A2(n_2120),
.B1(n_2123),
.B2(n_2122),
.C(n_2121),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2209),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2209),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_L g2240 ( 
.A(n_2211),
.B(n_2076),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2213),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2217),
.B(n_2112),
.Y(n_2242)
);

OAI211xp5_ASAP7_75t_L g2243 ( 
.A1(n_2228),
.A2(n_2215),
.B(n_2218),
.C(n_2222),
.Y(n_2243)
);

A2O1A1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_2227),
.A2(n_2203),
.B(n_2225),
.C(n_2214),
.Y(n_2244)
);

AOI221xp5_ASAP7_75t_L g2245 ( 
.A1(n_2227),
.A2(n_2225),
.B1(n_2214),
.B2(n_2223),
.C(n_2208),
.Y(n_2245)
);

AOI211xp5_ASAP7_75t_L g2246 ( 
.A1(n_2229),
.A2(n_2208),
.B(n_2223),
.C(n_2213),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2230),
.A2(n_2215),
.B1(n_2226),
.B2(n_2112),
.Y(n_2247)
);

NOR2x1_ASAP7_75t_L g2248 ( 
.A(n_2236),
.B(n_2226),
.Y(n_2248)
);

AOI32xp33_ASAP7_75t_L g2249 ( 
.A1(n_2231),
.A2(n_2128),
.A3(n_2114),
.B1(n_2107),
.B2(n_1993),
.Y(n_2249)
);

AOI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_2233),
.A2(n_1853),
.B1(n_1846),
.B2(n_1847),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2232),
.A2(n_2076),
.B1(n_1993),
.B2(n_2019),
.Y(n_2251)
);

NAND4xp75_ASAP7_75t_L g2252 ( 
.A(n_2240),
.B(n_1993),
.C(n_2128),
.D(n_2114),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2234),
.B(n_2242),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2235),
.B(n_2084),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2238),
.A2(n_1835),
.B1(n_2013),
.B2(n_1996),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2239),
.A2(n_1993),
.B1(n_1835),
.B2(n_2029),
.C(n_2060),
.Y(n_2256)
);

AOI21xp5_ASAP7_75t_L g2257 ( 
.A1(n_2243),
.A2(n_2241),
.B(n_2237),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2248),
.A2(n_2029),
.B(n_2022),
.Y(n_2258)
);

AOI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2251),
.A2(n_2013),
.B1(n_1996),
.B2(n_2027),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_2254),
.Y(n_2260)
);

AOI221xp5_ASAP7_75t_L g2261 ( 
.A1(n_2247),
.A2(n_1984),
.B1(n_2022),
.B2(n_2023),
.C(n_2071),
.Y(n_2261)
);

CKINVDCx20_ASAP7_75t_R g2262 ( 
.A(n_2253),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_2255),
.Y(n_2263)
);

NAND3xp33_ASAP7_75t_L g2264 ( 
.A(n_2246),
.B(n_2244),
.C(n_2245),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2249),
.B(n_2073),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2260),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_2258),
.Y(n_2267)
);

NAND3xp33_ASAP7_75t_L g2268 ( 
.A(n_2264),
.B(n_2250),
.C(n_2256),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2262),
.A2(n_1847),
.B1(n_1996),
.B2(n_2013),
.Y(n_2269)
);

NAND2x1p5_ASAP7_75t_L g2270 ( 
.A(n_2257),
.B(n_2259),
.Y(n_2270)
);

HB1xp67_ASAP7_75t_L g2271 ( 
.A(n_2263),
.Y(n_2271)
);

BUFx3_ASAP7_75t_L g2272 ( 
.A(n_2265),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_2261),
.B(n_2252),
.Y(n_2273)
);

NAND4xp25_ASAP7_75t_L g2274 ( 
.A(n_2268),
.B(n_2266),
.C(n_2272),
.D(n_2273),
.Y(n_2274)
);

INVxp67_ASAP7_75t_SL g2275 ( 
.A(n_2267),
.Y(n_2275)
);

NOR3xp33_ASAP7_75t_L g2276 ( 
.A(n_2271),
.B(n_1841),
.C(n_1913),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2267),
.Y(n_2277)
);

XOR2x2_ASAP7_75t_L g2278 ( 
.A(n_2270),
.B(n_1841),
.Y(n_2278)
);

NAND3x2_ASAP7_75t_L g2279 ( 
.A(n_2273),
.B(n_2019),
.C(n_1994),
.Y(n_2279)
);

NAND5xp2_ASAP7_75t_L g2280 ( 
.A(n_2270),
.B(n_2008),
.C(n_2027),
.D(n_2028),
.E(n_1903),
.Y(n_2280)
);

NOR3xp33_ASAP7_75t_L g2281 ( 
.A(n_2269),
.B(n_1913),
.C(n_2029),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_2275),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_2277),
.Y(n_2283)
);

AOI22xp33_ASAP7_75t_R g2284 ( 
.A1(n_2279),
.A2(n_2029),
.B1(n_2009),
.B2(n_2012),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2274),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_2282),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2282),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2286),
.B(n_2283),
.Y(n_2288)
);

OAI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_2287),
.A2(n_2285),
.B1(n_2284),
.B2(n_2278),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2288),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_2289),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2288),
.A2(n_2281),
.B1(n_2276),
.B2(n_2280),
.Y(n_2292)
);

INVxp33_ASAP7_75t_SL g2293 ( 
.A(n_2291),
.Y(n_2293)
);

AOI222xp33_ASAP7_75t_SL g2294 ( 
.A1(n_2290),
.A2(n_2014),
.B1(n_2021),
.B2(n_2012),
.C1(n_2009),
.C2(n_2083),
.Y(n_2294)
);

AOI222xp33_ASAP7_75t_L g2295 ( 
.A1(n_2293),
.A2(n_2292),
.B1(n_2083),
.B2(n_2081),
.C1(n_2080),
.C2(n_2079),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2294),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2296),
.Y(n_2297)
);

AOI221xp5_ASAP7_75t_L g2298 ( 
.A1(n_2297),
.A2(n_2295),
.B1(n_2081),
.B2(n_2080),
.C(n_2079),
.Y(n_2298)
);

AOI211xp5_ASAP7_75t_L g2299 ( 
.A1(n_2298),
.A2(n_2023),
.B(n_2074),
.C(n_2021),
.Y(n_2299)
);


endmodule