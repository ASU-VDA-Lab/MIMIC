module fake_jpeg_9915_n_108 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_12),
.B1(n_23),
.B2(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_42),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_12),
.B1(n_17),
.B2(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_20),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_17),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_10),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_9),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_39),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.C(n_66),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_37),
.B(n_34),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_18),
.B(n_26),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_52),
.B1(n_41),
.B2(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_72),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_48),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_66),
.C(n_69),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_41),
.B1(n_30),
.B2(n_45),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_65),
.B1(n_71),
.B2(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_80),
.C(n_76),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_74),
.A3(n_73),
.B1(n_80),
.B2(n_78),
.C(n_65),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_90),
.C(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_95),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_91),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_97),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_87),
.C(n_72),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_104),
.A3(n_102),
.B1(n_5),
.B2(n_7),
.C1(n_8),
.C2(n_11),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_101),
.B1(n_89),
.B2(n_45),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.B(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_4),
.Y(n_108)
);


endmodule