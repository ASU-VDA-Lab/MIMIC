module fake_jpeg_20868_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_1),
.Y(n_9)
);

BUFx10_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_10),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_21),
.B1(n_11),
.B2(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_22),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_18),
.B2(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_10),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_31),
.B(n_27),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_34),
.Y(n_39)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_14),
.B1(n_16),
.B2(n_10),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_38),
.B1(n_24),
.B2(n_27),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_44),
.B1(n_32),
.B2(n_10),
.Y(n_60)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_27),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_48),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_44),
.B(n_41),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_60),
.B1(n_54),
.B2(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_60),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_58),
.B1(n_59),
.B2(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

AOI31xp67_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_62),
.A3(n_64),
.B(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_4),
.B(n_7),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_7),
.B1(n_8),
.B2(n_3),
.Y(n_74)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_17),
.C1(n_73),
.C2(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_74),
.B(n_17),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_17),
.C(n_2),
.Y(n_78)
);


endmodule