module fake_jpeg_21500_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_30),
.B1(n_17),
.B2(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_44),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_54),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_34),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_95),
.B1(n_39),
.B2(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_65),
.B(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_40),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_71),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_72),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_77),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_53),
.B(n_35),
.Y(n_110)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_86),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_34),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_38),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_20),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_40),
.B1(n_44),
.B2(n_39),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_53),
.B1(n_52),
.B2(n_40),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_114),
.B1(n_109),
.B2(n_98),
.Y(n_135)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_67),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_40),
.B1(n_51),
.B2(n_35),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_78),
.B1(n_47),
.B2(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_111),
.B(n_22),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_0),
.B(n_1),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_84),
.B1(n_92),
.B2(n_82),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_69),
.B1(n_95),
.B2(n_77),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_29),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_99),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_22),
.Y(n_122)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_135),
.B1(n_139),
.B2(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_141),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_79),
.C(n_87),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_145),
.C(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_27),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_30),
.B1(n_80),
.B2(n_73),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_115),
.B(n_72),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_106),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_146),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_114),
.C(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_24),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_73),
.C(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_152),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_30),
.B1(n_47),
.B2(n_18),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_112),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_16),
.Y(n_170)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_23),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_25),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_142),
.A2(n_108),
.B1(n_113),
.B2(n_123),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_172),
.B1(n_174),
.B2(n_184),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_163),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_162),
.A2(n_182),
.B(n_0),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_29),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_30),
.B1(n_108),
.B2(n_123),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_19),
.B(n_1),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_180),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_18),
.A3(n_22),
.B1(n_32),
.B2(n_31),
.C1(n_19),
.C2(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_187),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_131),
.A2(n_136),
.B1(n_125),
.B2(n_145),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_124),
.C(n_74),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_176),
.C(n_165),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_96),
.B1(n_78),
.B2(n_18),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_93),
.C(n_74),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_96),
.B1(n_117),
.B2(n_101),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_178),
.B1(n_34),
.B2(n_29),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_32),
.B1(n_17),
.B2(n_24),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_17),
.B1(n_32),
.B2(n_28),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_29),
.B1(n_19),
.B2(n_31),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_31),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_137),
.A2(n_20),
.B(n_23),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_128),
.A2(n_152),
.B1(n_24),
.B2(n_25),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_128),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_193),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_190),
.B(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_154),
.C(n_56),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_200),
.C(n_208),
.Y(n_222)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_26),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_70),
.C(n_34),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_156),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_9),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_34),
.C(n_29),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_210),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_160),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_9),
.B1(n_13),
.B2(n_11),
.Y(n_211)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_162),
.Y(n_235)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_11),
.B1(n_10),
.B2(n_7),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_169),
.A2(n_11),
.B1(n_10),
.B2(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_180),
.C(n_155),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_238),
.C(n_239),
.Y(n_249)
);

FAx1_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_177),
.CI(n_169),
.CON(n_228),
.SN(n_228)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_230),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_170),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_235),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_185),
.B(n_159),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_159),
.C(n_168),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_166),
.C(n_160),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_157),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_214),
.B(n_215),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_195),
.B1(n_208),
.B2(n_217),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_234),
.B1(n_228),
.B2(n_233),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_200),
.C(n_203),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_256),
.C(n_258),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_205),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_166),
.C(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_205),
.C(n_202),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_188),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_262),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_216),
.B1(n_211),
.B2(n_184),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_221),
.B1(n_238),
.B2(n_222),
.Y(n_276)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_274),
.B1(n_248),
.B2(n_255),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_223),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_278),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_225),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_233),
.B1(n_228),
.B2(n_236),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_240),
.C(n_222),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_278),
.C(n_279),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_198),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_229),
.C(n_235),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_221),
.C(n_182),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_167),
.C(n_7),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_258),
.C(n_261),
.Y(n_284)
);

NAND2x1_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_245),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_248),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_287),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_254),
.B1(n_255),
.B2(n_247),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_247),
.C(n_5),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_2),
.C(n_3),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_5),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_0),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_0),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_4),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_296),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_302),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_285),
.B1(n_280),
.B2(n_283),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_304),
.B1(n_294),
.B2(n_292),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_264),
.B(n_2),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_282),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_291),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_307),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_313),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_281),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_289),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_4),
.C(n_2),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_3),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_310),
.A2(n_299),
.B(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_320),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_312),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_321),
.B(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_317),
.B(n_299),
.C(n_314),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_309),
.B(n_320),
.C(n_311),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_4),
.B(n_321),
.Y(n_328)
);


endmodule