module real_jpeg_8261_n_4 (n_3, n_1, n_0, n_2, n_4);

input n_3;
input n_1;
input n_0;
input n_2;

output n_4;

wire n_5;
wire n_8;
wire n_11;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_SL g5 ( 
.A1(n_1),
.A2(n_6),
.B(n_8),
.Y(n_5)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_3),
.B(n_7),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_7),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g4 ( 
.A1(n_5),
.A2(n_9),
.B(n_11),
.Y(n_4)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_5),
.B(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);


endmodule