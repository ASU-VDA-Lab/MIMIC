module fake_jpeg_26750_n_91 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_39),
.B1(n_33),
.B2(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_43),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_51),
.B(n_52),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_53),
.B1(n_5),
.B2(n_6),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_2),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_3),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_32),
.Y(n_56)
);

NAND2x1_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_5),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_67),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_18),
.C(n_30),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_6),
.A3(n_7),
.B1(n_11),
.B2(n_13),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_16),
.B1(n_27),
.B2(n_9),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_7),
.C(n_14),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_78),
.B1(n_66),
.B2(n_24),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_15),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_67),
.B(n_64),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_82),
.C(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_62),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_76),
.B1(n_73),
.B2(n_74),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_76),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_74),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_63),
.C(n_26),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_22),
.Y(n_91)
);


endmodule