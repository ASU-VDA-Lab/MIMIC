module fake_netlist_6_3962_n_1100 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1100);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1100;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g208 ( 
.A(n_68),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_88),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_5),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_108),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_22),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_38),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_26),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_139),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_35),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_41),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_15),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_16),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_47),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_160),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_143),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_119),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_166),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_37),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_19),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_159),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_16),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_150),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_82),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_52),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_7),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_123),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_29),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_185),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_76),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_71),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_204),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_75),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_205),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_54),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_39),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_25),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_72),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_200),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_207),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_146),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_183),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_14),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_170),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_77),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_106),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_178),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_121),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_98),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_66),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_46),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_105),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_114),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_214),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_225),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_223),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_227),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_225),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_244),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_263),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_245),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_210),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_237),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_217),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_218),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_231),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_219),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_213),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_221),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_213),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_226),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_234),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_250),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_229),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_230),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_243),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

OR2x6_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_252),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_253),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_256),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_209),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_251),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_255),
.B(n_243),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_319),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

OAI21x1_ASAP7_75t_L g346 ( 
.A1(n_312),
.A2(n_271),
.B(n_255),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_303),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

AND2x6_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_222),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_282),
.B(n_275),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_273),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_290),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_298),
.A2(n_272),
.B1(n_270),
.B2(n_269),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_317),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_294),
.B(n_222),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_222),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_292),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_304),
.B(n_233),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_293),
.A2(n_236),
.B(n_235),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g374 ( 
.A(n_287),
.B(n_222),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_283),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_319),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_302),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_280),
.A2(n_248),
.B1(n_240),
.B2(n_261),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_371),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_279),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_344),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_344),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_349),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_R g388 ( 
.A(n_376),
.B(n_313),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_376),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_335),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_286),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_339),
.B(n_313),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_335),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_378),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_342),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_R g401 ( 
.A(n_375),
.B(n_321),
.Y(n_401)
);

BUFx10_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_378),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_378),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_342),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_352),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_352),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_359),
.B(n_321),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_339),
.B(n_284),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_350),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_R g413 ( 
.A(n_377),
.B(n_285),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_355),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_332),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_379),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_334),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_374),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_341),
.B(n_280),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_372),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_349),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_374),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_374),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_330),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_374),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_374),
.B(n_285),
.Y(n_432)
);

AOI21x1_ASAP7_75t_L g433 ( 
.A1(n_343),
.A2(n_340),
.B(n_338),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_R g435 ( 
.A(n_374),
.B(n_286),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_R g436 ( 
.A(n_349),
.B(n_298),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_357),
.B(n_242),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_R g438 ( 
.A(n_373),
.B(n_0),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_333),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_364),
.B(n_268),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_333),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_333),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_333),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_357),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_349),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_351),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_338),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_361),
.Y(n_451)
);

NOR2x1p5_ASAP7_75t_L g452 ( 
.A(n_398),
.B(n_364),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_447),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_412),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_402),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_373),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_265),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_365),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_373),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_434),
.B(n_363),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_404),
.Y(n_472)
);

AND2x2_ASAP7_75t_SL g473 ( 
.A(n_446),
.B(n_265),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_443),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_430),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_394),
.B(n_265),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_365),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_411),
.B(n_348),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_364),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_397),
.B(n_363),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_414),
.B(n_366),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_400),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_436),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_381),
.B(n_366),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_417),
.B(n_366),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_407),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_436),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_450),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_413),
.B(n_348),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_422),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_426),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_444),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_410),
.A2(n_343),
.B1(n_365),
.B2(n_340),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_416),
.B(n_361),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_421),
.B(n_361),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_363),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_439),
.B(n_361),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_415),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_425),
.B(n_265),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_441),
.B(n_369),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_387),
.B(n_363),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_399),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_429),
.B(n_368),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_395),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_405),
.B(n_353),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_440),
.Y(n_518)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_393),
.B(n_368),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_442),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_406),
.B(n_369),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_413),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_388),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_432),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_408),
.B(n_369),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_409),
.B(n_368),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_384),
.B(n_353),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_345),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_445),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_386),
.B(n_354),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_391),
.B(n_354),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

AO22x2_ASAP7_75t_L g536 ( 
.A1(n_532),
.A2(n_438),
.B1(n_388),
.B2(n_2),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_454),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_475),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_497),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_511),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_490),
.B(n_328),
.Y(n_543)
);

NAND3x1_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_329),
.C(n_438),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_490),
.B(n_369),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_463),
.B(n_246),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_463),
.B(n_495),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_490),
.B(n_327),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_465),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_488),
.B(n_345),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_456),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_459),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_489),
.B(n_249),
.C(n_247),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_510),
.B(n_327),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_484),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_472),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_468),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_470),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_486),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_491),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_497),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_461),
.A2(n_260),
.B1(n_254),
.B2(n_213),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_531),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_516),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_533),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_471),
.B(n_480),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_496),
.B(n_500),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_497),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_524),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_478),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_478),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_531),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_485),
.B(n_343),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_520),
.B(n_3),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_524),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_525),
.B(n_326),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_469),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_506),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_453),
.B(n_346),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_533),
.B(n_346),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_501),
.B(n_326),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_512),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_453),
.B(n_326),
.Y(n_591)
);

AO22x2_ASAP7_75t_L g592 ( 
.A1(n_523),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_502),
.B(n_522),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_483),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_482),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_466),
.A2(n_527),
.B1(n_452),
.B2(n_464),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_493),
.B(n_6),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_528),
.B(n_326),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_498),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_474),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_535),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_572),
.A2(n_530),
.B(n_517),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_593),
.B(n_487),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_596),
.A2(n_526),
.B(n_504),
.C(n_508),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_575),
.B(n_519),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_571),
.B(n_518),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_589),
.B(n_467),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_552),
.B(n_467),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_540),
.B(n_515),
.Y(n_610)
);

O2A1O1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_581),
.A2(n_479),
.B(n_481),
.C(n_534),
.Y(n_611)
);

AO21x1_ASAP7_75t_L g612 ( 
.A1(n_567),
.A2(n_503),
.B(n_499),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_579),
.A2(n_509),
.B(n_473),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_540),
.Y(n_614)
);

INVx11_ASAP7_75t_L g615 ( 
.A(n_560),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_570),
.B(n_573),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_588),
.A2(n_474),
.B(n_464),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_553),
.A2(n_457),
.B(n_474),
.C(n_521),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_537),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_556),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_598),
.A2(n_514),
.B(n_505),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_551),
.A2(n_514),
.B(n_505),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_600),
.A2(n_479),
.B(n_516),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_541),
.A2(n_521),
.B1(n_529),
.B2(n_462),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_587),
.A2(n_529),
.B(n_462),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_550),
.B(n_521),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_597),
.B(n_483),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_544),
.A2(n_462),
.B(n_476),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_576),
.B(n_326),
.C(n_513),
.Y(n_630)
);

INVx11_ASAP7_75t_L g631 ( 
.A(n_583),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_557),
.B(n_462),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_537),
.A2(n_476),
.B(n_356),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_540),
.B(n_565),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_561),
.B(n_476),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_536),
.A2(n_476),
.B1(n_213),
.B2(n_507),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_542),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_538),
.A2(n_507),
.B(n_356),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_562),
.B(n_507),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_569),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_563),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_580),
.A2(n_584),
.B(n_547),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_586),
.A2(n_356),
.B(n_30),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_565),
.B(n_513),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_582),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_538),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_539),
.A2(n_356),
.B(n_31),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_566),
.B(n_356),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_539),
.A2(n_559),
.B(n_558),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_565),
.B(n_28),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_564),
.A2(n_33),
.B(n_32),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_590),
.A2(n_595),
.B(n_585),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_577),
.B(n_8),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_574),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_599),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_599),
.B(n_9),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_555),
.A2(n_36),
.B(n_34),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_583),
.A2(n_44),
.B(n_40),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_591),
.A2(n_546),
.B(n_549),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_549),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_620),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_641),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_607),
.A2(n_543),
.B(n_545),
.C(n_594),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_652),
.A2(n_583),
.B(n_543),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_SL g665 ( 
.A1(n_604),
.A2(n_583),
.B(n_578),
.C(n_568),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_622),
.A2(n_554),
.B(n_574),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_608),
.B(n_574),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_621),
.A2(n_554),
.B(n_568),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_614),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_616),
.B(n_578),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_603),
.A2(n_592),
.B(n_48),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_602),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_605),
.A2(n_592),
.B(n_11),
.C(n_12),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_606),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_SL g675 ( 
.A1(n_628),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_640),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_614),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_646),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_626),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_601),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_637),
.B(n_18),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_609),
.B(n_19),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_619),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_627),
.B(n_20),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_SL g685 ( 
.A(n_624),
.B(n_20),
.C(n_21),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_656),
.Y(n_686)
);

O2A1O1Ixp5_ASAP7_75t_SL g687 ( 
.A1(n_658),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_631),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_611),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_649),
.Y(n_690)
);

AND2x6_ASAP7_75t_SL g691 ( 
.A(n_644),
.B(n_24),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_SL g692 ( 
.A1(n_618),
.A2(n_632),
.B(n_629),
.C(n_635),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_26),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_649),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_613),
.A2(n_27),
.B1(n_45),
.B2(n_49),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_654),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_645),
.B(n_27),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_654),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_653),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_623),
.B(n_50),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_614),
.Y(n_701)
);

AOI21x1_ASAP7_75t_L g702 ( 
.A1(n_612),
.A2(n_51),
.B(n_53),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_650),
.B(n_55),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_634),
.B(n_56),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_617),
.B(n_57),
.Y(n_705)
);

OAI21x1_ASAP7_75t_L g706 ( 
.A1(n_652),
.A2(n_58),
.B(n_59),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_630),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_655),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_639),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_615),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_610),
.A2(n_67),
.B(n_69),
.C(n_70),
.Y(n_711)
);

CKINVDCx8_ASAP7_75t_R g712 ( 
.A(n_636),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_648),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_625),
.A2(n_74),
.B(n_78),
.C(n_79),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_659),
.B(n_80),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_659),
.A2(n_81),
.B(n_83),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_642),
.B(n_84),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_651),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_710),
.B(n_651),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_679),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_677),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_669),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_683),
.Y(n_723)
);

BUFx2_ASAP7_75t_R g724 ( 
.A(n_712),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_672),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_710),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_675),
.A2(n_647),
.B1(n_657),
.B2(n_643),
.Y(n_727)
);

BUFx4f_ASAP7_75t_SL g728 ( 
.A(n_676),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_677),
.Y(n_729)
);

CKINVDCx16_ASAP7_75t_R g730 ( 
.A(n_670),
.Y(n_730)
);

BUFx5_ASAP7_75t_L g731 ( 
.A(n_690),
.Y(n_731)
);

NAND2x1p5_ASAP7_75t_L g732 ( 
.A(n_688),
.B(n_657),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_701),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_688),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_667),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_669),
.Y(n_736)
);

CKINVDCx11_ASAP7_75t_R g737 ( 
.A(n_691),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_669),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_691),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_703),
.B(n_643),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_693),
.B(n_638),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_661),
.Y(n_742)
);

INVx3_ASAP7_75t_SL g743 ( 
.A(n_703),
.Y(n_743)
);

BUFx12f_ASAP7_75t_L g744 ( 
.A(n_703),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_696),
.Y(n_746)
);

BUFx4_ASAP7_75t_SL g747 ( 
.A(n_662),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_698),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_709),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_709),
.B(n_633),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_709),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_717),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_694),
.Y(n_753)
);

BUFx4_ASAP7_75t_SL g754 ( 
.A(n_699),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_681),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_718),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_697),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_717),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_686),
.B(n_633),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_713),
.Y(n_760)
);

INVx6_ASAP7_75t_SL g761 ( 
.A(n_663),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_692),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_702),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_706),
.Y(n_764)
);

NOR2x1_ASAP7_75t_SL g765 ( 
.A(n_715),
.B(n_700),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_682),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_664),
.B(n_85),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_695),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_768)
);

INVx5_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_704),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_673),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_684),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_705),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_671),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_675),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_708),
.A2(n_674),
.B1(n_680),
.B2(n_668),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_674),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_680),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_665),
.B(n_96),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_689),
.B(n_97),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_666),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_716),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_685),
.B(n_206),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_714),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_707),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_687),
.B(n_99),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_730),
.B(n_100),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_SL g788 ( 
.A1(n_783),
.A2(n_101),
.B(n_102),
.C(n_103),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_756),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_756),
.Y(n_790)
);

AOI221xp5_ASAP7_75t_SL g791 ( 
.A1(n_776),
.A2(n_104),
.B1(n_107),
.B2(n_109),
.C(n_110),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_754),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_764),
.A2(n_111),
.B(n_112),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_749),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_722),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_723),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_764),
.A2(n_113),
.B(n_115),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_727),
.A2(n_116),
.B(n_117),
.C(n_118),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_753),
.Y(n_799)
);

AOI221xp5_ASAP7_75t_L g800 ( 
.A1(n_771),
.A2(n_780),
.B1(n_778),
.B2(n_777),
.C(n_775),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_725),
.Y(n_801)
);

NOR2xp67_ASAP7_75t_L g802 ( 
.A(n_726),
.B(n_120),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_745),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_782),
.A2(n_122),
.B(n_124),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_727),
.A2(n_126),
.B(n_127),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_750),
.A2(n_128),
.B(n_129),
.Y(n_807)
);

NOR2x1_ASAP7_75t_L g808 ( 
.A(n_770),
.B(n_766),
.Y(n_808)
);

OAI221xp5_ASAP7_75t_L g809 ( 
.A1(n_757),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.C(n_134),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_772),
.B(n_135),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_749),
.Y(n_811)
);

BUFx2_ASAP7_75t_SL g812 ( 
.A(n_734),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_724),
.B(n_136),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_751),
.B(n_137),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_765),
.A2(n_140),
.B(n_141),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_735),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_735),
.B(n_142),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_728),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_730),
.B(n_144),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_763),
.A2(n_774),
.B(n_785),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_731),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_774),
.A2(n_145),
.B(n_148),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_767),
.A2(n_732),
.B(n_763),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_771),
.B(n_149),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_747),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_748),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_SL g827 ( 
.A1(n_739),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_781),
.A2(n_155),
.B(n_156),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_746),
.Y(n_829)
);

AO21x2_ASAP7_75t_L g830 ( 
.A1(n_785),
.A2(n_157),
.B(n_158),
.Y(n_830)
);

CKINVDCx12_ASAP7_75t_R g831 ( 
.A(n_740),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_755),
.A2(n_162),
.B(n_163),
.C(n_164),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_773),
.B(n_165),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_779),
.A2(n_743),
.B(n_740),
.C(n_786),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_731),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_731),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_733),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_719),
.A2(n_168),
.B(n_169),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_752),
.B(n_171),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_768),
.A2(n_172),
.B(n_173),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_772),
.A2(n_761),
.B1(n_769),
.B2(n_744),
.Y(n_841)
);

CKINVDCx11_ASAP7_75t_R g842 ( 
.A(n_818),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_789),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_790),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_799),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_800),
.A2(n_737),
.B1(n_761),
.B2(n_784),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_816),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_820),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_820),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_821),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_808),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_835),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_836),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_796),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_801),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_804),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_803),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_823),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_831),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_830),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_804),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_815),
.A2(n_759),
.B(n_741),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_830),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_829),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_805),
.Y(n_865)
);

NAND2x1_ASAP7_75t_L g866 ( 
.A(n_815),
.B(n_758),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_794),
.Y(n_867)
);

AO21x2_ASAP7_75t_L g868 ( 
.A1(n_806),
.A2(n_769),
.B(n_784),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_806),
.A2(n_784),
.B1(n_769),
.B2(n_752),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_824),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_804),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_839),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_837),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_839),
.Y(n_874)
);

AO21x2_ASAP7_75t_L g875 ( 
.A1(n_834),
.A2(n_781),
.B(n_762),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_822),
.A2(n_752),
.B(n_758),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_837),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_794),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_811),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_809),
.A2(n_762),
.B1(n_772),
.B2(n_760),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_833),
.Y(n_882)
);

BUFx4f_ASAP7_75t_SL g883 ( 
.A(n_795),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_795),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_824),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_826),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_787),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_838),
.B(n_762),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_846),
.A2(n_800),
.B(n_798),
.Y(n_889)
);

CKINVDCx11_ASAP7_75t_R g890 ( 
.A(n_842),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_848),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_R g892 ( 
.A(n_870),
.B(n_792),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_869),
.A2(n_828),
.B(n_832),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_847),
.B(n_841),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_873),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_843),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_876),
.B(n_812),
.Y(n_897)
);

AO31x2_ASAP7_75t_L g898 ( 
.A1(n_863),
.A2(n_828),
.A3(n_833),
.B(n_817),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_868),
.A2(n_809),
.B1(n_822),
.B2(n_827),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_873),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_873),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_843),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_877),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_881),
.A2(n_832),
.B(n_791),
.C(n_813),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_844),
.Y(n_905)
);

CKINVDCx16_ASAP7_75t_R g906 ( 
.A(n_871),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_871),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_868),
.A2(n_742),
.B1(n_819),
.B2(n_810),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_844),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_856),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_R g911 ( 
.A(n_883),
.B(n_825),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_877),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_877),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_R g914 ( 
.A(n_870),
.B(n_817),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_845),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_871),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_847),
.B(n_791),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_866),
.B(n_797),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_856),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_866),
.B(n_793),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_872),
.B(n_729),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_845),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_856),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_885),
.B(n_814),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_868),
.A2(n_840),
.B1(n_814),
.B2(n_802),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_914),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_891),
.B(n_895),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_914),
.Y(n_928)
);

AND2x4_ASAP7_75t_SL g929 ( 
.A(n_897),
.B(n_872),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_896),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_891),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_890),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_902),
.Y(n_933)
);

AO31x2_ASAP7_75t_L g934 ( 
.A1(n_905),
.A2(n_848),
.A3(n_849),
.B(n_860),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_903),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_900),
.B(n_850),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_909),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_915),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_922),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_901),
.B(n_885),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_912),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_889),
.A2(n_859),
.B1(n_887),
.B2(n_875),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_906),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_897),
.B(n_907),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_SL g945 ( 
.A1(n_893),
.A2(n_875),
.B1(n_872),
.B2(n_874),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_894),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_910),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_923),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_945),
.A2(n_899),
.B1(n_897),
.B2(n_859),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_926),
.B(n_921),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_946),
.B(n_928),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_934),
.Y(n_952)
);

OA21x2_ASAP7_75t_L g953 ( 
.A1(n_931),
.A2(n_849),
.B(n_917),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_942),
.A2(n_899),
.B1(n_908),
.B2(n_887),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_944),
.B(n_916),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_940),
.B(n_886),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_934),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_933),
.Y(n_958)
);

NAND2x1p5_ASAP7_75t_SL g959 ( 
.A(n_944),
.B(n_882),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_929),
.A2(n_904),
.B(n_875),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_927),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_934),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_934),
.Y(n_963)
);

AOI211xp5_ASAP7_75t_L g964 ( 
.A1(n_932),
.A2(n_788),
.B(n_924),
.C(n_851),
.Y(n_964)
);

AO21x2_ASAP7_75t_L g965 ( 
.A1(n_931),
.A2(n_860),
.B(n_863),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_961),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_949),
.A2(n_892),
.B1(n_929),
.B2(n_908),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_958),
.Y(n_968)
);

OAI33xp33_ASAP7_75t_L g969 ( 
.A1(n_950),
.A2(n_930),
.A3(n_937),
.B1(n_927),
.B2(n_852),
.B3(n_853),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_955),
.B(n_943),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_955),
.B(n_932),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_956),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_950),
.B(n_943),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_952),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_SL g975 ( 
.A1(n_960),
.A2(n_892),
.B1(n_921),
.B2(n_872),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_951),
.B(n_935),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_953),
.B(n_933),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_954),
.B(n_936),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_971),
.B(n_936),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_975),
.B(n_964),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_966),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_971),
.B(n_941),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_974),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_970),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_973),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_972),
.B(n_953),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_985),
.B(n_978),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_981),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_980),
.A2(n_967),
.B(n_975),
.C(n_976),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_982),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_984),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_991),
.B(n_979),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_988),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_987),
.B(n_983),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_968),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_989),
.B(n_986),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_990),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_990),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_991),
.B(n_986),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_991),
.B(n_959),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_988),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_995),
.B(n_959),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_996),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_994),
.Y(n_1005)
);

CKINVDCx16_ASAP7_75t_R g1006 ( 
.A(n_999),
.Y(n_1006)
);

AND2x2_ASAP7_75t_SL g1007 ( 
.A(n_998),
.B(n_911),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1000),
.B(n_977),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_998),
.B(n_911),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_993),
.B(n_1002),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_SL g1011 ( 
.A1(n_1007),
.A2(n_1001),
.B(n_997),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_R g1012 ( 
.A(n_1006),
.B(n_856),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_1009),
.A2(n_977),
.B(n_952),
.C(n_963),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1004),
.B(n_1005),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_1010),
.B(n_969),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1003),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1008),
.B(n_953),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1014),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_1011),
.B(n_969),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1016),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_1012),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1017),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1020),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1018),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1021),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1019),
.B(n_1015),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1022),
.B(n_1013),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1020),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1025),
.B(n_938),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_1026),
.A2(n_1028),
.B1(n_1023),
.B2(n_1027),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_L g1031 ( 
.A(n_1024),
.B(n_874),
.C(n_807),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1025),
.B(n_938),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1025),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_856),
.C(n_861),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_SL g1035 ( 
.A1(n_1033),
.A2(n_884),
.B(n_963),
.C(n_962),
.Y(n_1035)
);

AOI21xp33_ASAP7_75t_SL g1036 ( 
.A1(n_1030),
.A2(n_174),
.B(n_175),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1034),
.A2(n_861),
.B1(n_947),
.B2(n_957),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1029),
.Y(n_1038)
);

AOI211xp5_ASAP7_75t_L g1039 ( 
.A1(n_1032),
.A2(n_861),
.B(n_947),
.C(n_872),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_L g1040 ( 
.A(n_1036),
.B(n_1038),
.C(n_1039),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_1035),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_1037),
.A2(n_1031),
.B1(n_861),
.B2(n_947),
.Y(n_1042)
);

AOI221xp5_ASAP7_75t_L g1043 ( 
.A1(n_1036),
.A2(n_962),
.B1(n_957),
.B2(n_947),
.C(n_861),
.Y(n_1043)
);

AO22x2_ASAP7_75t_L g1044 ( 
.A1(n_1038),
.A2(n_884),
.B1(n_948),
.B2(n_874),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_L g1045 ( 
.A(n_1038),
.B(n_874),
.C(n_729),
.Y(n_1045)
);

AOI222xp33_ASAP7_75t_L g1046 ( 
.A1(n_1038),
.A2(n_947),
.B1(n_925),
.B2(n_864),
.C1(n_939),
.C2(n_910),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_1036),
.A2(n_736),
.B(n_939),
.C(n_923),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_1041),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_L g1050 ( 
.A(n_1043),
.B(n_738),
.C(n_722),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1045),
.Y(n_1051)
);

OAI321xp33_ASAP7_75t_L g1052 ( 
.A1(n_1042),
.A2(n_1046),
.A3(n_925),
.B1(n_722),
.B2(n_738),
.C(n_910),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1040),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1040),
.B(n_965),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_1040),
.B(n_919),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1041),
.B(n_965),
.Y(n_1056)
);

OAI311xp33_ASAP7_75t_L g1057 ( 
.A1(n_1054),
.A2(n_721),
.A3(n_858),
.B1(n_854),
.C1(n_855),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1055),
.Y(n_1058)
);

NAND4xp75_ASAP7_75t_L g1059 ( 
.A(n_1048),
.B(n_176),
.C(n_177),
.D(n_179),
.Y(n_1059)
);

XNOR2xp5_ASAP7_75t_L g1060 ( 
.A(n_1053),
.B(n_1049),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_L g1061 ( 
.A(n_1051),
.B(n_864),
.C(n_862),
.Y(n_1061)
);

OAI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1050),
.A2(n_918),
.B1(n_920),
.B2(n_738),
.C(n_882),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1052),
.B(n_180),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1056),
.A2(n_965),
.B1(n_888),
.B2(n_858),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_1053),
.B(n_898),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1055),
.B(n_898),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1055),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1055),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_SL g1069 ( 
.A1(n_1053),
.A2(n_920),
.B1(n_918),
.B2(n_888),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_L g1070 ( 
.A(n_1059),
.B(n_181),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_1060),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_1058),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1067),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1068),
.B(n_1063),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_1065),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_1066),
.Y(n_1076)
);

OAI221xp5_ASAP7_75t_SL g1077 ( 
.A1(n_1062),
.A2(n_920),
.B1(n_918),
.B2(n_880),
.C(n_867),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1069),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1073),
.A2(n_1057),
.B(n_1064),
.Y(n_1079)
);

AO22x2_ASAP7_75t_L g1080 ( 
.A1(n_1071),
.A2(n_1061),
.B1(n_880),
.B2(n_878),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1072),
.A2(n_888),
.B1(n_858),
.B2(n_879),
.Y(n_1081)
);

XNOR2xp5_ASAP7_75t_L g1082 ( 
.A(n_1070),
.B(n_182),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1078),
.A2(n_1077),
.B1(n_1074),
.B2(n_1075),
.Y(n_1083)
);

XNOR2xp5_ASAP7_75t_L g1084 ( 
.A(n_1076),
.B(n_186),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1084),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1082),
.B(n_188),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1083),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_1086),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1088),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1089),
.A2(n_1087),
.B(n_1079),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1090),
.A2(n_1085),
.B1(n_1080),
.B2(n_1081),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1090),
.Y(n_1092)
);

OAI222xp33_ASAP7_75t_L g1093 ( 
.A1(n_1092),
.A2(n_862),
.B1(n_858),
.B2(n_865),
.C1(n_878),
.C2(n_867),
.Y(n_1093)
);

AOI222xp33_ASAP7_75t_L g1094 ( 
.A1(n_1091),
.A2(n_888),
.B1(n_853),
.B2(n_852),
.C1(n_865),
.C2(n_195),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1094),
.A2(n_189),
.B1(n_191),
.B2(n_193),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1093),
.A2(n_854),
.B1(n_855),
.B2(n_857),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_1095),
.A2(n_1096),
.B(n_196),
.Y(n_1097)
);

AO21x2_ASAP7_75t_L g1098 ( 
.A1(n_1095),
.A2(n_194),
.B(n_197),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_198),
.B(n_199),
.Y(n_1099)
);

AOI211xp5_ASAP7_75t_L g1100 ( 
.A1(n_1099),
.A2(n_1098),
.B(n_201),
.C(n_203),
.Y(n_1100)
);


endmodule