module fake_jpeg_3684_n_230 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_33),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_90),
.Y(n_95)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_71),
.Y(n_99)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_80),
.B1(n_78),
.B2(n_56),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_94),
.B1(n_98),
.B2(n_100),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_89),
.B1(n_78),
.B2(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_79),
.B1(n_64),
.B2(n_62),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_81),
.B(n_59),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_79),
.B1(n_62),
.B2(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_74),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_67),
.B1(n_72),
.B2(n_68),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_55),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_101),
.Y(n_110)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_55),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_57),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_86),
.B1(n_75),
.B2(n_63),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_68),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_73),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_104),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_76),
.B(n_87),
.C(n_60),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_140),
.B(n_118),
.C(n_61),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_130),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_98),
.B(n_68),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_138),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_1),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_75),
.B(n_63),
.C(n_61),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_49),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_155),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_156),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_77),
.B(n_4),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_77),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_169),
.B1(n_173),
.B2(n_14),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_2),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_161),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_6),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_7),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_8),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_126),
.B(n_8),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_170),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_25),
.B1(n_42),
.B2(n_41),
.Y(n_168)
);

AOI22x1_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_23),
.C(n_40),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_43),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_15),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_173)
);

AO21x1_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_134),
.B(n_147),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_147),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_186),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_181),
.B1(n_188),
.B2(n_160),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_14),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_187),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_172),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_193),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_16),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_39),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_175),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_199),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_168),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_170),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_204),
.B1(n_178),
.B2(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_169),
.B1(n_148),
.B2(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_206),
.B(n_207),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_174),
.B1(n_190),
.B2(n_176),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_177),
.B1(n_193),
.B2(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_212),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_183),
.C(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_194),
.C(n_196),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_30),
.Y(n_216)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_19),
.B(n_20),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_216),
.C(n_218),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_211),
.C(n_209),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_21),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_213),
.C(n_26),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_21),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_224),
.B1(n_220),
.B2(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_29),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_31),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_34),
.B(n_37),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_38),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_205),
.Y(n_230)
);


endmodule