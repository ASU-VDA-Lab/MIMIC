module real_jpeg_16785_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_23;
wire n_14;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_1),
.A2(n_15),
.B1(n_16),
.B2(n_28),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_2),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_19),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_7),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_8),
.B(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_39),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_34),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_29),
.Y(n_13)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_25),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_24),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_43),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_42),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_26),
.C(n_27),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);


endmodule