module fake_jpeg_9448_n_194 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_194);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_35),
.B1(n_15),
.B2(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_22),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_45),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_28),
.C(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_24),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_46),
.B1(n_51),
.B2(n_32),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_36),
.B1(n_29),
.B2(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_30),
.B1(n_49),
.B2(n_47),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_27),
.B(n_22),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_42),
.C(n_41),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_68),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_33),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_34),
.B1(n_30),
.B2(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_34),
.B1(n_30),
.B2(n_31),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_47),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_34),
.B1(n_30),
.B2(n_26),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_52),
.B1(n_57),
.B2(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_76),
.B(n_79),
.Y(n_109)
);

OAI31xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_45),
.A3(n_42),
.B(n_39),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_85),
.B(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_93),
.B1(n_94),
.B2(n_54),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_33),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_16),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_49),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_0),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_1),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_47),
.B1(n_33),
.B2(n_25),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_16),
.B1(n_50),
.B2(n_22),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_115),
.B1(n_94),
.B2(n_80),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_54),
.B(n_68),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_111),
.B(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_102),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_67),
.B1(n_56),
.B2(n_61),
.Y(n_101)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_112),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_1),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_105),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_2),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_95),
.C(n_81),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_70),
.B1(n_61),
.B2(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_131),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_77),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.C(n_129),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_133),
.B1(n_104),
.B2(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_99),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_89),
.B(n_93),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_97),
.B1(n_72),
.B2(n_110),
.C(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_84),
.B1(n_81),
.B2(n_82),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_108),
.C(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_143),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_109),
.C(n_83),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_76),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_147),
.C(n_125),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_111),
.B(n_107),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_146),
.B(n_148),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_91),
.C(n_106),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_101),
.B1(n_91),
.B2(n_78),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_101),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_116),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_121),
.B1(n_123),
.B2(n_117),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_118),
.B1(n_128),
.B2(n_135),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_139),
.B1(n_70),
.B2(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_162),
.B(n_7),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_167),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_139),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_159),
.C(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_135),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_163),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B(n_9),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_7),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_6),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_158),
.B(n_155),
.C(n_163),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_178),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_164),
.B(n_12),
.Y(n_181)
);

NOR4xp25_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_161),
.C(n_7),
.D(n_8),
.Y(n_176)
);

AOI31xp67_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_180),
.A3(n_2),
.B(n_3),
.Y(n_182)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_2),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_180),
.B1(n_164),
.B2(n_177),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_3),
.C(n_4),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_5),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_185),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_5),
.C(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_5),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_191),
.C(n_5),
.Y(n_194)
);


endmodule