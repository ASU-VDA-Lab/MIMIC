module real_aes_8704_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g537 ( .A1(n_0), .A2(n_187), .B(n_538), .C(n_541), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_1), .B(n_526), .Y(n_542) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_3), .A2(n_745), .B1(n_748), .B2(n_749), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_3), .Y(n_749) );
INVx1_ASAP7_75t_L g205 ( .A(n_4), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_5), .B(n_176), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_6), .A2(n_441), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_7), .A2(n_152), .B(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_8), .A2(n_37), .B1(n_132), .B2(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_9), .B(n_152), .Y(n_216) );
AND2x6_ASAP7_75t_L g150 ( .A(n_10), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_11), .A2(n_150), .B(n_444), .C(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_12), .B(n_38), .Y(n_113) );
INVx1_ASAP7_75t_L g148 ( .A(n_13), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_14), .B(n_139), .Y(n_159) );
INVx1_ASAP7_75t_L g197 ( .A(n_15), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_16), .B(n_176), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_17), .B(n_153), .Y(n_221) );
AO32x2_ASAP7_75t_L g184 ( .A1(n_18), .A2(n_149), .A3(n_152), .B1(n_185), .B2(n_189), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_19), .B(n_141), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_20), .B(n_153), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_21), .A2(n_53), .B1(n_132), .B2(n_141), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g138 ( .A1(n_22), .A2(n_82), .B1(n_139), .B2(n_141), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_23), .B(n_141), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_24), .A2(n_149), .B(n_444), .C(n_446), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_25), .A2(n_149), .B(n_444), .C(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_26), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_27), .B(n_144), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_28), .A2(n_103), .B1(n_114), .B2(n_756), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_29), .A2(n_441), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_30), .B(n_144), .Y(n_182) );
INVx2_ASAP7_75t_L g134 ( .A(n_31), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_32), .A2(n_465), .B(n_474), .C(n_476), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_33), .B(n_141), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_34), .B(n_144), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_35), .A2(n_74), .B1(n_117), .B2(n_118), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_35), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_36), .B(n_161), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_39), .B(n_440), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_40), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_41), .B(n_176), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_42), .B(n_441), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_43), .A2(n_465), .B(n_474), .C(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_44), .A2(n_122), .B1(n_426), .B2(n_427), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_44), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_44), .A2(n_80), .B1(n_426), .B2(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_45), .B(n_141), .Y(n_211) );
INVx1_ASAP7_75t_L g539 ( .A(n_46), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_47), .A2(n_90), .B1(n_132), .B2(n_135), .Y(n_131) );
INVx1_ASAP7_75t_L g512 ( .A(n_48), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_49), .B(n_141), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_50), .B(n_141), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_51), .B(n_441), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_52), .B(n_203), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_54), .A2(n_59), .B1(n_139), .B2(n_141), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_55), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_56), .B(n_141), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_57), .B(n_141), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_58), .Y(n_753) );
INVx1_ASAP7_75t_L g151 ( .A(n_60), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_61), .B(n_441), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_62), .B(n_526), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_63), .A2(n_200), .B(n_203), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_64), .B(n_141), .Y(n_206) );
INVx1_ASAP7_75t_L g147 ( .A(n_65), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_66), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_67), .B(n_176), .Y(n_478) );
AO32x2_ASAP7_75t_L g129 ( .A1(n_68), .A2(n_130), .A3(n_143), .B1(n_149), .B2(n_152), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_69), .B(n_142), .Y(n_502) );
INVx1_ASAP7_75t_L g239 ( .A(n_70), .Y(n_239) );
INVx1_ASAP7_75t_L g174 ( .A(n_71), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_72), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_73), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g118 ( .A(n_74), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_75), .A2(n_444), .B(n_461), .C(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_76), .B(n_139), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_77), .Y(n_521) );
INVx1_ASAP7_75t_L g107 ( .A(n_78), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_79), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_80), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_81), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_83), .B(n_132), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_84), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_85), .B(n_139), .Y(n_179) );
INVx2_ASAP7_75t_L g145 ( .A(n_86), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_87), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_88), .B(n_136), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_89), .B(n_139), .Y(n_212) );
OR2x2_ASAP7_75t_L g109 ( .A(n_91), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g430 ( .A(n_91), .B(n_111), .Y(n_430) );
INVx2_ASAP7_75t_L g727 ( .A(n_91), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_92), .A2(n_101), .B1(n_139), .B2(n_140), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_93), .B(n_441), .Y(n_472) );
INVx1_ASAP7_75t_L g477 ( .A(n_94), .Y(n_477) );
INVxp67_ASAP7_75t_L g524 ( .A(n_95), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_96), .B(n_139), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_97), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g462 ( .A(n_98), .Y(n_462) );
INVx1_ASAP7_75t_L g498 ( .A(n_99), .Y(n_498) );
AND2x2_ASAP7_75t_L g514 ( .A(n_100), .B(n_144), .Y(n_514) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g757 ( .A(n_104), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_108), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g755 ( .A(n_109), .Y(n_755) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_110), .B(n_727), .Y(n_739) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g726 ( .A(n_111), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AO221x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_740), .B1(n_743), .B2(n_750), .C(n_752), .Y(n_114) );
OAI222xp33_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_119), .B1(n_728), .B2(n_729), .C1(n_735), .C2(n_736), .Y(n_115) );
INVx1_ASAP7_75t_L g728 ( .A(n_116), .Y(n_728) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_428), .B1(n_431), .B2(n_724), .Y(n_120) );
INVx1_ASAP7_75t_L g731 ( .A(n_121), .Y(n_731) );
INVx2_ASAP7_75t_L g427 ( .A(n_122), .Y(n_427) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
XOR2x2_ASAP7_75t_L g745 ( .A(n_123), .B(n_746), .Y(n_745) );
AND3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_346), .C(n_394), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_274), .C(n_319), .D(n_333), .Y(n_124) );
OAI311xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_190), .A3(n_217), .B1(n_227), .C1(n_242), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_154), .Y(n_126) );
OAI21xp33_ASAP7_75t_L g227 ( .A1(n_127), .A2(n_228), .B(n_230), .Y(n_227) );
AND2x2_ASAP7_75t_L g335 ( .A(n_127), .B(n_262), .Y(n_335) );
AND2x2_ASAP7_75t_L g392 ( .A(n_127), .B(n_278), .Y(n_392) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g285 ( .A(n_128), .B(n_183), .Y(n_285) );
AND2x2_ASAP7_75t_L g342 ( .A(n_128), .B(n_290), .Y(n_342) );
INVx1_ASAP7_75t_L g383 ( .A(n_128), .Y(n_383) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_129), .Y(n_251) );
AND2x2_ASAP7_75t_L g292 ( .A(n_129), .B(n_183), .Y(n_292) );
AND2x2_ASAP7_75t_L g296 ( .A(n_129), .B(n_184), .Y(n_296) );
INVx1_ASAP7_75t_L g308 ( .A(n_129), .Y(n_308) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_136), .B1(n_138), .B2(n_142), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx3_ASAP7_75t_L g135 ( .A(n_133), .Y(n_135) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
AND2x6_ASAP7_75t_L g444 ( .A(n_133), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx1_ASAP7_75t_L g204 ( .A(n_134), .Y(n_204) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_135), .Y(n_479) );
INVx2_ASAP7_75t_L g541 ( .A(n_135), .Y(n_541) );
INVx2_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_136), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_136), .A2(n_187), .B1(n_224), .B2(n_225), .Y(n_223) );
INVx4_ASAP7_75t_L g540 ( .A(n_136), .Y(n_540) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g142 ( .A(n_137), .Y(n_142) );
INVx1_ASAP7_75t_L g161 ( .A(n_137), .Y(n_161) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
AND2x2_ASAP7_75t_L g442 ( .A(n_137), .B(n_204), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_137), .Y(n_445) );
INVx2_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_141), .Y(n_464) );
INVx5_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx1_ASAP7_75t_L g451 ( .A(n_143), .Y(n_451) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_144), .A2(n_156), .B(n_166), .Y(n_155) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_144), .A2(n_171), .B(n_182), .Y(n_170) );
INVx1_ASAP7_75t_L g454 ( .A(n_144), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_144), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_144), .A2(n_509), .B(n_510), .Y(n_508) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_L g153 ( .A(n_145), .B(n_146), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_149), .B(n_223), .C(n_226), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_149), .A2(n_235), .B(n_238), .Y(n_234) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_150), .A2(n_157), .B(n_162), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_150), .A2(n_172), .B(n_177), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_150), .A2(n_196), .B(n_201), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_150), .A2(n_210), .B(n_213), .Y(n_209) );
AND2x4_ASAP7_75t_L g441 ( .A(n_150), .B(n_442), .Y(n_441) );
INVx4_ASAP7_75t_SL g466 ( .A(n_150), .Y(n_466) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_150), .B(n_442), .Y(n_499) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_152), .A2(n_209), .B(n_216), .Y(n_208) );
INVx4_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_152), .A2(n_489), .B(n_490), .Y(n_488) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_152), .Y(n_518) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_167), .Y(n_154) );
AND2x2_ASAP7_75t_L g229 ( .A(n_155), .B(n_183), .Y(n_229) );
INVx2_ASAP7_75t_L g263 ( .A(n_155), .Y(n_263) );
AND2x2_ASAP7_75t_L g278 ( .A(n_155), .B(n_184), .Y(n_278) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_155), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_155), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g298 ( .A(n_155), .B(n_261), .Y(n_298) );
INVx1_ASAP7_75t_L g310 ( .A(n_155), .Y(n_310) );
INVx1_ASAP7_75t_L g351 ( .A(n_155), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_155), .B(n_251), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_160), .Y(n_157) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_L g238 ( .A1(n_165), .A2(n_202), .B(n_239), .C(n_240), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g167 ( .A(n_168), .B(n_183), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g228 ( .A(n_169), .B(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_169), .Y(n_256) );
AND2x2_ASAP7_75t_SL g309 ( .A(n_169), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g313 ( .A(n_169), .B(n_183), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_169), .B(n_308), .Y(n_371) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g261 ( .A(n_170), .Y(n_261) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_170), .Y(n_277) );
OR2x2_ASAP7_75t_L g350 ( .A(n_170), .B(n_351), .Y(n_350) );
O2A1O1Ixp5_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_176), .Y(n_172) );
INVx2_ASAP7_75t_L g187 ( .A(n_176), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_176), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_176), .A2(n_236), .B(n_237), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_176), .B(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_177) );
INVx1_ASAP7_75t_L g200 ( .A(n_180), .Y(n_200) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g448 ( .A(n_181), .Y(n_448) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx2_ASAP7_75t_L g257 ( .A(n_184), .Y(n_257) );
AND2x2_ASAP7_75t_L g262 ( .A(n_184), .B(n_263), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_187), .A2(n_202), .B(n_205), .C(n_206), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_187), .A2(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g194 ( .A(n_189), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_189), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_190), .B(n_245), .Y(n_408) );
INVx1_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g378 ( .A(n_191), .B(n_219), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_208), .Y(n_191) );
AND2x2_ASAP7_75t_L g254 ( .A(n_192), .B(n_245), .Y(n_254) );
INVx2_ASAP7_75t_L g266 ( .A(n_192), .Y(n_266) );
AND2x2_ASAP7_75t_L g300 ( .A(n_192), .B(n_248), .Y(n_300) );
AND2x2_ASAP7_75t_L g367 ( .A(n_192), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_193), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g247 ( .A(n_193), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g287 ( .A(n_193), .B(n_208), .Y(n_287) );
AND2x2_ASAP7_75t_L g304 ( .A(n_193), .B(n_305), .Y(n_304) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_207), .Y(n_193) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_194), .A2(n_234), .B(n_241), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .C(n_200), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_198), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_198), .A2(n_502), .B(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_200), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_202), .A2(n_447), .B(n_449), .Y(n_446) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g230 ( .A(n_208), .B(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
AND2x2_ASAP7_75t_L g253 ( .A(n_208), .B(n_233), .Y(n_253) );
AND2x2_ASAP7_75t_L g326 ( .A(n_208), .B(n_305), .Y(n_326) );
AND2x2_ASAP7_75t_L g391 ( .A(n_208), .B(n_381), .Y(n_391) );
OAI311xp33_ASAP7_75t_L g274 ( .A1(n_217), .A2(n_275), .A3(n_279), .B1(n_281), .C1(n_301), .Y(n_274) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g286 ( .A(n_218), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g345 ( .A(n_218), .B(n_253), .Y(n_345) );
AND2x2_ASAP7_75t_L g419 ( .A(n_218), .B(n_300), .Y(n_419) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_219), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g354 ( .A(n_219), .Y(n_354) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g245 ( .A(n_220), .Y(n_245) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_220), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g374 ( .A(n_220), .B(n_248), .Y(n_374) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
AO21x1_ASAP7_75t_L g270 ( .A1(n_223), .A2(n_226), .B(n_271), .Y(n_270) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_226), .A2(n_459), .B(n_468), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_226), .B(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_226), .B(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_226), .A2(n_497), .B(n_504), .Y(n_496) );
INVx3_ASAP7_75t_L g526 ( .A(n_226), .Y(n_526) );
AND2x2_ASAP7_75t_L g249 ( .A(n_229), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g302 ( .A(n_229), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g382 ( .A(n_229), .B(n_383), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_230), .A2(n_262), .B1(n_282), .B2(n_286), .C(n_288), .Y(n_281) );
INVx1_ASAP7_75t_L g406 ( .A(n_231), .Y(n_406) );
OR2x2_ASAP7_75t_L g372 ( .A(n_232), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g267 ( .A(n_233), .B(n_248), .Y(n_267) );
OR2x2_ASAP7_75t_L g269 ( .A(n_233), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g294 ( .A(n_233), .Y(n_294) );
INVx2_ASAP7_75t_L g305 ( .A(n_233), .Y(n_305) );
AND2x2_ASAP7_75t_L g332 ( .A(n_233), .B(n_270), .Y(n_332) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_233), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_249), .B1(n_252), .B2(n_255), .C(n_258), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g343 ( .A(n_245), .B(n_253), .Y(n_343) );
AND2x2_ASAP7_75t_L g393 ( .A(n_245), .B(n_247), .Y(n_393) );
INVx2_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g280 ( .A(n_247), .B(n_251), .Y(n_280) );
AND2x2_ASAP7_75t_L g359 ( .A(n_247), .B(n_332), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_248), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g318 ( .A(n_248), .Y(n_318) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_249), .A2(n_329), .B(n_331), .Y(n_328) );
OR2x2_ASAP7_75t_L g272 ( .A(n_250), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g338 ( .A(n_250), .B(n_298), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_250), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g315 ( .A(n_251), .B(n_284), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_251), .B(n_398), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_252), .B(n_278), .Y(n_388) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g311 ( .A(n_253), .B(n_266), .Y(n_311) );
INVx1_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .B1(n_268), .B2(n_272), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g290 ( .A(n_261), .Y(n_290) );
INVx1_ASAP7_75t_L g303 ( .A(n_261), .Y(n_303) );
INVx1_ASAP7_75t_L g273 ( .A(n_262), .Y(n_273) );
AND2x2_ASAP7_75t_L g344 ( .A(n_262), .B(n_290), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_262), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
OR2x2_ASAP7_75t_L g268 ( .A(n_265), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_265), .B(n_381), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_265), .B(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g415 ( .A(n_267), .B(n_367), .Y(n_415) );
INVx1_ASAP7_75t_SL g381 ( .A(n_269), .Y(n_381) );
AND2x2_ASAP7_75t_L g321 ( .A(n_270), .B(n_305), .Y(n_321) );
INVx1_ASAP7_75t_L g368 ( .A(n_270), .Y(n_368) );
OAI222xp33_ASAP7_75t_L g409 ( .A1(n_275), .A2(n_365), .B1(n_410), .B2(n_411), .C1(n_414), .C2(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
AND2x2_ASAP7_75t_L g341 ( .A(n_278), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_278), .B(n_383), .Y(n_410) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_280), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g385 ( .A(n_282), .Y(n_385) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g323 ( .A(n_285), .Y(n_323) );
AND2x2_ASAP7_75t_L g402 ( .A(n_285), .B(n_363), .Y(n_402) );
AND2x2_ASAP7_75t_L g425 ( .A(n_285), .B(n_309), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_287), .B(n_321), .Y(n_320) );
OAI32xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .A3(n_293), .B1(n_295), .B2(n_299), .Y(n_288) );
BUFx2_ASAP7_75t_L g363 ( .A(n_290), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_291), .B(n_309), .Y(n_390) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g329 ( .A(n_292), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g397 ( .A(n_292), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g386 ( .A(n_293), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g357 ( .A(n_296), .B(n_330), .Y(n_357) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OAI221xp5_ASAP7_75t_SL g319 ( .A1(n_298), .A2(n_320), .B1(n_322), .B2(n_324), .C(n_328), .Y(n_319) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g331 ( .A(n_300), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g337 ( .A(n_300), .B(n_321), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_304), .B1(n_306), .B2(n_311), .C(n_312), .Y(n_301) );
INVx1_ASAP7_75t_L g420 ( .A(n_302), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_303), .B(n_397), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_304), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_309), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g375 ( .A(n_309), .Y(n_375) );
BUFx3_ASAP7_75t_L g398 ( .A(n_310), .Y(n_398) );
INVx1_ASAP7_75t_SL g339 ( .A(n_311), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_311), .B(n_353), .Y(n_352) );
AOI21xp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_314), .B(n_316), .Y(n_312) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_313), .A2(n_414), .B1(n_418), .B2(n_420), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_321), .Y(n_360) );
INVx1_ASAP7_75t_L g424 ( .A(n_318), .Y(n_424) );
INVx2_ASAP7_75t_L g413 ( .A(n_321), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_321), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g366 ( .A(n_326), .B(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B1(n_338), .B2(n_339), .C(n_340), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_342), .A2(n_404), .B1(n_405), .B2(n_407), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_345), .A2(n_422), .B(n_425), .Y(n_421) );
NOR4xp25_ASAP7_75t_SL g346 ( .A(n_347), .B(n_355), .C(n_364), .D(n_384), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B1(n_361), .B2(n_362), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B1(n_372), .B2(n_375), .C(n_376), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g387 ( .A(n_367), .Y(n_387) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_379), .B(n_382), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_388), .C(n_389), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_389) );
CKINVDCx14_ASAP7_75t_R g399 ( .A(n_393), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_409), .C(n_417), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B1(n_400), .B2(n_401), .C(n_403), .Y(n_395) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g732 ( .A(n_429), .Y(n_732) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g733 ( .A(n_432), .Y(n_733) );
AND3x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_628), .C(n_685), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_573), .C(n_609), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_482), .B(n_528), .C(n_560), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_455), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g531 ( .A(n_437), .B(n_532), .Y(n_531) );
INVx5_ASAP7_75t_L g559 ( .A(n_437), .Y(n_559) );
AND2x2_ASAP7_75t_L g632 ( .A(n_437), .B(n_548), .Y(n_632) );
AND2x2_ASAP7_75t_L g670 ( .A(n_437), .B(n_576), .Y(n_670) );
AND2x2_ASAP7_75t_L g690 ( .A(n_437), .B(n_533), .Y(n_690) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_452), .Y(n_437) );
AOI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_443), .B(n_451), .Y(n_438) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx5_ASAP7_75t_L g475 ( .A(n_444), .Y(n_475) );
INVx2_ASAP7_75t_L g450 ( .A(n_448), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_450), .A2(n_477), .B(n_478), .C(n_479), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_450), .A2(n_479), .B(n_512), .C(n_513), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_455), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_470), .Y(n_455) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_456), .Y(n_571) );
AND2x2_ASAP7_75t_L g585 ( .A(n_456), .B(n_532), .Y(n_585) );
INVx1_ASAP7_75t_L g608 ( .A(n_456), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_456), .B(n_559), .Y(n_647) );
OR2x2_ASAP7_75t_L g684 ( .A(n_456), .B(n_530), .Y(n_684) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_457), .Y(n_620) );
AND2x2_ASAP7_75t_L g627 ( .A(n_457), .B(n_533), .Y(n_627) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g548 ( .A(n_458), .B(n_533), .Y(n_548) );
BUFx2_ASAP7_75t_L g576 ( .A(n_458), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_466), .A2(n_475), .B(n_521), .C(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_466), .A2(n_475), .B(n_536), .C(n_537), .Y(n_535) );
INVx5_ASAP7_75t_L g530 ( .A(n_470), .Y(n_530) );
BUFx2_ASAP7_75t_L g552 ( .A(n_470), .Y(n_552) );
AND2x2_ASAP7_75t_L g709 ( .A(n_470), .B(n_563), .Y(n_709) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_515), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_484), .A2(n_610), .B1(n_617), .B2(n_618), .C(n_621), .Y(n_609) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
AND2x2_ASAP7_75t_L g516 ( .A(n_485), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_485), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g544 ( .A(n_486), .B(n_495), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_486), .B(n_496), .Y(n_554) );
OR2x2_ASAP7_75t_L g565 ( .A(n_486), .B(n_517), .Y(n_565) );
AND2x2_ASAP7_75t_L g568 ( .A(n_486), .B(n_556), .Y(n_568) );
AND2x2_ASAP7_75t_L g584 ( .A(n_486), .B(n_506), .Y(n_584) );
OR2x2_ASAP7_75t_L g600 ( .A(n_486), .B(n_496), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_486), .B(n_517), .Y(n_662) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_487), .B(n_506), .Y(n_654) );
AND2x2_ASAP7_75t_L g657 ( .A(n_487), .B(n_496), .Y(n_657) );
OR2x2_ASAP7_75t_L g578 ( .A(n_494), .B(n_565), .Y(n_578) );
INVx2_ASAP7_75t_L g604 ( .A(n_494), .Y(n_604) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
AND2x2_ASAP7_75t_L g527 ( .A(n_495), .B(n_507), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_495), .B(n_517), .Y(n_583) );
OR2x2_ASAP7_75t_L g594 ( .A(n_495), .B(n_507), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_495), .B(n_556), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_495), .A2(n_687), .B1(n_689), .B2(n_691), .C(n_694), .Y(n_686) );
INVx5_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_496), .B(n_517), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_506), .B(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_506), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g572 ( .A(n_506), .B(n_544), .Y(n_572) );
OR2x2_ASAP7_75t_L g616 ( .A(n_506), .B(n_517), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_506), .B(n_568), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_506), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g681 ( .A(n_506), .B(n_682), .Y(n_681) );
INVx5_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_507), .B(n_516), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_507), .A2(n_550), .B(n_553), .C(n_557), .Y(n_549) );
OR2x2_ASAP7_75t_L g587 ( .A(n_507), .B(n_583), .Y(n_587) );
OR2x2_ASAP7_75t_L g623 ( .A(n_507), .B(n_565), .Y(n_623) );
OAI311xp33_ASAP7_75t_L g629 ( .A1(n_507), .A2(n_568), .A3(n_630), .B1(n_633), .C1(n_640), .Y(n_629) );
AND2x2_ASAP7_75t_L g680 ( .A(n_507), .B(n_517), .Y(n_680) );
AND2x2_ASAP7_75t_L g688 ( .A(n_507), .B(n_543), .Y(n_688) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_507), .Y(n_706) );
AND2x2_ASAP7_75t_L g723 ( .A(n_507), .B(n_544), .Y(n_723) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_527), .Y(n_515) );
AND2x2_ASAP7_75t_L g551 ( .A(n_516), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g707 ( .A(n_516), .Y(n_707) );
AND2x2_ASAP7_75t_L g543 ( .A(n_517), .B(n_544), .Y(n_543) );
INVx3_ASAP7_75t_L g556 ( .A(n_517), .Y(n_556) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_517), .Y(n_599) );
INVxp67_ASAP7_75t_L g638 ( .A(n_517), .Y(n_638) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_517) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_526), .A2(n_534), .B(n_542), .Y(n_533) );
AND2x2_ASAP7_75t_L g716 ( .A(n_527), .B(n_564), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_543), .B1(n_545), .B2(n_546), .C(n_549), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_530), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g569 ( .A(n_530), .B(n_559), .Y(n_569) );
AND2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_532), .Y(n_577) );
OR2x2_ASAP7_75t_L g589 ( .A(n_530), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g607 ( .A(n_530), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g631 ( .A(n_530), .B(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_530), .Y(n_651) );
AND2x2_ASAP7_75t_L g703 ( .A(n_530), .B(n_627), .Y(n_703) );
OAI31xp33_ASAP7_75t_L g711 ( .A1(n_530), .A2(n_580), .A3(n_679), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_531), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g675 ( .A(n_531), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_531), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g563 ( .A(n_532), .B(n_559), .Y(n_563) );
INVx1_ASAP7_75t_L g650 ( .A(n_532), .Y(n_650) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g700 ( .A(n_533), .B(n_559), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_SL g710 ( .A(n_543), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_544), .B(n_615), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_545), .A2(n_657), .B1(n_695), .B2(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g558 ( .A(n_548), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g617 ( .A(n_548), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_548), .B(n_569), .Y(n_722) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g692 ( .A(n_551), .B(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_552), .A2(n_611), .B(n_613), .Y(n_610) );
OR2x2_ASAP7_75t_L g618 ( .A(n_552), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g639 ( .A(n_552), .B(n_627), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_552), .B(n_650), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_552), .B(n_690), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g666 ( .A1(n_553), .A2(n_667), .B1(n_672), .B2(n_675), .C(n_676), .Y(n_666) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OR2x2_ASAP7_75t_L g643 ( .A(n_554), .B(n_616), .Y(n_643) );
INVx1_ASAP7_75t_L g682 ( .A(n_554), .Y(n_682) );
INVx2_ASAP7_75t_L g658 ( .A(n_555), .Y(n_658) );
INVx1_ASAP7_75t_L g592 ( .A(n_556), .Y(n_592) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g597 ( .A(n_559), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_559), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g626 ( .A(n_559), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g714 ( .A(n_559), .B(n_684), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B1(n_566), .B2(n_569), .C1(n_570), .C2(n_572), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g570 ( .A(n_563), .B(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_563), .A2(n_613), .B1(n_641), .B2(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_563), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OAI21xp33_ASAP7_75t_SL g601 ( .A1(n_572), .A2(n_602), .B(n_605), .Y(n_601) );
OAI211xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_578), .B(n_579), .C(n_601), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_577), .A2(n_580), .B1(n_585), .B2(n_586), .C(n_588), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_577), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g671 ( .A(n_577), .Y(n_671) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g673 ( .A(n_582), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g590 ( .A(n_585), .Y(n_590) );
AND2x2_ASAP7_75t_L g596 ( .A(n_585), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B1(n_595), .B2(n_598), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_592), .B(n_604), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_593), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g693 ( .A(n_597), .Y(n_693) );
AND2x2_ASAP7_75t_L g712 ( .A(n_597), .B(n_627), .Y(n_712) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_604), .B(n_661), .Y(n_720) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_607), .B(n_675), .Y(n_718) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g641 ( .A(n_619), .Y(n_641) );
BUFx2_ASAP7_75t_L g665 ( .A(n_620), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_624), .B(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_644), .C(n_666), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_648), .B(n_652), .C(n_655), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_645), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NOR2xp67_ASAP7_75t_SL g649 ( .A(n_650), .B(n_651), .Y(n_649) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_SL g674 ( .A(n_654), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B(n_663), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AND2x2_ASAP7_75t_L g679 ( .A(n_657), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B1(n_681), .B2(n_683), .Y(n_676) );
INVx2_ASAP7_75t_SL g697 ( .A(n_684), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_701), .C(n_713), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_697), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_708), .B2(n_710), .C(n_711), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_702), .A2(n_714), .B(n_715), .C(n_717), .Y(n_713) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_721), .B2(n_723), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g734 ( .A(n_725), .Y(n_734) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_730) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_SL g751 ( .A(n_741), .Y(n_751) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g748 ( .A(n_745), .Y(n_748) );
BUFx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
endmodule