module fake_jpeg_1950_n_494 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g112 ( 
.A(n_48),
.Y(n_112)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_51),
.Y(n_135)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_39),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_95),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_41),
.Y(n_102)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_22),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_27),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_20),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_101),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_146),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_21),
.B1(n_28),
.B2(n_25),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_107),
.A2(n_143),
.B1(n_24),
.B2(n_26),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_60),
.A2(n_16),
.B1(n_41),
.B2(n_45),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_131),
.B1(n_149),
.B2(n_154),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_63),
.A2(n_16),
.B1(n_41),
.B2(n_32),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_38),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_145),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_65),
.A2(n_40),
.B1(n_32),
.B2(n_35),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_55),
.B(n_23),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_45),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_66),
.A2(n_37),
.B1(n_23),
.B2(n_35),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_47),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_109),
.A2(n_75),
.B1(n_93),
.B2(n_92),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_157),
.A2(n_168),
.B1(n_170),
.B2(n_184),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_158),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_22),
.B1(n_88),
.B2(n_81),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_160),
.A2(n_172),
.B1(n_182),
.B2(n_196),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_118),
.A2(n_40),
.B1(n_67),
.B2(n_97),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_162),
.A2(n_179),
.B1(n_183),
.B2(n_140),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_112),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_165),
.Y(n_235)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_84),
.B1(n_49),
.B2(n_68),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_185),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_78),
.B1(n_74),
.B2(n_73),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_103),
.B(n_48),
.C(n_69),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_114),
.C(n_122),
.Y(n_206)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_178),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_40),
.B1(n_25),
.B2(n_33),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_107),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_136),
.A2(n_33),
.B1(n_83),
.B2(n_91),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_107),
.A2(n_125),
.B1(n_116),
.B2(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_106),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_188),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_105),
.A2(n_48),
.A3(n_69),
.B1(n_72),
.B2(n_51),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_32),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_198),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_129),
.A2(n_91),
.B1(n_83),
.B2(n_35),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_200),
.B1(n_104),
.B2(n_133),
.Y(n_234)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_119),
.A2(n_85),
.B1(n_21),
.B2(n_35),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_0),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_129),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_142),
.B(n_1),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_116),
.B1(n_148),
.B2(n_144),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_204),
.A2(n_185),
.B1(n_192),
.B2(n_190),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_171),
.C(n_165),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_209),
.A2(n_214),
.B1(n_224),
.B2(n_193),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_163),
.A2(n_153),
.B1(n_147),
.B2(n_121),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_161),
.A2(n_111),
.B1(n_155),
.B2(n_99),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_234),
.B1(n_157),
.B2(n_200),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_151),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_231),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_163),
.A2(n_122),
.B1(n_104),
.B2(n_113),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_155),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_139),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_184),
.Y(n_241)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_191),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_241),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_257),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_232),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_243),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_195),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_181),
.B(n_201),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_244),
.A2(n_240),
.B(n_264),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_195),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_217),
.B(n_195),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_174),
.C(n_186),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_252),
.C(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_207),
.B(n_186),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_250),
.B(n_264),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_227),
.B(n_207),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_237),
.B(n_233),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_156),
.C(n_177),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_227),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_254),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_218),
.B(n_164),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_215),
.A2(n_161),
.B1(n_172),
.B2(n_181),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_267),
.B1(n_203),
.B2(n_132),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_202),
.Y(n_259)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_212),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_211),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_216),
.A2(n_170),
.B1(n_181),
.B2(n_196),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_263),
.A2(n_126),
.B1(n_99),
.B2(n_169),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_188),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_235),
.B1(n_213),
.B2(n_234),
.Y(n_265)
);

AO21x2_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_199),
.B(n_228),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_192),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_204),
.A2(n_132),
.B1(n_139),
.B2(n_126),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

AO22x1_ASAP7_75t_SL g270 ( 
.A1(n_256),
.A2(n_213),
.B1(n_236),
.B2(n_203),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_270),
.B(n_279),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_284),
.B1(n_286),
.B2(n_292),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_261),
.C(n_242),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_283),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_277),
.A2(n_289),
.B(n_290),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_245),
.A3(n_242),
.B1(n_252),
.B2(n_238),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_225),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_282),
.B(n_272),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_212),
.C(n_226),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_285),
.A2(n_275),
.B1(n_263),
.B2(n_287),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_228),
.B1(n_219),
.B2(n_229),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_295),
.B1(n_239),
.B2(n_263),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_233),
.B(n_219),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_229),
.B(n_223),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_226),
.C(n_223),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_293),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_180),
.B1(n_178),
.B2(n_220),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_230),
.C(n_220),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_244),
.B(n_243),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_239),
.A2(n_230),
.B1(n_205),
.B2(n_211),
.Y(n_295)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_252),
.B(n_244),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_245),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_305),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_260),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_254),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_306),
.B(n_309),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_SL g349 ( 
.A(n_307),
.B(n_286),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_257),
.B(n_250),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_318),
.B(n_285),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_255),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_311),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_290),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_323),
.B1(n_285),
.B2(n_205),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_281),
.B(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_319),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_277),
.A2(n_271),
.B(n_281),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_246),
.C(n_276),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_271),
.A2(n_260),
.B1(n_241),
.B2(n_267),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_313),
.B1(n_314),
.B2(n_321),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_259),
.B1(n_266),
.B2(n_248),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_321),
.A2(n_285),
.B1(n_295),
.B2(n_284),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_322),
.B(n_292),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_278),
.A2(n_285),
.B1(n_288),
.B2(n_270),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_284),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_325),
.Y(n_341)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_282),
.C(n_272),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_335),
.C(n_338),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_293),
.C(n_279),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_336),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_337),
.A2(n_349),
.B(n_327),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_299),
.C(n_270),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_247),
.C(n_268),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_358),
.C(n_307),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_344),
.B(n_346),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_304),
.B(n_315),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_348),
.A2(n_356),
.B1(n_258),
.B2(n_175),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_351),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_222),
.Y(n_353)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_303),
.B(n_305),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_355),
.B(n_300),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_222),
.B1(n_258),
.B2(n_176),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_222),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_361),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_197),
.C(n_194),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_310),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_306),
.Y(n_365)
);

AOI21xp33_ASAP7_75t_L g361 ( 
.A1(n_308),
.A2(n_258),
.B(n_159),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_309),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_362),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_369),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_380),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_367),
.A2(n_368),
.B(n_371),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_337),
.A2(n_318),
.B(n_327),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_341),
.A2(n_311),
.B(n_325),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_329),
.C(n_317),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_377),
.C(n_379),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_329),
.B(n_320),
.Y(n_371)
);

AO21x1_ASAP7_75t_L g372 ( 
.A1(n_352),
.A2(n_314),
.B(n_328),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_349),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_382),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_324),
.C(n_330),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_378),
.A2(n_387),
.B1(n_336),
.B2(n_359),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_173),
.C(n_167),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_14),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_342),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_381)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_12),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_348),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_383),
.A2(n_389),
.B1(n_343),
.B2(n_354),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_0),
.C(n_1),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_388),
.C(n_346),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_333),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_386),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_11),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_358),
.C(n_345),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_342),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_390),
.B(n_392),
.Y(n_429)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_391),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_350),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_365),
.B(n_332),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_399),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_343),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_397),
.Y(n_417)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_403),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_345),
.C(n_334),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_404),
.C(n_409),
.Y(n_421)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_411),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_334),
.C(n_332),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_356),
.C(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_387),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_383),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_354),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_347),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_412),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_372),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_10),
.Y(n_432)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_388),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_418),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_406),
.A2(n_375),
.B1(n_370),
.B2(n_385),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_400),
.A2(n_412),
.B1(n_391),
.B2(n_409),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_420),
.Y(n_440)
);

NAND2xp67_ASAP7_75t_SL g420 ( 
.A(n_407),
.B(n_367),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_397),
.A2(n_368),
.B1(n_382),
.B2(n_374),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_425),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_407),
.A2(n_364),
.B1(n_347),
.B2(n_360),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_404),
.A2(n_389),
.B1(n_360),
.B2(n_380),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_395),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_403),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_401),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_393),
.A2(n_364),
.B(n_386),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_431),
.A2(n_405),
.B(n_408),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_432),
.A2(n_410),
.B(n_399),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_439),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_438),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_398),
.C(n_411),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_423),
.A2(n_405),
.B(n_408),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_429),
.B(n_398),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_441),
.B(n_427),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_449),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_395),
.C(n_5),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_SL g456 ( 
.A(n_443),
.B(n_446),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_444),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_11),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_445),
.B(n_424),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_3),
.C(n_5),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_428),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_415),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_417),
.A2(n_5),
.B(n_6),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_448),
.A2(n_425),
.B1(n_430),
.B2(n_433),
.Y(n_460)
);

FAx1_ASAP7_75t_SL g449 ( 
.A(n_420),
.B(n_5),
.CI(n_6),
.CON(n_449),
.SN(n_449)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_437),
.A2(n_418),
.B(n_416),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_451),
.B(n_454),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_452),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_440),
.A2(n_424),
.B(n_417),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_458),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_438),
.B(n_443),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_460),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_415),
.C(n_433),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_462),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_426),
.C(n_422),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_431),
.C(n_414),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_435),
.C(n_450),
.Y(n_468)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_436),
.C(n_446),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_471),
.Y(n_482)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_442),
.B(n_448),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_470),
.A2(n_7),
.B(n_9),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_461),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_449),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_472),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_449),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_475),
.B(n_465),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g485 ( 
.A1(n_477),
.A2(n_478),
.B(n_473),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_473),
.A2(n_457),
.B1(n_452),
.B2(n_463),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_456),
.C(n_7),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_479),
.B(n_7),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g484 ( 
.A1(n_481),
.A2(n_474),
.B(n_466),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_484),
.Y(n_489)
);

AO21x1_ASAP7_75t_L g490 ( 
.A1(n_485),
.A2(n_486),
.B(n_487),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_482),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_483),
.C(n_468),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_488),
.B(n_467),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_490),
.B(n_480),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_480),
.C(n_489),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_472),
.Y(n_494)
);


endmodule