module real_aes_10657_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_884, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_884;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_880;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g582 ( .A(n_0), .B(n_158), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_1), .A2(n_86), .B1(n_151), .B2(n_153), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_2), .B(n_168), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_3), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_4), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_5), .B(n_201), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_6), .A2(n_41), .B1(n_145), .B2(n_180), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_7), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_8), .B(n_153), .Y(n_626) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g120 ( .A(n_9), .B(n_89), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_10), .B(n_180), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_11), .B(n_143), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_12), .A2(n_64), .B1(n_178), .B2(n_180), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g250 ( .A(n_13), .B(n_180), .C(n_197), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_14), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_15), .Y(n_881) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_16), .B(n_180), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_17), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_18), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_19), .B(n_152), .Y(n_210) );
NAND3xp33_ASAP7_75t_L g245 ( .A(n_20), .B(n_143), .C(n_149), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_21), .B(n_180), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_22), .A2(n_29), .B1(n_143), .B2(n_145), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_23), .B(n_212), .Y(n_266) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_24), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_25), .B(n_153), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_26), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_27), .B(n_192), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_28), .B(n_540), .Y(n_568) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_30), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_31), .B(n_143), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_32), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_33), .B(n_564), .Y(n_563) );
NAND2xp33_ASAP7_75t_SL g538 ( .A(n_34), .B(n_152), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_35), .A2(n_54), .B1(n_178), .B2(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_36), .B(n_183), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_37), .B(n_149), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_38), .B(n_265), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_39), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g119 ( .A(n_39), .Y(n_119) );
OAI21x1_ASAP7_75t_L g160 ( .A1(n_40), .A2(n_69), .B(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_42), .A2(n_132), .B1(n_133), .B2(n_516), .Y(n_131) );
INVx1_ASAP7_75t_L g516 ( .A(n_42), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_42), .A2(n_82), .B1(n_516), .B2(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_43), .B(n_183), .Y(n_613) );
AND2x2_ASAP7_75t_L g182 ( .A(n_44), .B(n_183), .Y(n_182) );
AND2x6_ASAP7_75t_L g164 ( .A(n_45), .B(n_165), .Y(n_164) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_46), .B(n_183), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_47), .B(n_531), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_48), .B(n_531), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_49), .B(n_597), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_50), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_51), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_52), .B(n_152), .Y(n_268) );
INVx1_ASAP7_75t_L g165 ( .A(n_53), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_55), .B(n_178), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_56), .B(n_183), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_57), .B(n_143), .Y(n_217) );
NAND2xp33_ASAP7_75t_L g536 ( .A(n_58), .B(n_152), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_59), .A2(n_129), .B1(n_130), .B2(n_858), .Y(n_128) );
INVx1_ASAP7_75t_L g858 ( .A(n_59), .Y(n_858) );
AND2x2_ASAP7_75t_L g108 ( .A(n_60), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_61), .B(n_143), .Y(n_199) );
NAND2x1_ASAP7_75t_L g273 ( .A(n_62), .B(n_183), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_63), .B(n_197), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_65), .B(n_540), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_66), .B(n_235), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_67), .B(n_179), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_68), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_70), .B(n_143), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_71), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_72), .B(n_197), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_73), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_74), .B(n_597), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_75), .A2(n_79), .B1(n_143), .B2(n_145), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_76), .B(n_183), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_77), .Y(n_233) );
BUFx10_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
INVx1_ASAP7_75t_SL g169 ( .A(n_80), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_81), .Y(n_298) );
INVx1_ASAP7_75t_L g868 ( .A(n_82), .Y(n_868) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_83), .B(n_143), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_84), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_85), .B(n_145), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_87), .B(n_264), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_88), .B(n_180), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_89), .B(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g161 ( .A(n_90), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_91), .B(n_197), .Y(n_247) );
INVx1_ASAP7_75t_L g110 ( .A(n_92), .Y(n_110) );
OR2x2_ASAP7_75t_L g116 ( .A(n_92), .B(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g519 ( .A(n_92), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_92), .B(n_118), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_93), .B(n_231), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_94), .B(n_564), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_95), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g109 ( .A(n_96), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_97), .B(n_153), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_98), .B(n_146), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_99), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_111), .B(n_880), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx3_ASAP7_75t_L g882 ( .A(n_103), .Y(n_882) );
AND2x6_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_110), .Y(n_107) );
OR2x6_ASAP7_75t_L g111 ( .A(n_112), .B(n_121), .Y(n_111) );
INVx1_ASAP7_75t_L g873 ( .A(n_112), .Y(n_873) );
NOR2xp67_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .Y(n_112) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx4_ASAP7_75t_L g865 ( .A(n_115), .Y(n_865) );
INVx5_ASAP7_75t_L g872 ( .A(n_115), .Y(n_872) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x6_ASAP7_75t_L g125 ( .A(n_118), .B(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI21x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_128), .B(n_859), .Y(n_121) );
INVx2_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx12f_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g878 ( .A(n_126), .B(n_879), .Y(n_878) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
BUFx12f_ASAP7_75t_L g861 ( .A(n_127), .Y(n_861) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_517), .B(n_520), .Y(n_130) );
INVx2_ASAP7_75t_SL g869 ( .A(n_132), .Y(n_869) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_421), .Y(n_133) );
NAND4xp25_ASAP7_75t_L g134 ( .A(n_135), .B(n_325), .C(n_372), .D(n_409), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_257), .B(n_274), .Y(n_135) );
AO22x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_204), .B1(n_236), .B2(n_256), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_185), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_138), .B(n_186), .Y(n_338) );
AND2x2_ASAP7_75t_L g441 ( .A(n_138), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_139), .B(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g477 ( .A(n_139), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_170), .Y(n_139) );
AND2x2_ASAP7_75t_L g252 ( .A(n_140), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g281 ( .A(n_140), .Y(n_281) );
INVx1_ASAP7_75t_L g304 ( .A(n_140), .Y(n_304) );
INVx1_ASAP7_75t_L g334 ( .A(n_140), .Y(n_334) );
AO31x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_157), .A3(n_162), .B(n_166), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B1(n_150), .B2(n_155), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_143), .A2(n_195), .B(n_196), .C(n_197), .Y(n_194) );
OAI321xp33_ASAP7_75t_L g222 ( .A1(n_143), .A2(n_149), .A3(n_151), .B1(n_223), .B2(n_224), .C(n_225), .Y(n_222) );
INVx2_ASAP7_75t_SL g249 ( .A(n_143), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_143), .A2(n_265), .B1(n_577), .B2(n_578), .Y(n_576) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_144), .Y(n_146) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
INVx1_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
INVx2_ASAP7_75t_L g265 ( .A(n_144), .Y(n_265) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g201 ( .A(n_146), .Y(n_201) );
INVx2_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
INVx2_ASAP7_75t_L g540 ( .A(n_146), .Y(n_540) );
INVx2_ASAP7_75t_L g564 ( .A(n_146), .Y(n_564) );
OA22x2_ASAP7_75t_L g175 ( .A1(n_147), .A2(n_155), .B1(n_176), .B2(n_177), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_147), .A2(n_293), .B1(n_294), .B2(n_295), .Y(n_292) );
CKINVDCx6p67_ASAP7_75t_R g147 ( .A(n_148), .Y(n_147) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_148), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_148), .A2(n_227), .B(n_232), .Y(n_226) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_148), .A2(n_263), .B(n_266), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_148), .A2(n_534), .B(n_535), .C(n_536), .Y(n_533) );
INVx2_ASAP7_75t_SL g541 ( .A(n_148), .Y(n_541) );
INVx2_ASAP7_75t_SL g552 ( .A(n_148), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_148), .A2(n_563), .B(n_565), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_148), .A2(n_596), .B(n_598), .Y(n_595) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx12f_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx5_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_149), .A2(n_214), .B1(n_215), .B2(n_217), .Y(n_213) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g216 ( .A(n_152), .Y(n_216) );
INVx2_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_152), .B(n_233), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_153), .A2(n_197), .B(n_586), .C(n_587), .Y(n_585) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_156), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21x1_ASAP7_75t_L g267 ( .A1(n_156), .A2(n_268), .B(n_269), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_156), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_156), .A2(n_580), .B(n_581), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_156), .A2(n_589), .B(n_590), .Y(n_588) );
INVx3_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g240 ( .A(n_158), .Y(n_240) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_158), .Y(n_254) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_158), .A2(n_584), .B(n_591), .Y(n_583) );
BUFx4f_ASAP7_75t_L g602 ( .A(n_158), .Y(n_602) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_159), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
AND2x2_ASAP7_75t_L g291 ( .A(n_162), .B(n_240), .Y(n_291) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_162), .A2(n_562), .B(n_566), .Y(n_561) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_162), .A2(n_621), .B(n_624), .Y(n_620) );
INVx8_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_163), .A2(n_225), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_SL g542 ( .A(n_163), .Y(n_542) );
INVx8_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_164), .A2(n_209), .B(n_213), .Y(n_208) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_164), .A2(n_242), .B(n_246), .Y(n_241) );
BUFx2_ASAP7_75t_L g272 ( .A(n_164), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_164), .A2(n_541), .B(n_576), .C(n_579), .Y(n_575) );
OAI21x1_ASAP7_75t_SL g584 ( .A1(n_164), .A2(n_585), .B(n_588), .Y(n_584) );
OAI21x1_ASAP7_75t_L g606 ( .A1(n_164), .A2(n_607), .B(n_610), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
INVx1_ASAP7_75t_L g192 ( .A(n_167), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_167), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_SL g531 ( .A(n_167), .Y(n_531) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx5_ASAP7_75t_L g173 ( .A(n_168), .Y(n_173) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_168), .Y(n_235) );
INVx1_ASAP7_75t_L g332 ( .A(n_170), .Y(n_332) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_170), .Y(n_350) );
INVx1_ASAP7_75t_L g377 ( .A(n_170), .Y(n_377) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_170), .Y(n_407) );
INVx1_ASAP7_75t_L g456 ( .A(n_170), .Y(n_456) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_175), .B(n_181), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_174), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI21x1_ASAP7_75t_L g547 ( .A1(n_173), .A2(n_548), .B(n_557), .Y(n_547) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_173), .A2(n_561), .B(n_569), .Y(n_560) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_173), .A2(n_575), .B(n_582), .Y(n_574) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_173), .A2(n_620), .B(n_627), .Y(n_619) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_175), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx5_ASAP7_75t_L g597 ( .A(n_180), .Y(n_597) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVxp67_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g472 ( .A(n_186), .B(n_252), .Y(n_472) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp67_ASAP7_75t_L g303 ( .A(n_187), .B(n_304), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_187), .B(n_376), .C(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g455 ( .A(n_187), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g277 ( .A(n_188), .B(n_253), .Y(n_277) );
AND2x2_ASAP7_75t_L g378 ( .A(n_188), .B(n_342), .Y(n_378) );
AND2x2_ASAP7_75t_L g386 ( .A(n_188), .B(n_304), .Y(n_386) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g336 ( .A(n_189), .B(n_238), .Y(n_336) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g310 ( .A(n_190), .Y(n_310) );
AND2x2_ASAP7_75t_L g420 ( .A(n_190), .B(n_238), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_198), .B(n_202), .Y(n_193) );
O2A1O1Ixp5_ASAP7_75t_L g553 ( .A1(n_197), .A2(n_554), .B(n_555), .C(n_556), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_197), .A2(n_608), .B(n_609), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_197), .A2(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g555 ( .A(n_201), .Y(n_555) );
AND2x2_ASAP7_75t_L g413 ( .A(n_204), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_219), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_205), .B(n_323), .Y(n_328) );
INVx1_ASAP7_75t_L g396 ( .A(n_205), .Y(n_396) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g285 ( .A(n_206), .Y(n_285) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_218), .Y(n_206) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_207), .A2(n_261), .B(n_273), .Y(n_260) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_207), .A2(n_261), .B(n_273), .Y(n_322) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_207), .A2(n_208), .B(n_218), .Y(n_357) );
INVxp67_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_216), .B(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g256 ( .A(n_219), .Y(n_256) );
AND2x4_ASAP7_75t_L g438 ( .A(n_219), .B(n_383), .Y(n_438) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_220), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g390 ( .A(n_220), .B(n_322), .Y(n_390) );
AND2x2_ASAP7_75t_L g504 ( .A(n_220), .B(n_399), .Y(n_504) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g288 ( .A(n_221), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g301 ( .A(n_221), .Y(n_301) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_226), .B(n_234), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI32xp33_ASAP7_75t_L g313 ( .A1(n_236), .A2(n_307), .A3(n_314), .B1(n_315), .B2(n_318), .Y(n_313) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_252), .Y(n_236) );
NOR2xp67_ASAP7_75t_L g278 ( .A(n_237), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_237), .B(n_334), .Y(n_371) );
OAI32xp33_ASAP7_75t_L g423 ( .A1(n_237), .A2(n_331), .A3(n_424), .B1(n_427), .B2(n_429), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_237), .B(n_324), .C(n_459), .Y(n_458) );
BUFx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_241), .B(n_251), .Y(n_238) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_239), .A2(n_241), .B(n_251), .Y(n_306) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_245), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_250), .Y(n_246) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_252), .B(n_408), .Y(n_513) );
AND2x2_ASAP7_75t_L g305 ( .A(n_253), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g314 ( .A(n_256), .Y(n_314) );
INVx1_ASAP7_75t_L g482 ( .A(n_256), .Y(n_482) );
OR2x2_ASAP7_75t_L g509 ( .A(n_257), .B(n_425), .Y(n_509) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g283 ( .A(n_258), .B(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g329 ( .A(n_258), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_258), .B(n_284), .Y(n_426) );
AND2x2_ASAP7_75t_L g448 ( .A(n_258), .B(n_349), .Y(n_448) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g312 ( .A(n_259), .B(n_289), .Y(n_312) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_259), .Y(n_502) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g364 ( .A(n_260), .Y(n_364) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_267), .B(n_272), .Y(n_261) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g296 ( .A(n_265), .Y(n_296) );
INVx1_ASAP7_75t_L g535 ( .A(n_265), .Y(n_535) );
INVx4_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_313), .Y(n_274) );
AOI322xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_282), .A3(n_286), .B1(n_299), .B2(n_302), .C1(n_307), .C2(n_311), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g370 ( .A(n_277), .Y(n_370) );
AND2x2_ASAP7_75t_L g497 ( .A(n_277), .B(n_341), .Y(n_497) );
INVxp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g486 ( .A(n_280), .B(n_310), .Y(n_486) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g309 ( .A(n_281), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g341 ( .A(n_281), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_283), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g490 ( .A(n_284), .B(n_395), .Y(n_490) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_SL g324 ( .A(n_285), .Y(n_324) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_287), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g382 ( .A(n_288), .B(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g446 ( .A(n_288), .Y(n_446) );
AND2x2_ASAP7_75t_L g467 ( .A(n_288), .B(n_384), .Y(n_467) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
INVx2_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g399 ( .A(n_290), .Y(n_399) );
AOI21x1_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_297), .Y(n_290) );
AND2x2_ASAP7_75t_L g356 ( .A(n_301), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g367 ( .A(n_301), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g425 ( .A(n_301), .B(n_399), .Y(n_425) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_301), .Y(n_440) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g417 ( .A(n_304), .Y(n_417) );
AND2x4_ASAP7_75t_L g485 ( .A(n_305), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_305), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g342 ( .A(n_306), .Y(n_342) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
AND2x2_ASAP7_75t_L g387 ( .A(n_309), .B(n_377), .Y(n_387) );
BUFx2_ASAP7_75t_L g450 ( .A(n_309), .Y(n_450) );
INVx1_ASAP7_75t_L g507 ( .A(n_309), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_310), .B(n_342), .Y(n_393) );
INVx2_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_316), .A2(n_386), .B1(n_455), .B2(n_457), .C(n_458), .Y(n_454) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_317), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g457 ( .A(n_317), .Y(n_457) );
INVx1_ASAP7_75t_L g346 ( .A(n_318), .Y(n_346) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
INVx2_ASAP7_75t_L g431 ( .A(n_320), .Y(n_431) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx2_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g360 ( .A(n_323), .Y(n_360) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_323), .Y(n_389) );
AND2x2_ASAP7_75t_L g343 ( .A(n_324), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g379 ( .A(n_324), .B(n_358), .Y(n_379) );
AND2x2_ASAP7_75t_L g463 ( .A(n_324), .B(n_366), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_330), .B1(n_337), .B2(n_343), .C(n_345), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_328), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
OR2x2_ASAP7_75t_L g339 ( .A(n_331), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g427 ( .A(n_331), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g385 ( .A(n_332), .B(n_386), .Y(n_385) );
NOR2x1_ASAP7_75t_L g481 ( .A(n_332), .B(n_417), .Y(n_481) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g353 ( .A(n_334), .Y(n_353) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_334), .Y(n_374) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g400 ( .A(n_336), .B(n_377), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NOR2x1p5_ASAP7_75t_L g487 ( .A(n_340), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g349 ( .A(n_342), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_344), .B(n_356), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_352), .B2(n_354), .C(n_361), .Y(n_345) );
OAI222xp33_ASAP7_75t_L g510 ( .A1(n_347), .A2(n_412), .B1(n_511), .B2(n_512), .C1(n_513), .C2(n_514), .Y(n_510) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
OR2x2_ASAP7_75t_L g352 ( .A(n_348), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
OR2x6_ASAP7_75t_L g495 ( .A(n_351), .B(n_456), .Y(n_495) );
INVx2_ASAP7_75t_L g468 ( .A(n_352), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_355), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g368 ( .A(n_357), .Y(n_368) );
INVx2_ASAP7_75t_L g384 ( .A(n_357), .Y(n_384) );
INVx1_ASAP7_75t_L g412 ( .A(n_358), .Y(n_412) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g366 ( .A(n_359), .Y(n_366) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_359), .Y(n_414) );
AND2x2_ASAP7_75t_L g479 ( .A(n_359), .B(n_378), .Y(n_479) );
AND2x2_ASAP7_75t_L g395 ( .A(n_360), .B(n_364), .Y(n_395) );
OAI21xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_369), .Y(n_361) );
BUFx2_ASAP7_75t_L g453 ( .A(n_364), .Y(n_453) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_364), .Y(n_515) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g397 ( .A(n_367), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g430 ( .A(n_367), .Y(n_430) );
NOR2x1p5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AOI211xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_379), .B(n_380), .C(n_401), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx2_ASAP7_75t_L g466 ( .A(n_375), .Y(n_466) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
AO22x1_ASAP7_75t_L g480 ( .A1(n_376), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_480) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
AND2x2_ASAP7_75t_L g491 ( .A(n_378), .B(n_477), .Y(n_491) );
INVx1_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
NAND2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_391), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B1(n_387), .B2(n_388), .Y(n_381) );
INVx2_ASAP7_75t_SL g402 ( .A(n_382), .Y(n_402) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g508 ( .A(n_385), .Y(n_508) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g459 ( .A(n_390), .Y(n_459) );
AOI32xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .A3(n_396), .B1(n_397), .B2(n_400), .Y(n_391) );
INVx1_ASAP7_75t_L g408 ( .A(n_393), .Y(n_408) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g434 ( .A(n_395), .Y(n_434) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g465 ( .A(n_400), .Y(n_465) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_404), .Y(n_401) );
OAI321xp33_ASAP7_75t_L g444 ( .A1(n_402), .A2(n_445), .A3(n_447), .B1(n_449), .B2(n_451), .C(n_454), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_406), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_413), .B(n_415), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g443 ( .A(n_420), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_469), .Y(n_421) );
NOR4xp25_ASAP7_75t_L g422 ( .A(n_423), .B(n_432), .C(n_444), .D(n_460), .Y(n_422) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx2_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx2_ASAP7_75t_L g483 ( .A(n_430), .Y(n_483) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_439), .C(n_441), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_436), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx4_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_445), .A2(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_446), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g473 ( .A(n_452), .B(n_467), .Y(n_473) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g488 ( .A(n_455), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_457), .A2(n_462), .B1(n_485), .B2(n_487), .Y(n_484) );
AO22x1_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B1(n_467), .B2(n_468), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g512 ( .A(n_462), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_492), .C(n_510), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_478), .C(n_484), .D(n_489), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_474), .B2(n_476), .Y(n_471) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_490), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g511 ( .A(n_491), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_505), .B1(n_508), .B2(n_509), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx8_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx8_ASAP7_75t_SL g857 ( .A(n_519), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_856), .Y(n_520) );
AND4x1_ASAP7_75t_L g521 ( .A(n_522), .B(n_760), .C(n_802), .D(n_824), .Y(n_521) );
NOR2x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_704), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_648), .C(n_680), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_570), .B1(n_614), .B2(n_629), .C1(n_638), .C2(n_644), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_526), .A2(n_672), .B(n_676), .Y(n_671) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_544), .Y(n_526) );
OR2x2_ASAP7_75t_L g721 ( .A(n_527), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g759 ( .A(n_527), .Y(n_759) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_528), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g714 ( .A(n_528), .B(n_616), .Y(n_714) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g628 ( .A(n_529), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_529), .B(n_643), .Y(n_660) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_529), .Y(n_766) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_530), .Y(n_692) );
AND2x2_ASAP7_75t_L g745 ( .A(n_530), .B(n_617), .Y(n_745) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_543), .Y(n_530) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_531), .A2(n_606), .B(n_613), .Y(n_605) );
OAI21x1_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_537), .B(n_542), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B(n_541), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_541), .A2(n_567), .B(n_568), .Y(n_566) );
AOI21x1_ASAP7_75t_L g599 ( .A1(n_541), .A2(n_600), .B(n_601), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_542), .A2(n_549), .B(n_553), .Y(n_548) );
OAI21x1_ASAP7_75t_L g594 ( .A1(n_542), .A2(n_595), .B(n_599), .Y(n_594) );
INVx1_ASAP7_75t_L g743 ( .A(n_544), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_558), .Y(n_544) );
INVx1_ASAP7_75t_L g717 ( .A(n_545), .Y(n_717) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g639 ( .A(n_546), .B(n_618), .Y(n_639) );
INVx2_ASAP7_75t_L g658 ( .A(n_546), .Y(n_658) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g723 ( .A(n_547), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_552), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_552), .A2(n_611), .B(n_612), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_552), .A2(n_622), .B(n_623), .Y(n_621) );
AND2x2_ASAP7_75t_L g683 ( .A(n_558), .B(n_632), .Y(n_683) );
BUFx2_ASAP7_75t_L g813 ( .A(n_558), .Y(n_813) );
AND2x2_ASAP7_75t_L g849 ( .A(n_558), .B(n_573), .Y(n_849) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx3_ASAP7_75t_L g713 ( .A(n_559), .Y(n_713) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g643 ( .A(n_560), .Y(n_643) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_592), .Y(n_572) );
INVx1_ASAP7_75t_L g843 ( .A(n_573), .Y(n_843) );
AND2x2_ASAP7_75t_L g850 ( .A(n_573), .B(n_664), .Y(n_850) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_583), .Y(n_573) );
INVx3_ASAP7_75t_L g632 ( .A(n_574), .Y(n_632) );
AND2x2_ASAP7_75t_L g645 ( .A(n_574), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g663 ( .A(n_574), .Y(n_663) );
INVx3_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
INVx1_ASAP7_75t_L g741 ( .A(n_592), .Y(n_741) );
INVx2_ASAP7_75t_L g785 ( .A(n_592), .Y(n_785) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_604), .Y(n_592) );
BUFx2_ASAP7_75t_L g635 ( .A(n_593), .Y(n_635) );
AND2x2_ASAP7_75t_L g695 ( .A(n_593), .B(n_605), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_602), .B(n_603), .Y(n_593) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_594), .A2(n_602), .B(n_603), .Y(n_647) );
INVx1_ASAP7_75t_L g633 ( .A(n_604), .Y(n_633) );
NOR2xp67_ASAP7_75t_L g652 ( .A(n_604), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g670 ( .A(n_604), .B(n_637), .Y(n_670) );
AND2x2_ASAP7_75t_L g708 ( .A(n_604), .B(n_709), .Y(n_708) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_604), .Y(n_727) );
INVx1_ASAP7_75t_L g734 ( .A(n_604), .Y(n_734) );
INVx1_ASAP7_75t_L g855 ( .A(n_604), .Y(n_855) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g836 ( .A(n_615), .Y(n_836) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_628), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g668 ( .A(n_618), .B(n_658), .Y(n_668) );
INVx1_ASAP7_75t_L g691 ( .A(n_618), .Y(n_691) );
INVx1_ASAP7_75t_L g719 ( .A(n_618), .Y(n_719) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g675 ( .A(n_628), .Y(n_675) );
AND2x2_ASAP7_75t_L g769 ( .A(n_628), .B(n_643), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_629), .A2(n_639), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
AND2x4_ASAP7_75t_L g700 ( .A(n_630), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_630), .B(n_634), .Y(n_794) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
AND2x2_ASAP7_75t_L g679 ( .A(n_631), .B(n_637), .Y(n_679) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g707 ( .A(n_632), .B(n_646), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_632), .B(n_637), .Y(n_775) );
AND2x2_ASAP7_75t_L g787 ( .A(n_632), .B(n_709), .Y(n_787) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx2_ASAP7_75t_L g678 ( .A(n_635), .Y(n_678) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_635), .Y(n_842) );
INVx1_ASAP7_75t_L g751 ( .A(n_636), .Y(n_751) );
AND2x2_ASAP7_75t_L g825 ( .A(n_636), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g653 ( .A(n_637), .Y(n_653) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_637), .Y(n_694) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_637), .Y(n_702) );
INVx2_ASAP7_75t_SL g709 ( .A(n_637), .Y(n_709) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g768 ( .A(n_639), .B(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g833 ( .A(n_639), .B(n_813), .Y(n_833) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g688 ( .A(n_642), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g722 ( .A(n_642), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2x1_ASAP7_75t_L g726 ( .A(n_645), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g832 ( .A(n_645), .B(n_708), .Y(n_832) );
INVx2_ASAP7_75t_SL g664 ( .A(n_646), .Y(n_664) );
AND2x4_ASAP7_75t_L g733 ( .A(n_646), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_R g703 ( .A(n_647), .Y(n_703) );
NOR2xp33_ASAP7_75t_SL g648 ( .A(n_649), .B(n_671), .Y(n_648) );
OAI31xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_654), .A3(n_661), .B(n_665), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g830 ( .A(n_652), .B(n_707), .Y(n_830) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_653), .Y(n_763) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g749 ( .A(n_658), .Y(n_749) );
AND2x2_ASAP7_75t_L g771 ( .A(n_658), .B(n_719), .Y(n_771) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g698 ( .A(n_660), .Y(n_698) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2x1_ASAP7_75t_L g732 ( .A(n_663), .B(n_733), .Y(n_732) );
INVx4_ASAP7_75t_L g740 ( .A(n_663), .Y(n_740) );
AND2x4_ASAP7_75t_L g669 ( .A(n_664), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g773 ( .A(n_664), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
AND2x2_ASAP7_75t_L g681 ( .A(n_666), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g699 ( .A(n_667), .Y(n_699) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g673 ( .A(n_668), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g765 ( .A(n_668), .B(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g809 ( .A(n_669), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g685 ( .A(n_670), .Y(n_685) );
AND2x2_ASAP7_75t_L g780 ( .A(n_670), .B(n_703), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_670), .B(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g821 ( .A(n_670), .B(n_740), .Y(n_821) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_673), .B(n_778), .Y(n_777) );
AOI31xp33_ASAP7_75t_L g803 ( .A1(n_673), .A2(n_751), .A3(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g736 ( .A(n_675), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g839 ( .A(n_675), .Y(n_839) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_678), .B(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g778 ( .A(n_678), .B(n_708), .Y(n_778) );
INVx1_ASAP7_75t_L g804 ( .A(n_678), .Y(n_804) );
AND2x2_ASAP7_75t_L g755 ( .A(n_679), .B(n_695), .Y(n_755) );
AND2x2_ASAP7_75t_L g806 ( .A(n_679), .B(n_733), .Y(n_806) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B1(n_686), .B2(n_693), .C1(n_696), .C2(n_700), .Y(n_680) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
OR2x2_ASAP7_75t_L g791 ( .A(n_688), .B(n_690), .Y(n_791) );
OA211x2_ASAP7_75t_L g802 ( .A1(n_688), .A2(n_803), .B(n_807), .C(n_811), .Y(n_802) );
OAI21xp33_ASAP7_75t_L g851 ( .A1(n_689), .A2(n_699), .B(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_694), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_695), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g816 ( .A(n_695), .Y(n_816) );
AND2x2_ASAP7_75t_L g835 ( .A(n_695), .B(n_787), .Y(n_835) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
AND2x2_ASAP7_75t_L g818 ( .A(n_697), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g805 ( .A(n_699), .B(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_702), .B(n_855), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_730), .C(n_746), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_710), .B1(n_720), .B2(n_724), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g801 ( .A(n_707), .Y(n_801) );
INVx1_ASAP7_75t_L g752 ( .A(n_708), .Y(n_752) );
NAND2xp33_ASAP7_75t_SL g710 ( .A(n_711), .B(n_715), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
AND2x4_ASAP7_75t_SL g753 ( .A(n_712), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_SL g797 ( .A(n_712), .Y(n_797) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g716 ( .A(n_713), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g757 ( .A(n_713), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g754 ( .A(n_714), .Y(n_754) );
OAI22xp33_ASAP7_75t_R g847 ( .A1(n_714), .A2(n_741), .B1(n_773), .B2(n_848), .Y(n_847) );
NAND2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g737 ( .A(n_716), .Y(n_737) );
AND2x2_ASAP7_75t_L g845 ( .A(n_716), .B(n_754), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_717), .B(n_719), .Y(n_822) );
AND2x4_ASAP7_75t_L g781 ( .A(n_718), .B(n_782), .Y(n_781) );
OAI32xp33_ASAP7_75t_L g812 ( .A1(n_718), .A2(n_732), .A3(n_813), .B1(n_814), .B2(n_816), .Y(n_812) );
INVx1_ASAP7_75t_L g848 ( .A(n_718), .Y(n_848) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g782 ( .A(n_722), .Y(n_782) );
INVx1_ASAP7_75t_L g815 ( .A(n_722), .Y(n_815) );
OAI22xp33_ASAP7_75t_SL g747 ( .A1(n_723), .A2(n_748), .B1(n_750), .B2(n_752), .Y(n_747) );
INVx2_ASAP7_75t_L g758 ( .A(n_723), .Y(n_758) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
OR2x2_ASAP7_75t_L g762 ( .A(n_726), .B(n_763), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_735), .B1(n_738), .B2(n_742), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_733), .Y(n_826) );
OAI21xp33_ASAP7_75t_L g807 ( .A1(n_735), .A2(n_808), .B(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI221xp5_ASAP7_75t_L g761 ( .A1(n_739), .A2(n_758), .B1(n_762), .B2(n_764), .C(n_767), .Y(n_761) );
OR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
AOI33xp33_ASAP7_75t_L g746 ( .A1(n_740), .A2(n_747), .A3(n_753), .B1(n_755), .B2(n_756), .B3(n_759), .Y(n_746) );
INVx1_ASAP7_75t_L g810 ( .A(n_740), .Y(n_810) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx2_ASAP7_75t_L g789 ( .A(n_743), .Y(n_789) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_745), .A2(n_789), .B(n_790), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_745), .B(n_815), .Y(n_814) );
INVxp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI32xp33_ASAP7_75t_L g834 ( .A1(n_757), .A2(n_835), .A3(n_836), .B1(n_837), .B2(n_884), .Y(n_834) );
AND2x4_ASAP7_75t_SL g793 ( .A(n_758), .B(n_769), .Y(n_793) );
NOR3x1_ASAP7_75t_L g760 ( .A(n_761), .B(n_776), .C(n_783), .Y(n_760) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g827 ( .A(n_765), .B(n_813), .Y(n_827) );
AND2x2_ASAP7_75t_L g770 ( .A(n_766), .B(n_771), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_770), .B(n_772), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_768), .A2(n_847), .B1(n_849), .B2(n_850), .Y(n_846) );
AND2x2_ASAP7_75t_L g796 ( .A(n_771), .B(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_778), .A2(n_793), .B1(n_832), .B2(n_833), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g819 ( .A(n_782), .Y(n_819) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_788), .B1(n_792), .B2(n_794), .C(n_795), .Y(n_783) );
OR2x6_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g808 ( .A(n_789), .Y(n_808) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .Y(n_795) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OR2x6_ASAP7_75t_L g853 ( .A(n_801), .B(n_854), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_817), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_820), .B1(n_822), .B2(n_823), .Y(n_817) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVxp33_ASAP7_75t_L g823 ( .A(n_821), .Y(n_823) );
OR2x2_ASAP7_75t_L g838 ( .A(n_822), .B(n_839), .Y(n_838) );
AOI211x1_ASAP7_75t_SL g824 ( .A1(n_825), .A2(n_827), .B(n_828), .C(n_840), .Y(n_824) );
NAND3xp33_ASAP7_75t_SL g828 ( .A(n_829), .B(n_831), .C(n_834), .Y(n_828) );
INVx1_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
OAI211xp5_ASAP7_75t_SL g840 ( .A1(n_841), .A2(n_844), .B(n_846), .C(n_851), .Y(n_840) );
OR2x2_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_862), .B(n_874), .Y(n_859) );
INVx3_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_869), .B(n_870), .C(n_873), .Y(n_862) );
NAND2xp5_ASAP7_75t_SL g863 ( .A(n_864), .B(n_866), .Y(n_863) );
INVx5_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g870 ( .A(n_867), .B(n_869), .C(n_871), .Y(n_870) );
INVx6_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
BUFx6f_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
BUFx12f_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
endmodule