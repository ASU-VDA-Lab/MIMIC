module fake_jpeg_27002_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_55),
.B1(n_59),
.B2(n_68),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_65),
.B1(n_66),
.B2(n_49),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_53),
.B1(n_50),
.B2(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_83),
.B1(n_89),
.B2(n_66),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_53),
.B1(n_75),
.B2(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_62),
.B1(n_54),
.B2(n_68),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_0),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_103),
.B1(n_86),
.B2(n_83),
.Y(n_104)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_57),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_56),
.B(n_48),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_69),
.B1(n_61),
.B2(n_58),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_63),
.B1(n_51),
.B2(n_65),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_98),
.B1(n_95),
.B2(n_6),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_117),
.B(n_43),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_16),
.B1(n_40),
.B2(n_39),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_15),
.C(n_36),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_2),
.C(n_3),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_14),
.B1(n_34),
.B2(n_33),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_26),
.B(n_32),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_123),
.B(n_127),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_5),
.C(n_7),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_124),
.B1(n_125),
.B2(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_4),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_4),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_9),
.B(n_10),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_115),
.C(n_106),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_137),
.Y(n_148)
);

NOR2x1_ASAP7_75t_R g132 ( 
.A(n_120),
.B(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_140),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_28),
.B(n_27),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_132),
.B1(n_138),
.B2(n_134),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_149),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_142),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_150),
.B(n_146),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_146),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_131),
.B(n_130),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_148),
.B1(n_17),
.B2(n_19),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_148),
.Y(n_160)
);


endmodule