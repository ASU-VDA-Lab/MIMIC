module real_aes_9189_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_0), .B(n_89), .C(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
INVx1_ASAP7_75t_L g526 ( .A(n_1), .Y(n_526) );
INVx1_ASAP7_75t_L g162 ( .A(n_2), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_3), .A2(n_751), .B1(n_754), .B2(n_755), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_3), .Y(n_755) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_4), .A2(n_21), .B1(n_131), .B2(n_132), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_4), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_5), .A2(n_39), .B1(n_187), .B2(n_482), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g206 ( .A1(n_6), .A2(n_178), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_7), .B(n_176), .Y(n_537) );
AND2x6_ASAP7_75t_L g155 ( .A(n_8), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_9), .A2(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_10), .B(n_40), .Y(n_128) );
INVx1_ASAP7_75t_L g212 ( .A(n_11), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_12), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g147 ( .A(n_13), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_14), .B(n_168), .Y(n_490) );
INVx1_ASAP7_75t_L g266 ( .A(n_15), .Y(n_266) );
INVx1_ASAP7_75t_L g520 ( .A(n_16), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_17), .B(n_143), .Y(n_542) );
AO32x2_ASAP7_75t_L g509 ( .A1(n_18), .A2(n_142), .A3(n_176), .B1(n_484), .B2(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_19), .B(n_187), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_20), .B(n_183), .Y(n_254) );
INVxp67_ASAP7_75t_L g131 ( .A(n_21), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_21), .B(n_143), .Y(n_528) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_22), .A2(n_32), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_22), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_23), .A2(n_53), .B1(n_187), .B2(n_482), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_24), .B(n_178), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_25), .A2(n_80), .B1(n_168), .B2(n_187), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_26), .B(n_187), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_27), .B(n_190), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_28), .A2(n_264), .B(n_265), .C(n_267), .Y(n_263) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_29), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_30), .B(n_173), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_31), .B(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_32), .Y(n_455) );
INVx1_ASAP7_75t_L g201 ( .A(n_33), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_34), .B(n_173), .Y(n_507) );
INVx2_ASAP7_75t_L g153 ( .A(n_35), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_36), .B(n_187), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_37), .B(n_173), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_38), .A2(n_155), .B(n_158), .C(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_40), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g199 ( .A(n_41), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_42), .B(n_166), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_43), .B(n_459), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_44), .A2(n_463), .B1(n_746), .B2(n_747), .C1(n_756), .C2(n_758), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_45), .B(n_187), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_46), .A2(n_105), .B1(n_116), .B2(n_763), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_47), .A2(n_90), .B1(n_230), .B2(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_48), .B(n_187), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_49), .B(n_187), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_50), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_51), .B(n_525), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_52), .B(n_178), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_54), .A2(n_64), .B1(n_168), .B2(n_187), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_55), .A2(n_158), .B1(n_168), .B2(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_56), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_57), .B(n_187), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_58), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_59), .B(n_187), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_60), .A2(n_186), .B(n_210), .C(n_211), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_61), .Y(n_257) );
INVx1_ASAP7_75t_L g208 ( .A(n_62), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_63), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_63), .Y(n_748) );
INVx1_ASAP7_75t_L g156 ( .A(n_65), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_66), .B(n_187), .Y(n_527) );
INVx1_ASAP7_75t_L g146 ( .A(n_67), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_68), .Y(n_121) );
AO32x2_ASAP7_75t_L g479 ( .A1(n_69), .A2(n_176), .A3(n_235), .B1(n_480), .B2(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g559 ( .A(n_70), .Y(n_559) );
INVx1_ASAP7_75t_L g502 ( .A(n_71), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_72), .A2(n_79), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_72), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_SL g182 ( .A1(n_73), .A2(n_183), .B(n_184), .C(n_186), .Y(n_182) );
INVxp67_ASAP7_75t_L g185 ( .A(n_74), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_75), .B(n_168), .Y(n_503) );
INVx1_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_77), .Y(n_204) );
INVx1_ASAP7_75t_L g250 ( .A(n_78), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_79), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_81), .A2(n_155), .B(n_158), .C(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_82), .B(n_482), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_83), .B(n_168), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_84), .B(n_163), .Y(n_226) );
INVx2_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_86), .B(n_183), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_87), .B(n_168), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_88), .A2(n_155), .B(n_158), .C(n_161), .Y(n_157) );
OR2x2_ASAP7_75t_L g124 ( .A(n_89), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g466 ( .A(n_89), .B(n_126), .Y(n_466) );
INVx2_ASAP7_75t_L g470 ( .A(n_89), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_91), .A2(n_103), .B1(n_168), .B2(n_169), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_92), .B(n_173), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_93), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_94), .A2(n_155), .B(n_158), .C(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_95), .Y(n_245) );
INVx1_ASAP7_75t_L g181 ( .A(n_96), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_97), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_98), .B(n_163), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_99), .B(n_168), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_100), .B(n_176), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_101), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_102), .A2(n_178), .B(n_179), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_108), .Y(n_764) );
CKINVDCx9p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_461), .Y(n_116) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g762 ( .A(n_120), .Y(n_762) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_129), .B(n_458), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_124), .Y(n_460) );
NOR2x2_ASAP7_75t_L g760 ( .A(n_125), .B(n_470), .Y(n_760) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g469 ( .A(n_126), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_133), .B1(n_134), .B2(n_457), .Y(n_129) );
INVx1_ASAP7_75t_L g457 ( .A(n_130), .Y(n_457) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_452), .B1(n_453), .B2(n_456), .Y(n_134) );
INVx2_ASAP7_75t_L g456 ( .A(n_135), .Y(n_456) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_135), .A2(n_464), .B1(n_472), .B2(n_757), .Y(n_756) );
OR4x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_341), .C(n_401), .D(n_428), .Y(n_135) );
NAND4xp25_ASAP7_75t_SL g136 ( .A(n_137), .B(n_289), .C(n_320), .D(n_337), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_214), .B(n_216), .C(n_269), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_192), .Y(n_138) );
INVx1_ASAP7_75t_L g331 ( .A(n_139), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_139), .A2(n_372), .B1(n_420), .B2(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_174), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_140), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g282 ( .A(n_140), .B(n_194), .Y(n_282) );
AND2x2_ASAP7_75t_L g324 ( .A(n_140), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_140), .B(n_215), .Y(n_336) );
INVx1_ASAP7_75t_L g376 ( .A(n_140), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_140), .B(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g304 ( .A(n_141), .B(n_194), .Y(n_304) );
INVx3_ASAP7_75t_L g308 ( .A(n_141), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_141), .B(n_366), .Y(n_365) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_148), .B(n_170), .Y(n_141) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_142), .A2(n_195), .B(n_203), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_142), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g231 ( .A(n_142), .Y(n_231) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_144), .B(n_145), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_157), .Y(n_148) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_150), .A2(n_188), .B1(n_196), .B2(n_202), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_150), .A2(n_250), .B(n_251), .Y(n_249) );
NAND2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
AND2x4_ASAP7_75t_L g178 ( .A(n_151), .B(n_155), .Y(n_178) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
INVx1_ASAP7_75t_L g525 ( .A(n_152), .Y(n_525) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
INVx1_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
INVx1_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
INVx3_ASAP7_75t_L g164 ( .A(n_154), .Y(n_164) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_154), .Y(n_166) );
INVx1_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_154), .Y(n_198) );
INVx4_ASAP7_75t_SL g188 ( .A(n_155), .Y(n_188) );
BUFx3_ASAP7_75t_L g484 ( .A(n_155), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_155), .A2(n_488), .B(n_492), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_155), .A2(n_501), .B(n_504), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_155), .A2(n_519), .B(n_523), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_155), .A2(n_531), .B(n_534), .Y(n_530) );
INVx5_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
AND2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
BUFx3_ASAP7_75t_L g230 ( .A(n_159), .Y(n_230) );
INVx1_ASAP7_75t_L g482 ( .A(n_159), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_165), .C(n_167), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_SL g501 ( .A1(n_163), .A2(n_186), .B(n_502), .C(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g512 ( .A(n_163), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_163), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_163), .A2(n_556), .B(n_557), .Y(n_555) );
INVx5_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_164), .B(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_164), .B(n_212), .Y(n_211) );
OAI22xp5_ASAP7_75t_SL g480 ( .A1(n_164), .A2(n_166), .B1(n_481), .B2(n_483), .Y(n_480) );
INVx2_ASAP7_75t_L g210 ( .A(n_166), .Y(n_210) );
INVx4_ASAP7_75t_L g241 ( .A(n_166), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_166), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_166), .A2(n_512), .B1(n_545), .B2(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_167), .A2(n_520), .B(n_521), .C(n_522), .Y(n_519) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_172), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_172), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g235 ( .A(n_173), .Y(n_235) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_173), .A2(n_259), .B(n_268), .Y(n_258) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_173), .A2(n_487), .B(n_495), .Y(n_486) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_173), .A2(n_500), .B(n_507), .Y(n_499) );
AND2x2_ASAP7_75t_L g395 ( .A(n_174), .B(n_205), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_174), .B(n_308), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_174), .B(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g215 ( .A(n_175), .B(n_194), .Y(n_215) );
INVx1_ASAP7_75t_L g277 ( .A(n_175), .Y(n_277) );
BUFx2_ASAP7_75t_L g281 ( .A(n_175), .Y(n_281) );
AND2x2_ASAP7_75t_L g325 ( .A(n_175), .B(n_193), .Y(n_325) );
OR2x2_ASAP7_75t_L g364 ( .A(n_175), .B(n_193), .Y(n_364) );
AND2x2_ASAP7_75t_L g389 ( .A(n_175), .B(n_205), .Y(n_389) );
AND2x2_ASAP7_75t_L g448 ( .A(n_175), .B(n_278), .Y(n_448) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_189), .Y(n_175) );
INVx4_ASAP7_75t_L g191 ( .A(n_176), .Y(n_191) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_176), .A2(n_530), .B(n_537), .Y(n_529) );
BUFx2_ASAP7_75t_L g260 ( .A(n_178), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_188), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_180), .A2(n_188), .B(n_208), .C(n_209), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_180), .A2(n_188), .B(n_262), .C(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g491 ( .A(n_183), .Y(n_491) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_187), .Y(n_242) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_190), .A2(n_206), .B(n_213), .Y(n_205) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_191), .B(n_233), .Y(n_232) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_191), .B(n_484), .C(n_544), .Y(n_543) );
AO21x1_ASAP7_75t_L g590 ( .A1(n_191), .A2(n_544), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g423 ( .A(n_192), .Y(n_423) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_205), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_193), .B(n_205), .Y(n_309) );
AND2x2_ASAP7_75t_L g319 ( .A(n_193), .B(n_308), .Y(n_319) );
BUFx2_ASAP7_75t_L g330 ( .A(n_193), .Y(n_330) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g352 ( .A(n_194), .B(n_205), .Y(n_352) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_194), .Y(n_407) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_198), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g200 ( .A(n_198), .Y(n_200) );
INVx4_ASAP7_75t_L g264 ( .A(n_198), .Y(n_264) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_205), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_SL g278 ( .A(n_205), .Y(n_278) );
BUFx2_ASAP7_75t_L g303 ( .A(n_205), .Y(n_303) );
INVx2_ASAP7_75t_L g322 ( .A(n_205), .Y(n_322) );
AND2x2_ASAP7_75t_L g384 ( .A(n_205), .B(n_308), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_210), .A2(n_493), .B(n_494), .Y(n_492) );
O2A1O1Ixp5_ASAP7_75t_L g558 ( .A1(n_210), .A2(n_524), .B(n_559), .C(n_560), .Y(n_558) );
AOI321xp33_ASAP7_75t_L g403 ( .A1(n_214), .A2(n_404), .A3(n_405), .B1(n_406), .B2(n_408), .C(n_409), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_215), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_215), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g397 ( .A(n_215), .B(n_376), .Y(n_397) );
AND2x2_ASAP7_75t_L g430 ( .A(n_215), .B(n_322), .Y(n_430) );
INVx1_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_246), .Y(n_217) );
OR2x2_ASAP7_75t_L g332 ( .A(n_218), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_234), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g284 ( .A(n_221), .Y(n_284) );
AND2x2_ASAP7_75t_L g294 ( .A(n_221), .B(n_248), .Y(n_294) );
AND2x2_ASAP7_75t_L g299 ( .A(n_221), .B(n_274), .Y(n_299) );
INVx1_ASAP7_75t_L g316 ( .A(n_221), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_221), .B(n_297), .Y(n_335) );
AND2x2_ASAP7_75t_L g340 ( .A(n_221), .B(n_273), .Y(n_340) );
OR2x2_ASAP7_75t_L g372 ( .A(n_221), .B(n_361), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_221), .B(n_285), .Y(n_411) );
AND2x2_ASAP7_75t_L g445 ( .A(n_221), .B(n_271), .Y(n_445) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_232), .Y(n_221) );
AOI21xp5_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_224), .B(n_231), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_228), .A2(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g267 ( .A(n_230), .Y(n_267) );
INVx1_ASAP7_75t_L g255 ( .A(n_231), .Y(n_255) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_231), .A2(n_518), .B(n_528), .Y(n_517) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_231), .A2(n_554), .B(n_561), .Y(n_553) );
INVx1_ASAP7_75t_L g272 ( .A(n_234), .Y(n_272) );
INVx2_ASAP7_75t_L g287 ( .A(n_234), .Y(n_287) );
AND2x2_ASAP7_75t_L g327 ( .A(n_234), .B(n_298), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_234), .B(n_274), .Y(n_349) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_242), .Y(n_238) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g433 ( .A(n_247), .B(n_284), .Y(n_433) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_258), .Y(n_247) );
INVx2_ASAP7_75t_L g274 ( .A(n_248), .Y(n_274) );
AND2x2_ASAP7_75t_L g427 ( .A(n_248), .B(n_287), .Y(n_427) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_255), .B(n_256), .Y(n_248) );
AND2x2_ASAP7_75t_L g273 ( .A(n_258), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g288 ( .A(n_258), .Y(n_288) );
INVx1_ASAP7_75t_L g298 ( .A(n_258), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_264), .B(n_266), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_264), .A2(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g522 ( .A(n_264), .Y(n_522) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_275), .B1(n_279), .B2(n_283), .Y(n_269) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_270), .A2(n_388), .B1(n_425), .B2(n_426), .Y(n_424) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g339 ( .A(n_272), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_273), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g334 ( .A(n_274), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_274), .B(n_287), .Y(n_361) );
INVx1_ASAP7_75t_L g377 ( .A(n_274), .Y(n_377) );
AND2x2_ASAP7_75t_L g318 ( .A(n_276), .B(n_319), .Y(n_318) );
INVx3_ASAP7_75t_SL g357 ( .A(n_276), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_276), .B(n_282), .Y(n_434) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g443 ( .A(n_279), .Y(n_443) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_280), .B(n_376), .Y(n_418) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx3_ASAP7_75t_SL g323 ( .A(n_282), .Y(n_323) );
NAND2x1_ASAP7_75t_SL g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g344 ( .A(n_284), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g351 ( .A(n_284), .B(n_288), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_284), .B(n_297), .Y(n_356) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_284), .Y(n_405) );
OAI311xp33_ASAP7_75t_L g428 ( .A1(n_285), .A2(n_429), .A3(n_431), .B1(n_432), .C1(n_442), .Y(n_428) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g441 ( .A(n_286), .B(n_314), .Y(n_441) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g297 ( .A(n_287), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g345 ( .A(n_287), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g400 ( .A(n_287), .Y(n_400) );
INVx1_ASAP7_75t_L g293 ( .A(n_288), .Y(n_293) );
INVx1_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_288), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g346 ( .A(n_288), .Y(n_346) );
AOI221xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_292), .B1(n_300), .B2(n_305), .C(n_310), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx4_ASAP7_75t_L g314 ( .A(n_294), .Y(n_314) );
AND2x2_ASAP7_75t_L g408 ( .A(n_294), .B(n_327), .Y(n_408) );
AND2x2_ASAP7_75t_L g415 ( .A(n_294), .B(n_297), .Y(n_415) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_297), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g326 ( .A(n_299), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_302), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g451 ( .A(n_304), .B(n_395), .Y(n_451) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g436 ( .A(n_308), .B(n_364), .Y(n_436) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_309), .A2(n_402), .B(n_403), .C(n_416), .Y(n_401) );
AOI21xp33_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_315), .B(n_317), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g380 ( .A(n_314), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_315), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_413), .Y(n_409) );
AND2x2_ASAP7_75t_L g386 ( .A(n_316), .B(n_327), .Y(n_386) );
AND2x2_ASAP7_75t_L g439 ( .A(n_316), .B(n_334), .Y(n_439) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_319), .B(n_357), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .B(n_326), .C(n_328), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g367 ( .A(n_322), .B(n_325), .Y(n_367) );
OR2x2_ASAP7_75t_L g410 ( .A(n_322), .B(n_364), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_323), .B(n_389), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_323), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g354 ( .A(n_324), .Y(n_354) );
INVx1_ASAP7_75t_L g420 ( .A(n_327), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B1(n_335), .B2(n_336), .Y(n_328) );
INVx1_ASAP7_75t_L g343 ( .A(n_329), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_330), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g406 ( .A(n_331), .B(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g392 ( .A(n_333), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_334), .B(n_420), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_335), .A2(n_394), .B1(n_396), .B2(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g402 ( .A(n_338), .Y(n_402) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x2_ASAP7_75t_L g444 ( .A(n_339), .B(n_439), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_374), .B1(n_377), .B2(n_378), .C1(n_381), .C2(n_382), .Y(n_373) );
NAND4xp25_ASAP7_75t_SL g341 ( .A(n_342), .B(n_362), .C(n_373), .D(n_385), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_347), .B2(n_352), .C(n_353), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_345), .B(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_347), .A2(n_417), .B1(n_419), .B2(n_421), .C(n_424), .Y(n_416) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g359 ( .A(n_351), .B(n_360), .Y(n_359) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_352), .A2(n_414), .B(n_415), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_357), .B2(n_358), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_368), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_376), .B(n_395), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_376), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_380), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g412 ( .A(n_384), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_390), .B2(n_392), .C(n_393), .Y(n_385) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_395), .A2(n_433), .B1(n_434), .B2(n_435), .C1(n_437), .C2(n_440), .Y(n_432) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_399), .B(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVxp33_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_445), .B2(n_446), .C(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_456), .A2(n_464), .B1(n_467), .B2(n_471), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_458), .B(n_462), .C(n_761), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g757 ( .A(n_468), .Y(n_757) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND3x1_ASAP7_75t_L g473 ( .A(n_474), .B(n_666), .C(n_714), .Y(n_473) );
NOR4xp25_ASAP7_75t_L g474 ( .A(n_475), .B(n_594), .C(n_639), .D(n_653), .Y(n_474) );
OAI311xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_514), .A3(n_538), .B1(n_547), .C1(n_562), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_485), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_477), .A2(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g655 ( .A(n_477), .B(n_582), .Y(n_655) );
AND2x2_ASAP7_75t_L g712 ( .A(n_477), .B(n_598), .Y(n_712) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g605 ( .A(n_478), .B(n_508), .Y(n_605) );
AND2x2_ASAP7_75t_L g662 ( .A(n_478), .B(n_610), .Y(n_662) );
INVx1_ASAP7_75t_L g703 ( .A(n_478), .Y(n_703) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_479), .Y(n_571) );
AND2x2_ASAP7_75t_L g612 ( .A(n_479), .B(n_508), .Y(n_612) );
AND2x2_ASAP7_75t_L g616 ( .A(n_479), .B(n_509), .Y(n_616) );
INVx1_ASAP7_75t_L g628 ( .A(n_479), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_484), .A2(n_555), .B(n_558), .Y(n_554) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
AND2x2_ASAP7_75t_L g549 ( .A(n_486), .B(n_508), .Y(n_549) );
INVx2_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
AND2x2_ASAP7_75t_L g598 ( .A(n_486), .B(n_509), .Y(n_598) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_486), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_486), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g618 ( .A(n_486), .B(n_581), .Y(n_618) );
INVx1_ASAP7_75t_L g630 ( .A(n_486), .Y(n_630) );
INVx1_ASAP7_75t_L g671 ( .A(n_486), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_486), .B(n_571), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_491), .Y(n_488) );
NOR2xp67_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g548 ( .A(n_498), .B(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_498), .Y(n_576) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_498), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g633 ( .A(n_498), .B(n_508), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_498), .B(n_628), .Y(n_691) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g581 ( .A(n_499), .Y(n_581) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_499), .Y(n_597) );
OR2x2_ASAP7_75t_L g670 ( .A(n_499), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g577 ( .A(n_509), .Y(n_577) );
AND2x2_ASAP7_75t_L g582 ( .A(n_509), .B(n_583), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_512), .A2(n_524), .B(n_526), .C(n_527), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_512), .A2(n_535), .B(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_514), .B(n_565), .Y(n_728) );
INVx1_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g698 ( .A(n_515), .B(n_540), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_529), .Y(n_515) );
AND2x2_ASAP7_75t_L g574 ( .A(n_516), .B(n_565), .Y(n_574) );
INVx2_ASAP7_75t_L g586 ( .A(n_516), .Y(n_586) );
AND2x2_ASAP7_75t_L g620 ( .A(n_516), .B(n_568), .Y(n_620) );
AND2x2_ASAP7_75t_L g687 ( .A(n_516), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_517), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g567 ( .A(n_517), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g607 ( .A(n_517), .B(n_529), .Y(n_607) );
AND2x2_ASAP7_75t_L g624 ( .A(n_517), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g550 ( .A(n_529), .B(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g568 ( .A(n_529), .Y(n_568) );
AND2x2_ASAP7_75t_L g573 ( .A(n_529), .B(n_553), .Y(n_573) );
AND2x2_ASAP7_75t_L g646 ( .A(n_529), .B(n_625), .Y(n_646) );
AND2x2_ASAP7_75t_L g711 ( .A(n_529), .B(n_701), .Y(n_711) );
OAI311xp33_ASAP7_75t_L g594 ( .A1(n_538), .A2(n_595), .A3(n_599), .B1(n_601), .C1(n_621), .Y(n_594) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g606 ( .A(n_539), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g665 ( .A(n_539), .B(n_573), .Y(n_665) );
AND2x2_ASAP7_75t_L g739 ( .A(n_539), .B(n_620), .Y(n_739) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_540), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g674 ( .A(n_540), .Y(n_674) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx3_ASAP7_75t_L g565 ( .A(n_541), .Y(n_565) );
NOR2x1_ASAP7_75t_L g637 ( .A(n_541), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g694 ( .A(n_541), .B(n_568), .Y(n_694) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g591 ( .A(n_542), .Y(n_591) );
AND2x2_ASAP7_75t_L g569 ( .A(n_549), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g622 ( .A(n_549), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g702 ( .A(n_549), .B(n_703), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_550), .A2(n_582), .B1(n_602), .B2(n_606), .C(n_608), .Y(n_601) );
INVx1_ASAP7_75t_L g726 ( .A(n_551), .Y(n_726) );
OR2x2_ASAP7_75t_L g692 ( .A(n_552), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g587 ( .A(n_553), .B(n_568), .Y(n_587) );
OR2x2_ASAP7_75t_L g589 ( .A(n_553), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g614 ( .A(n_553), .Y(n_614) );
INVx2_ASAP7_75t_L g625 ( .A(n_553), .Y(n_625) );
AND2x2_ASAP7_75t_L g652 ( .A(n_553), .B(n_590), .Y(n_652) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_553), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_569), .B1(n_572), .B2(n_575), .C(n_578), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g663 ( .A(n_565), .B(n_573), .Y(n_663) );
AND2x2_ASAP7_75t_L g713 ( .A(n_565), .B(n_567), .Y(n_713) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g600 ( .A(n_567), .B(n_571), .Y(n_600) );
AND2x2_ASAP7_75t_L g679 ( .A(n_567), .B(n_652), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_568), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g638 ( .A(n_568), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g648 ( .A1(n_569), .A2(n_649), .B(n_651), .Y(n_648) );
OR2x2_ASAP7_75t_L g592 ( .A(n_570), .B(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g658 ( .A(n_570), .B(n_618), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_570), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g635 ( .A(n_571), .B(n_604), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_571), .B(n_718), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_572), .B(n_598), .Y(n_708) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g631 ( .A(n_573), .B(n_586), .Y(n_631) );
INVx1_ASAP7_75t_L g647 ( .A(n_574), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_584), .B1(n_588), .B2(n_592), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g610 ( .A(n_581), .Y(n_610) );
INVx1_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
INVx1_ASAP7_75t_L g593 ( .A(n_582), .Y(n_593) );
AND2x2_ASAP7_75t_L g664 ( .A(n_582), .B(n_610), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_582), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
OR2x2_ASAP7_75t_L g588 ( .A(n_585), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_585), .B(n_701), .Y(n_700) );
NOR2xp67_ASAP7_75t_L g732 ( .A(n_585), .B(n_733), .Y(n_732) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g735 ( .A(n_587), .B(n_687), .Y(n_735) );
INVx1_ASAP7_75t_SL g701 ( .A(n_589), .Y(n_701) );
AND2x2_ASAP7_75t_L g641 ( .A(n_590), .B(n_625), .Y(n_641) );
INVx1_ASAP7_75t_L g688 ( .A(n_590), .Y(n_688) );
OAI222xp33_ASAP7_75t_L g729 ( .A1(n_595), .A2(n_685), .B1(n_730), .B2(n_731), .C1(n_734), .C2(n_736), .Y(n_729) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g650 ( .A(n_597), .Y(n_650) );
AND2x2_ASAP7_75t_L g661 ( .A(n_598), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_598), .B(n_703), .Y(n_730) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_600), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g705 ( .A(n_602), .Y(n_705) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g643 ( .A(n_605), .Y(n_643) );
AND2x2_ASAP7_75t_L g722 ( .A(n_605), .B(n_683), .Y(n_722) );
AND2x2_ASAP7_75t_L g745 ( .A(n_605), .B(n_629), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_607), .B(n_641), .Y(n_640) );
OAI32xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .A3(n_613), .B1(n_615), .B2(n_619), .Y(n_608) );
BUFx2_ASAP7_75t_L g683 ( .A(n_610), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_611), .B(n_629), .Y(n_710) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g649 ( .A(n_612), .B(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g717 ( .A(n_612), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g706 ( .A(n_613), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g677 ( .A(n_616), .B(n_650), .Y(n_677) );
INVx2_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g639 ( .A1(n_618), .A2(n_640), .B1(n_642), .B2(n_644), .C(n_648), .Y(n_639) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g651 ( .A(n_620), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g657 ( .A(n_620), .B(n_641), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_626), .B2(n_631), .C(n_632), .Y(n_621) );
INVx1_ASAP7_75t_L g740 ( .A(n_622), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_623), .B(n_717), .Y(n_716) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_624), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_629), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g695 ( .A(n_629), .Y(n_695) );
BUFx3_ASAP7_75t_L g718 ( .A(n_630), .Y(n_718) );
INVx1_ASAP7_75t_SL g659 ( .A(n_631), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_631), .B(n_673), .Y(n_672) );
AOI21xp33_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_634), .B(n_636), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_633), .A2(n_734), .B1(n_738), .B2(n_740), .C(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g680 ( .A(n_638), .B(n_641), .Y(n_680) );
INVx1_ASAP7_75t_L g744 ( .A(n_638), .Y(n_744) );
INVx2_ASAP7_75t_L g733 ( .A(n_641), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_641), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g686 ( .A(n_646), .B(n_687), .Y(n_686) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B1(n_658), .B2(n_659), .C(n_660), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_662), .A2(n_724), .B1(n_725), .B2(n_727), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_665), .A2(n_742), .B(n_745), .Y(n_741) );
NOR4xp25_ASAP7_75t_SL g666 ( .A(n_667), .B(n_675), .C(n_684), .D(n_704), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_672), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B1(n_681), .B2(n_682), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g720 ( .A(n_680), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B1(n_692), .B2(n_695), .C(n_696), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g707 ( .A(n_687), .Y(n_707) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI21xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_699), .B(n_702), .Y(n_696) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B(n_708), .C(n_709), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_709) );
CKINVDCx14_ASAP7_75t_R g719 ( .A(n_713), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_729), .C(n_737), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .B1(n_720), .B2(n_721), .C(n_723), .Y(n_715) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx16_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
CKINVDCx16_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g754 ( .A(n_751), .Y(n_754) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
endmodule