module fake_jpeg_3698_n_6 (n_0, n_1, n_6);

input n_0;
input n_1;

output n_6;

wire n_3;
wire n_2;
wire n_4;
wire n_5;

INVx1_ASAP7_75t_SL g2 ( 
.A(n_0),
.Y(n_2)
);

INVx8_ASAP7_75t_L g3 ( 
.A(n_0),
.Y(n_3)
);

A2O1A1Ixp33_ASAP7_75t_SL g4 ( 
.A1(n_2),
.A2(n_1),
.B(n_3),
.C(n_0),
.Y(n_4)
);

MAJIxp5_ASAP7_75t_L g5 ( 
.A(n_4),
.B(n_2),
.C(n_1),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);


endmodule