module fake_jpeg_31409_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_65),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_51),
.Y(n_85)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_1),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_66),
.B1(n_65),
.B2(n_49),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_90),
.B1(n_68),
.B2(n_42),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_64),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_55),
.B(n_63),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_68),
.C(n_41),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_49),
.B1(n_69),
.B2(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_70),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_79),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_69),
.B1(n_52),
.B2(n_58),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_106),
.B1(n_111),
.B2(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_107),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_67),
.B1(n_61),
.B2(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_112),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_68),
.B1(n_17),
.B2(n_18),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_9),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_37),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_2),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_86),
.C(n_38),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_125),
.C(n_134),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_29),
.B1(n_34),
.B2(n_33),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_128),
.B1(n_9),
.B2(n_10),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_124),
.Y(n_136)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_4),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_32),
.C(n_28),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_7),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_8),
.Y(n_132)
);

NOR4xp25_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_133),
.C(n_134),
.D(n_12),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_8),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_26),
.C(n_22),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_10),
.B(n_11),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_11),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_127),
.B(n_113),
.C(n_115),
.D(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_140),
.C(n_136),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_148),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_139),
.C(n_156),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_141),
.C(n_116),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_158),
.B(n_144),
.C(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_155),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_152),
.B(n_157),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_138),
.A3(n_154),
.B1(n_147),
.B2(n_142),
.C1(n_165),
.C2(n_128),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_135),
.B(n_121),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_13),
.Y(n_171)
);


endmodule