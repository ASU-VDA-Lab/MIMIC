module fake_jpeg_3083_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_0),
.B(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_54),
.Y(n_108)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_7),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g116 ( 
.A(n_55),
.Y(n_116)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx4f_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_11),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_24),
.B(n_5),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_74),
.Y(n_126)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_19),
.B(n_12),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_19),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_88),
.Y(n_130)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_93),
.Y(n_132)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_2),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_52),
.A2(n_31),
.B1(n_21),
.B2(n_44),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_111),
.A2(n_115),
.B1(n_15),
.B2(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_78),
.B1(n_84),
.B2(n_80),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_135),
.B1(n_142),
.B2(n_31),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_41),
.B1(n_45),
.B2(n_44),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_36),
.B1(n_33),
.B2(n_42),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_61),
.B(n_40),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_40),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_145),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_58),
.A2(n_45),
.B1(n_41),
.B2(n_42),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_57),
.B(n_36),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_16),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_148),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_55),
.B(n_2),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_149),
.B(n_162),
.Y(n_211)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_104),
.A2(n_62),
.B1(n_96),
.B2(n_59),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_163),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_21),
.B1(n_90),
.B2(n_89),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_182),
.B1(n_156),
.B2(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_63),
.B1(n_85),
.B2(n_35),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_160),
.A2(n_169),
.B1(n_187),
.B2(n_99),
.Y(n_212)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_71),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_0),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_178),
.Y(n_197)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_71),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_167),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_53),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_116),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_91),
.B1(n_88),
.B2(n_53),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_4),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_98),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_173),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_176),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_0),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_145),
.C(n_97),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_4),
.Y(n_176)
);

BUFx6f_ASAP7_75t_SL g177 ( 
.A(n_116),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_4),
.Y(n_178)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_185),
.C(n_186),
.Y(n_199)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_207)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

AOI22x1_ASAP7_75t_L g182 ( 
.A1(n_123),
.A2(n_29),
.B1(n_46),
.B2(n_13),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_15),
.B(n_46),
.C(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_107),
.B1(n_113),
.B2(n_127),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_198),
.B1(n_210),
.B2(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_194),
.C(n_213),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_153),
.A2(n_132),
.B(n_105),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_201),
.B(n_122),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_132),
.C(n_144),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_150),
.A2(n_100),
.B1(n_144),
.B2(n_124),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_120),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_134),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_171),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_206),
.B1(n_198),
.B2(n_189),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_152),
.B1(n_150),
.B2(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_109),
.C(n_133),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_182),
.B1(n_156),
.B2(n_183),
.Y(n_216)
);

AO22x1_ASAP7_75t_SL g245 ( 
.A1(n_216),
.A2(n_206),
.B1(n_210),
.B2(n_194),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_164),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_175),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_223),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_165),
.B(n_172),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_229),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_197),
.B(n_181),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_161),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_233),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_180),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_235),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_191),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_151),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_208),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_206),
.B1(n_201),
.B2(n_205),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_226),
.B1(n_225),
.B2(n_216),
.C(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_199),
.B1(n_204),
.B2(n_200),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_213),
.B1(n_195),
.B2(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_255),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_232),
.B(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_192),
.C(n_195),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_254),
.C(n_219),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_204),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_258),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_257),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_217),
.A3(n_230),
.B1(n_222),
.B2(n_236),
.C1(n_237),
.C2(n_229),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_242),
.A3(n_244),
.B1(n_241),
.B2(n_245),
.C1(n_258),
.C2(n_257),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_266),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_273),
.B1(n_274),
.B2(n_253),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_243),
.B(n_220),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_270),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_226),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_218),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_249),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_245),
.A2(n_216),
.B1(n_227),
.B2(n_224),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_240),
.B1(n_246),
.B2(n_248),
.Y(n_284)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_231),
.B(n_216),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_216),
.B(n_202),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_202),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_275),
.A2(n_250),
.B1(n_245),
.B2(n_256),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_271),
.B1(n_284),
.B2(n_279),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_253),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_284),
.B1(n_286),
.B2(n_289),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_259),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_264),
.B1(n_262),
.B2(n_242),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_267),
.C(n_266),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_299),
.C(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_298),
.Y(n_307)
);

AND3x1_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_262),
.C(n_268),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_277),
.B(n_196),
.C(n_214),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_295),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_296),
.A2(n_134),
.B1(n_98),
.B2(n_143),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_252),
.B(n_208),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_276),
.B1(n_281),
.B2(n_280),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_196),
.B(n_179),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_214),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_297),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_306),
.B1(n_296),
.B2(n_297),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_290),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_184),
.B1(n_177),
.B2(n_109),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_298),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_302),
.C(n_293),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_307),
.B(n_301),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_313),
.B(n_299),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_319),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_311),
.A2(n_306),
.B1(n_292),
.B2(n_304),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_310),
.Y(n_321)
);

AOI21x1_ASAP7_75t_SL g324 ( 
.A1(n_321),
.A2(n_322),
.B(n_316),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_316),
.C(n_308),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_324),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_143),
.Y(n_327)
);


endmodule