module fake_jpeg_8086_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_8),
.C(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_52),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_20),
.B1(n_16),
.B2(n_32),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_53),
.B1(n_16),
.B2(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_51),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_16),
.B1(n_20),
.B2(n_24),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_24),
.B1(n_25),
.B2(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_20),
.B1(n_33),
.B2(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_52),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_66),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_25),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_17),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_24),
.B(n_23),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_89),
.B(n_18),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_79),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_53),
.B1(n_30),
.B2(n_26),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_29),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_21),
.B1(n_62),
.B2(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_101),
.A2(n_69),
.B1(n_31),
.B2(n_22),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_66),
.B1(n_88),
.B2(n_86),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_110),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_80),
.B1(n_65),
.B2(n_70),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_46),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.C(n_83),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_46),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_128),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_83),
.A3(n_71),
.B1(n_79),
.B2(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_130),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_128),
.CI(n_132),
.CON(n_171),
.SN(n_171)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_129),
.B1(n_109),
.B2(n_115),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_90),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_138),
.C(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_146),
.Y(n_162)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_97),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_56),
.B1(n_84),
.B2(n_69),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_137),
.A2(n_94),
.B1(n_116),
.B2(n_117),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_57),
.C(n_64),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_31),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_147),
.B(n_94),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_73),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_107),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_151),
.C(n_156),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_161),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_98),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_169),
.B1(n_177),
.B2(n_77),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_113),
.C(n_92),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_158),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_98),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_163),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_92),
.C(n_97),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_96),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_109),
.B1(n_112),
.B2(n_99),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_99),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_27),
.B(n_33),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_175),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_13),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_111),
.B1(n_33),
.B2(n_91),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_143),
.B1(n_123),
.B2(n_144),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_143),
.B1(n_144),
.B2(n_133),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_187),
.B1(n_189),
.B2(n_177),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_125),
.B1(n_77),
.B2(n_68),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_149),
.A2(n_125),
.B1(n_77),
.B2(n_68),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_173),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_30),
.B(n_28),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_157),
.B(n_10),
.C(n_15),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_206),
.C(n_156),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_159),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_28),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_10),
.C(n_15),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_171),
.C(n_150),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_SL g244 ( 
.A(n_207),
.B(n_209),
.C(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_201),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_167),
.B1(n_161),
.B2(n_170),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_163),
.B1(n_160),
.B2(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_153),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_214),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_150),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_193),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_148),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_220),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_151),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_171),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_198),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_200),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_229),
.C(n_204),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_177),
.B1(n_174),
.B2(n_178),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_178),
.B1(n_28),
.B2(n_26),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_22),
.B1(n_26),
.B2(n_2),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_27),
.C(n_26),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_185),
.B1(n_199),
.B2(n_180),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_189),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_210),
.B(n_229),
.Y(n_256)
);

FAx1_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_194),
.CI(n_190),
.CON(n_233),
.SN(n_233)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_218),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_182),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_241),
.B(n_15),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_248),
.C(n_251),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_243),
.A2(n_247),
.B1(n_227),
.B2(n_221),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_223),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_199),
.B1(n_9),
.B2(n_11),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_27),
.C(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_8),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_27),
.C(n_3),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_233),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_246),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_256),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_233),
.B(n_245),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_261),
.C(n_263),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_228),
.B1(n_207),
.B2(n_213),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_238),
.B1(n_243),
.B2(n_235),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_217),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_244),
.A2(n_224),
.B1(n_9),
.B2(n_12),
.Y(n_262)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_27),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_0),
.C(n_3),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_248),
.C(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_257),
.Y(n_268)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_14),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_263),
.B(n_3),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_276),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_0),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_261),
.C(n_234),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_265),
.C(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_285),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_290),
.C(n_270),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_291),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_278),
.A2(n_262),
.B1(n_267),
.B2(n_266),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_13),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_3),
.C(n_4),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_277),
.B(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_293),
.B(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_297),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_285),
.B(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_279),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_300),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_272),
.C(n_269),
.Y(n_300)
);

OA21x2_ASAP7_75t_SL g301 ( 
.A1(n_299),
.A2(n_289),
.B(n_286),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_281),
.B(n_269),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_292),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_309),
.B(n_304),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_306),
.B(n_308),
.C(n_302),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_4),
.C(n_6),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_4),
.C(n_6),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_7),
.Y(n_314)
);


endmodule