module real_jpeg_18091_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_288;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_197;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_195;
wire n_110;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_0),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_0),
.B(n_135),
.Y(n_134)
);

AND2x4_ASAP7_75t_SL g180 ( 
.A(n_0),
.B(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_2),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_2),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_2),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_2),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_3),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_4),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_4),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_5),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_5),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_7),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_7),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_7),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_7),
.B(n_114),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_7),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_7),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_8),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_8),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_8),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_8),
.B(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_8),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_8),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_8),
.B(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_9),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_10),
.A2(n_14),
.B1(n_60),
.B2(n_63),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_11),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_115),
.Y(n_152)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_13),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g265 ( 
.A(n_13),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_14),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_14),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_14),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_14),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_15),
.Y(n_147)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_188),
.B1(n_295),
.B2(n_296),
.Y(n_17)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_18),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_186),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_141),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_20),
.B(n_141),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_122),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_21),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_22),
.B(n_44),
.C(n_66),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.C(n_38),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_23),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_24),
.B(n_28),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_24),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_24),
.A2(n_239),
.B1(n_240),
.B2(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_27),
.Y(n_206)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_31),
.Y(n_242)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_33),
.Y(n_282)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_41),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_66),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_53),
.B(n_59),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_51),
.Y(n_179)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_59),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_67),
.B(n_71),
.C(n_74),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_73),
.B(n_196),
.C(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_74),
.B(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_78),
.B(n_122),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_95),
.C(n_111),
.Y(n_78)
);

XOR2x1_ASAP7_75t_L g286 ( 
.A(n_79),
.B(n_287),
.Y(n_286)
);

XOR2x1_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_86),
.C(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_94),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_86),
.A2(n_94),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_86),
.B(n_246),
.C(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_96),
.B(n_112),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.C(n_106),
.Y(n_96)
);

XOR2x1_ASAP7_75t_L g232 ( 
.A(n_97),
.B(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_101),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_102),
.Y(n_234)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_106),
.A2(n_107),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_116),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

XNOR2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_138),
.Y(n_122)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_134),
.C(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_130),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_159),
.C(n_160),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_157),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_173),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2x2_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_180),
.B1(n_184),
.B2(n_185),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_188),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_290),
.B(n_294),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_275),
.B(n_289),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_235),
.B(n_274),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_218),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_193),
.B(n_218),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.C(n_208),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_194),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_200),
.A2(n_201),
.B1(n_208),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_202),
.B(n_207),
.Y(n_251)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

AO22x1_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_216),
.Y(n_220)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_230),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_219),
.B(n_231),
.C(n_232),
.Y(n_288)
);

XOR2x1_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_268),
.B(n_273),
.Y(n_235)
);

OAI21x1_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_252),
.B(n_267),
.Y(n_236)
);

NOR2x1_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_243),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_250),
.B2(n_251),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI21x1_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_259),
.B(n_266),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

NOR2x1_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_272),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_288),
.Y(n_275)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_288),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_286),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_284),
.C(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_293),
.Y(n_294)
);


endmodule