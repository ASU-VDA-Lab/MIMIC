module real_jpeg_24011_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_1),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_158),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_158),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_35),
.B1(n_52),
.B2(n_53),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_2),
.A2(n_35),
.B1(n_69),
.B2(n_70),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_112),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_3),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_24),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_155),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_65),
.C(n_70),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_3),
.B(n_51),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_3),
.A2(n_89),
.B1(n_245),
.B2(n_252),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_6),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_149),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_6),
.A2(n_69),
.B1(n_70),
.B2(n_149),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_6),
.A2(n_111),
.B1(n_112),
.B2(n_149),
.Y(n_286)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_8),
.A2(n_33),
.B1(n_147),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_147),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_8),
.A2(n_69),
.B1(n_70),
.B2(n_147),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_9),
.A2(n_56),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_9),
.A2(n_56),
.B1(n_69),
.B2(n_70),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_10),
.A2(n_39),
.B1(n_52),
.B2(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_10),
.A2(n_39),
.B1(n_69),
.B2(n_70),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_12),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_12),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_73),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_73),
.Y(n_118)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_15),
.Y(n_141)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_19),
.B(n_105),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.C(n_85),
.Y(n_19)
);

FAx1_ASAP7_75t_L g328 ( 
.A(n_20),
.B(n_74),
.CI(n_85),
.CON(n_328),
.SN(n_328)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_43),
.B2(n_44),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_21),
.A2(n_22),
.B1(n_107),
.B2(n_120),
.Y(n_106)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_46),
.C(n_60),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B(n_36),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_23),
.B(n_38),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_23),
.A2(n_151),
.B1(n_152),
.B2(n_156),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_23),
.B(n_103),
.Y(n_305)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_24),
.A2(n_40),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_24),
.A2(n_40),
.B1(n_157),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_24),
.A2(n_40),
.B1(n_165),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_25),
.A2(n_26),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_25),
.A2(n_29),
.B(n_154),
.C(n_172),
.Y(n_171)
);

HAxp5_ASAP7_75t_SL g200 ( 
.A(n_25),
.B(n_155),
.CON(n_200),
.SN(n_200)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_26),
.B(n_28),
.C(n_167),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_26),
.A2(n_50),
.A3(n_53),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_29),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_31),
.Y(n_109)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_34),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_40),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_40),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_40),
.A2(n_286),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B(n_57),
.Y(n_46)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_47),
.B(n_59),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_47),
.A2(n_51),
.B1(n_191),
.B2(n_200),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_49),
.B(n_52),
.Y(n_201)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_51),
.B(n_118),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_53),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_53),
.B(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_58),
.A2(n_76),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_61),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_68),
.B(n_71),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_72),
.B(n_99),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_63),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_63),
.A2(n_81),
.B(n_207),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_63),
.A2(n_206),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_63),
.A2(n_205),
.B1(n_206),
.B2(n_225),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_63),
.A2(n_98),
.B1(n_206),
.B2(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_84),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_68),
.A2(n_82),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_68),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_68),
.B(n_155),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_69),
.B(n_256),
.Y(n_255)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_74),
.A2(n_75),
.B(n_79),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_78),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_76),
.A2(n_117),
.B(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_76),
.A2(n_78),
.B1(n_146),
.B2(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_77),
.A2(n_78),
.B(n_119),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_100),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_86),
.B(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_87),
.A2(n_88),
.B1(n_97),
.B2(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_87),
.A2(n_88),
.B1(n_100),
.B2(n_101),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B(n_95),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_89),
.A2(n_95),
.B(n_138),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_89),
.A2(n_235),
.B(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_89),
.A2(n_93),
.B1(n_242),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_90),
.A2(n_91),
.B1(n_137),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_90),
.B(n_139),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_90),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_93),
.B(n_155),
.Y(n_256)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_96),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_97),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_121),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_113),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_118),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_325),
.B(n_329),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_312),
.B(n_324),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_294),
.B(n_311),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_192),
.B(n_271),
.C(n_293),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_177),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_177),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_161),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_142),
.B1(n_159),
.B2(n_160),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_132),
.B(n_160),
.C(n_161),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_133),
.B(n_135),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_134),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_141),
.Y(n_237)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_150),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_170),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_164),
.B(n_168),
.C(n_170),
.Y(n_291)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_178),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_181),
.B(n_183),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_212),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_186),
.B(n_236),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_266),
.B(n_270),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_219),
.B(n_265),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_197),
.B(n_208),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.C(n_204),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_198),
.B(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_202),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_203),
.B(n_204),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_216),
.C(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_260),
.B(n_264),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_238),
.B(n_259),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_222),
.B(n_228),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_226),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_248),
.B(n_258),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_247),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_253),
.B(n_257),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_273),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_291),
.B2(n_292),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_282),
.C(n_292),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_281),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_279),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_287),
.C(n_290),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_296),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_310),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_300),
.B1(n_308),
.B2(n_309),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_309),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_304),
.C(n_306),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_314),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_322),
.B2(n_323),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_321),
.C(n_323),
.Y(n_327)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_327),
.B(n_328),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_328),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule