module fake_ariane_689_n_104 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_104);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_104;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_53;
wire n_66;
wire n_71;
wire n_96;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_91;
wire n_72;
wire n_82;
wire n_57;
wire n_70;
wire n_85;
wire n_94;
wire n_101;
wire n_58;
wire n_65;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_61;
wire n_102;
wire n_81;
wire n_87;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_78;
wire n_59;
wire n_63;
wire n_99;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

OR2x6_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_28),
.Y(n_60)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_49),
.B(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_0),
.B1(n_44),
.B2(n_31),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_46),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_18),
.B(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_1),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_8),
.Y(n_76)
);

OR2x6_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_14),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_15),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

AOI22x1_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_67),
.B1(n_70),
.B2(n_68),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_63),
.B1(n_56),
.B2(n_57),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_53),
.B(n_60),
.C(n_64),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_66),
.B1(n_58),
.B2(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_58),
.B1(n_20),
.B2(n_24),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_16),
.B(n_26),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_78),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_34),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_89),
.B1(n_93),
.B2(n_86),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);

AOI21x1_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_92),
.B(n_90),
.Y(n_102)
);

AOI222xp33_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_84),
.B1(n_87),
.B2(n_96),
.C1(n_47),
.C2(n_36),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_104)
);


endmodule