module fake_aes_9862_n_30 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_30);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_L g8 ( .A(n_4), .B(n_1), .Y(n_8) );
BUFx10_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
BUFx10_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
BUFx6f_ASAP7_75t_SL g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
OAI21x1_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_0), .B(n_1), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_10), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
AO32x2_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_5), .A3(n_6), .B1(n_7), .B2(n_13), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_10), .B(n_5), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_11), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_18), .B(n_15), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_20), .Y(n_24) );
AOI321xp33_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_17), .A3(n_8), .B1(n_18), .B2(n_19), .C(n_13), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_21), .B1(n_23), .B2(n_8), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_23), .B1(n_21), .B2(n_19), .C(n_9), .Y(n_27) );
AOI222xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_9), .B1(n_16), .B2(n_19), .C1(n_24), .C2(n_22), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_19), .B(n_28), .Y(n_30) );
endmodule