module fake_jpeg_208_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_34),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_39),
.B1(n_40),
.B2(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_38),
.B1(n_42),
.B2(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_45),
.B1(n_46),
.B2(n_3),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_67),
.Y(n_81)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_14),
.B1(n_27),
.B2(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_65),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_31),
.B(n_10),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_11),
.B(n_25),
.Y(n_88)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_9),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_83),
.C(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_3),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_94),
.B(n_24),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_6),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_74),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_100),
.B1(n_102),
.B2(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_16),
.B(n_19),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_22),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_107),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_93),
.B1(n_87),
.B2(n_23),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_98),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_109),
.B(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_115),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_118),
.B(n_104),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_110),
.Y(n_120)
);


endmodule