module fake_jpeg_958_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_81),
.Y(n_87)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_54),
.B1(n_71),
.B2(n_60),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_91),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_69),
.B1(n_66),
.B2(n_61),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_57),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_57),
.B1(n_71),
.B2(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_94),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_51),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_58),
.C(n_53),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_89),
.C(n_64),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_55),
.B(n_70),
.C(n_62),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_59),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_112),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_0),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_65),
.B(n_52),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_113),
.B1(n_90),
.B2(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_124),
.B1(n_44),
.B2(n_41),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_90),
.B1(n_69),
.B2(n_60),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_96),
.B(n_90),
.C(n_72),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_23),
.B(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_67),
.B(n_63),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_46),
.B(n_45),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_0),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_48),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_29),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_72),
.B1(n_67),
.B2(n_47),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_33),
.B1(n_31),
.B2(n_30),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_7),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_142),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_149),
.B(n_153),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_146),
.B1(n_149),
.B2(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_39),
.C(n_38),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_14),
.C(n_15),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_36),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_1),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_2),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_4),
.B(n_5),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_158),
.B(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_5),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_6),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_6),
.B(n_7),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_8),
.B(n_10),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_134),
.B(n_117),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_173),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_168),
.B(n_170),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_166),
.B(n_172),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_132),
.B(n_9),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_8),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_158),
.B(n_140),
.C(n_145),
.D(n_149),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_15),
.C(n_16),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_154),
.B1(n_153),
.B2(n_160),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_163),
.B1(n_161),
.B2(n_178),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_16),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_17),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_193),
.B1(n_195),
.B2(n_192),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_161),
.B1(n_163),
.B2(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

AOI31xp67_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_178),
.A3(n_183),
.B(n_169),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_187),
.B(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_197),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_188),
.C(n_180),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_180),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_200),
.A2(n_165),
.B1(n_177),
.B2(n_20),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_203),
.B(n_165),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_176),
.B(n_199),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_201),
.C(n_17),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_19),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_19),
.Y(n_208)
);


endmodule