module fake_jpeg_31769_n_438 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_438);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_65),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_66),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_14),
.CON(n_58),
.SN(n_58)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_89),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_31),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_71),
.Y(n_112)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_31),
.B(n_0),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_88),
.Y(n_100)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_81),
.Y(n_115)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_90),
.Y(n_128)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_85),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_86),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_87),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_19),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_42),
.B1(n_43),
.B2(n_39),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_92),
.A2(n_116),
.B1(n_134),
.B2(n_2),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_58),
.B(n_35),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_121),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_42),
.B1(n_18),
.B2(n_43),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_108),
.A2(n_117),
.B1(n_129),
.B2(n_131),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_54),
.B1(n_85),
.B2(n_56),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_59),
.A2(n_18),
.B1(n_43),
.B2(n_39),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_61),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_48),
.A2(n_27),
.B1(n_39),
.B2(n_41),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_125),
.A2(n_141),
.B1(n_4),
.B2(n_9),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_49),
.A2(n_27),
.B1(n_46),
.B2(n_44),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_57),
.A2(n_46),
.B1(n_37),
.B2(n_38),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_41),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_67),
.A2(n_37),
.B1(n_38),
.B2(n_34),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_29),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_70),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_73),
.B1(n_82),
.B2(n_76),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_143),
.A2(n_152),
.B1(n_166),
.B2(n_186),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_100),
.A2(n_84),
.B(n_36),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_144),
.A2(n_130),
.B(n_114),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_79),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_146),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_36),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_36),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_159),
.Y(n_197)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_110),
.A2(n_81),
.B1(n_36),
.B2(n_72),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_154),
.Y(n_215)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_95),
.A2(n_36),
.B1(n_33),
.B2(n_3),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_176),
.B(n_12),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_111),
.B1(n_98),
.B2(n_101),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_158),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_95),
.B(n_4),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_136),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_162),
.C(n_181),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_33),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_104),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_164),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_4),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_96),
.A2(n_33),
.B1(n_5),
.B2(n_6),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_103),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_171),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_112),
.A2(n_128),
.B(n_115),
.C(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_174),
.Y(n_190)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_115),
.A2(n_33),
.B1(n_5),
.B2(n_6),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_182),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_180),
.A2(n_187),
.B1(n_118),
.B2(n_126),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_4),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_121),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_114),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_96),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_14),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_191),
.B(n_218),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_193),
.A2(n_194),
.B1(n_210),
.B2(n_161),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_111),
.B1(n_98),
.B2(n_132),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_159),
.B(n_185),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_156),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_99),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_130),
.C(n_137),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_224),
.C(n_162),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_146),
.B(n_113),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_113),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_160),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_137),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_172),
.B1(n_154),
.B2(n_162),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_132),
.B1(n_126),
.B2(n_105),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_222),
.A2(n_229),
.B1(n_154),
.B2(n_175),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_160),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_226),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_124),
.C(n_135),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_163),
.B(n_124),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_151),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_181),
.A2(n_135),
.B1(n_93),
.B2(n_140),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_248),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_239),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_181),
.B1(n_176),
.B2(n_147),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_232),
.Y(n_282)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_234),
.A2(n_264),
.B(n_190),
.C(n_195),
.D(n_198),
.Y(n_292)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_238),
.B(n_256),
.C(n_213),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_183),
.C(n_169),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_240),
.A2(n_254),
.B1(n_261),
.B2(n_231),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_199),
.A2(n_182),
.B1(n_155),
.B2(n_171),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_241),
.A2(n_204),
.B1(n_226),
.B2(n_227),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_253),
.Y(n_267)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_150),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_250),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_167),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_222),
.B1(n_210),
.B2(n_229),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_192),
.B(n_170),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_192),
.B(n_197),
.CI(n_205),
.CON(n_255),
.SN(n_255)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_258),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_173),
.C(n_174),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_191),
.B(n_142),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_259),
.B(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_205),
.B(n_93),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_223),
.B(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_179),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_197),
.B(n_179),
.Y(n_263)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_211),
.A2(n_149),
.A3(n_179),
.B1(n_212),
.B2(n_219),
.Y(n_264)
);

INVx2_ASAP7_75t_R g265 ( 
.A(n_218),
.Y(n_265)
);

OAI21x1_ASAP7_75t_R g294 ( 
.A1(n_265),
.A2(n_215),
.B(n_196),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_272),
.A2(n_286),
.B1(n_291),
.B2(n_282),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_216),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_280),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_277),
.A2(n_286),
.B(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_209),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_247),
.B(n_207),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_285),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_297),
.C(n_238),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_207),
.Y(n_285)
);

OAI22x1_ASAP7_75t_L g286 ( 
.A1(n_239),
.A2(n_200),
.B1(n_194),
.B2(n_193),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_189),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_293),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_236),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_251),
.A2(n_198),
.B1(n_215),
.B2(n_206),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_240),
.B1(n_260),
.B2(n_259),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_292),
.A2(n_232),
.B(n_234),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_233),
.B(n_206),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_298),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_265),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_246),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_196),
.C(n_202),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_268),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_299),
.B(n_300),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_268),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_327),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_255),
.C(n_256),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_261),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_309),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_263),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_247),
.C(n_262),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_231),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_313),
.Y(n_340)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_264),
.C(n_232),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_316),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_294),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_235),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_319),
.Y(n_345)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_237),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_288),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_324),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_296),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_326),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_275),
.Y(n_336)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_302),
.A2(n_282),
.B1(n_272),
.B2(n_292),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_338),
.A2(n_349),
.B1(n_352),
.B2(n_305),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_302),
.A2(n_279),
.B(n_298),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_314),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_344),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_293),
.Y(n_342)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_267),
.Y(n_343)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_301),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_270),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_321),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_279),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_351),
.A2(n_303),
.B(n_267),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_302),
.A2(n_281),
.B1(n_284),
.B2(n_232),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_308),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_356),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_354),
.A2(n_337),
.B1(n_338),
.B2(n_333),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_332),
.A2(n_327),
.B1(n_317),
.B2(n_319),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_355),
.A2(n_360),
.B1(n_352),
.B2(n_349),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_340),
.B(n_309),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_306),
.C(n_310),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_368),
.C(n_370),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_347),
.A2(n_271),
.B1(n_331),
.B2(n_329),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_311),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_362),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_313),
.Y(n_362)
);

NAND2x1_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_303),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_365),
.B(n_373),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_366),
.A2(n_351),
.B(n_336),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_321),
.Y(n_370)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_334),
.B(n_280),
.CI(n_287),
.CON(n_371),
.SN(n_371)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_371),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_276),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_375),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_383),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_358),
.A2(n_350),
.B1(n_346),
.B2(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_369),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_379),
.B(n_269),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_328),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_380),
.Y(n_391)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_SL g387 ( 
.A1(n_365),
.A2(n_343),
.B(n_342),
.C(n_345),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_387),
.A2(n_243),
.B(n_295),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_364),
.A2(n_345),
.B1(n_346),
.B2(n_331),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_243),
.Y(n_400)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

AO221x1_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_326),
.B1(n_318),
.B2(n_312),
.C(n_372),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_370),
.C(n_357),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_394),
.C(n_397),
.Y(n_403)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_362),
.C(n_353),
.Y(n_394)
);

OAI321xp33_ASAP7_75t_L g395 ( 
.A1(n_382),
.A2(n_371),
.A3(n_355),
.B1(n_364),
.B2(n_368),
.C(n_373),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_399),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_356),
.C(n_361),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_380),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_402),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_273),
.Y(n_411)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_391),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_408),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_386),
.C(n_388),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_402),
.B(n_396),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_377),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_381),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_413),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_412),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_398),
.B(n_385),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_269),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_385),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_394),
.C(n_384),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_421),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_416),
.A2(n_417),
.B(n_422),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_405),
.A2(n_384),
.B(n_387),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_400),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_419),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_269),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_406),
.A2(n_403),
.B(n_407),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_420),
.A2(n_403),
.B(n_414),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_425),
.B(n_426),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_407),
.B1(n_387),
.B2(n_295),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_419),
.A2(n_387),
.B1(n_257),
.B2(n_244),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_423),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_431),
.B(n_432),
.Y(n_435)
);

OAI321xp33_ASAP7_75t_L g432 ( 
.A1(n_424),
.A2(n_428),
.A3(n_423),
.B1(n_429),
.B2(n_273),
.C(n_245),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_SL g433 ( 
.A(n_429),
.B(n_273),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_227),
.C(n_273),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_434),
.Y(n_436)
);

NOR3xp33_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_435),
.C(n_430),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_245),
.Y(n_438)
);


endmodule