module fake_jpeg_11048_n_564 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_564);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_564;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_20),
.B(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_79),
.B(n_90),
.Y(n_153)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_40),
.B(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_40),
.Y(n_156)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_103),
.Y(n_165)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_156),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_50),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_113),
.B(n_118),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_75),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_116),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_50),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_120),
.B(n_121),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_19),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_37),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_33),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_60),
.A2(n_19),
.B1(n_46),
.B2(n_45),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_49),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_162),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_62),
.B(n_49),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_96),
.B(n_19),
.C(n_44),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_25),
.C(n_36),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_108),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_170),
.B(n_145),
.C(n_136),
.Y(n_250)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_172),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_208),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_174),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_46),
.B1(n_45),
.B2(n_38),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_175),
.A2(n_181),
.B1(n_184),
.B2(n_190),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_121),
.A2(n_84),
.B1(n_72),
.B2(n_70),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_176),
.A2(n_182),
.B1(n_216),
.B2(n_226),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_38),
.B(n_30),
.C(n_28),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_177),
.B(n_186),
.Y(n_235)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_180),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_46),
.B1(n_30),
.B2(n_28),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_102),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_83),
.B1(n_93),
.B2(n_85),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_108),
.A2(n_26),
.B(n_38),
.C(n_30),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

BUFx4f_ASAP7_75t_SL g256 ( 
.A(n_188),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_189),
.A2(n_195),
.B(n_202),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_112),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_191),
.A2(n_196),
.B1(n_207),
.B2(n_224),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_61),
.B1(n_76),
.B2(n_74),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_192),
.A2(n_200),
.B1(n_14),
.B2(n_16),
.Y(n_282)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_115),
.B(n_101),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_141),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_139),
.A2(n_66),
.B(n_65),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_0),
.Y(n_260)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_137),
.A2(n_59),
.B1(n_44),
.B2(n_43),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_124),
.B(n_0),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_132),
.B(n_134),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_229),
.Y(n_238)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_165),
.A2(n_25),
.B1(n_36),
.B2(n_34),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_211),
.B(n_213),
.Y(n_271)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_43),
.B1(n_34),
.B2(n_2),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_219),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g218 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g269 ( 
.A1(n_218),
.A2(n_6),
.B1(n_8),
.B2(n_13),
.Y(n_269)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_221),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_122),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_119),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_223),
.Y(n_263)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_138),
.A2(n_10),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_225),
.B(n_227),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_150),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_151),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_110),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_230),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_127),
.B(n_12),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_140),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_111),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_173),
.B(n_163),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_239),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_170),
.B(n_199),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_149),
.B1(n_163),
.B2(n_135),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_243),
.A2(n_247),
.B1(n_254),
.B2(n_262),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_185),
.A2(n_126),
.B(n_136),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_246),
.A2(n_221),
.B(n_231),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_215),
.A2(n_135),
.B1(n_111),
.B2(n_131),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_178),
.B(n_13),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_250),
.C(n_279),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_188),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_252),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_189),
.A2(n_145),
.B1(n_0),
.B2(n_5),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_204),
.A2(n_12),
.B(n_4),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_272),
.B(n_195),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_260),
.B(n_172),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_261),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_184),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_177),
.B(n_186),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_268),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_216),
.A2(n_225),
.B1(n_193),
.B2(n_218),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_266),
.A2(n_267),
.B1(n_273),
.B2(n_282),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_218),
.A2(n_6),
.B1(n_8),
.B2(n_12),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_6),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_269),
.B(n_267),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_202),
.A2(n_6),
.B(n_8),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_218),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_187),
.B(n_13),
.C(n_14),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_206),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_211),
.B(n_16),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_284),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_220),
.B1(n_214),
.B2(n_213),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_SL g292 ( 
.A1(n_264),
.A2(n_218),
.B(n_183),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_292),
.A2(n_301),
.B(n_252),
.Y(n_362)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_295),
.Y(n_361)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_223),
.B1(n_231),
.B2(n_228),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_299),
.A2(n_303),
.B1(n_306),
.B2(n_308),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_263),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_219),
.B1(n_205),
.B2(n_179),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_235),
.A2(n_180),
.B1(n_171),
.B2(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_271),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_307),
.B(n_309),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_275),
.A2(n_222),
.B1(n_194),
.B2(n_212),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_271),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_310),
.B(n_314),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_198),
.B(n_195),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_316),
.B(n_319),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_245),
.A2(n_217),
.B1(n_208),
.B2(n_201),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_315),
.B1(n_324),
.B2(n_281),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_253),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_325),
.Y(n_342)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_266),
.A2(n_234),
.B1(n_236),
.B2(n_238),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_233),
.A2(n_236),
.B(n_250),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_239),
.B(n_233),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_321),
.C(n_254),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_233),
.A2(n_246),
.B(n_272),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_320),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_260),
.B(n_259),
.C(n_248),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_242),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_322),
.B(n_255),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_243),
.A2(n_232),
.B1(n_257),
.B2(n_262),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_268),
.A2(n_269),
.B(n_279),
.C(n_242),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_270),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_327),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_269),
.A3(n_258),
.B1(n_263),
.B2(n_247),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_244),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_244),
.A2(n_270),
.B1(n_255),
.B2(n_240),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_256),
.B(n_312),
.Y(n_370)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_273),
.B(n_232),
.CI(n_269),
.CON(n_335),
.SN(n_335)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_281),
.C(n_277),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_283),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_340),
.C(n_344),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_258),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_287),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_343),
.B(n_353),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_289),
.B(n_276),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_347),
.B(n_366),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_240),
.C(n_277),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_349),
.B(n_357),
.C(n_368),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_321),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_302),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_286),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_354),
.B(n_375),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_355),
.A2(n_374),
.B(n_301),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_276),
.C(n_265),
.Y(n_357)
);

OAI32xp33_ASAP7_75t_L g396 ( 
.A1(n_358),
.A2(n_307),
.A3(n_300),
.B1(n_326),
.B2(n_333),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_265),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_364),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_304),
.B(n_237),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_365),
.A2(n_378),
.B1(n_379),
.B2(n_318),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_296),
.B(n_237),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_296),
.B(n_256),
.C(n_300),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_333),
.C(n_313),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_370),
.A2(n_337),
.B(n_374),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_329),
.A2(n_256),
.B1(n_318),
.B2(n_327),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_352),
.B1(n_351),
.B2(n_358),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_319),
.A2(n_256),
.B(n_305),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_291),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_293),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_295),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_325),
.Y(n_377)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_324),
.A2(n_303),
.B1(n_335),
.B2(n_306),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_335),
.A2(n_323),
.B1(n_332),
.B2(n_311),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_381),
.A2(n_384),
.B1(n_389),
.B2(n_405),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_372),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_379),
.A2(n_378),
.B1(n_352),
.B2(n_365),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_364),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_388),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_387),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_363),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_329),
.B1(n_314),
.B2(n_310),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_390),
.A2(n_400),
.B(n_412),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_373),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_393),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_355),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_376),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_394),
.B(n_396),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_345),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_403),
.C(n_407),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_337),
.A2(n_289),
.B1(n_313),
.B2(n_331),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_290),
.C(n_330),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_404),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_342),
.A2(n_294),
.B1(n_309),
.B2(n_320),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_367),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_341),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_339),
.C(n_350),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_377),
.A2(n_328),
.B1(n_351),
.B2(n_359),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_415),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_357),
.Y(n_409)
);

NAND3xp33_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_414),
.C(n_416),
.Y(n_426)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_411),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_344),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_362),
.C(n_346),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_371),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_348),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_349),
.Y(n_416)
);

OAI21x1_ASAP7_75t_SL g452 ( 
.A1(n_418),
.A2(n_382),
.B(n_412),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_420),
.B(n_434),
.C(n_440),
.Y(n_450)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_427),
.B(n_441),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_394),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_428),
.B(n_435),
.Y(n_458)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_411),
.Y(n_429)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_429),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_346),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_402),
.B(n_361),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_436),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_361),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_444),
.Y(n_463)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_380),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_439),
.B(n_418),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_370),
.C(n_338),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_401),
.B(n_391),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_392),
.A2(n_360),
.B(n_338),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_442),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_359),
.C(n_356),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_447),
.C(n_403),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_385),
.B(n_356),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_401),
.B(n_402),
.Y(n_446)
);

OAI22xp33_ASAP7_75t_SL g475 ( 
.A1(n_446),
.A2(n_449),
.B1(n_425),
.B2(n_438),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_397),
.B(n_385),
.C(n_399),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_383),
.B(n_388),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_420),
.B(n_397),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_451),
.B(n_465),
.Y(n_487)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_452),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_381),
.B1(n_384),
.B2(n_408),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_456),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_423),
.A2(n_393),
.B1(n_386),
.B2(n_390),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_421),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_461),
.C(n_437),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_419),
.B(n_392),
.C(n_389),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_445),
.A2(n_400),
.B(n_396),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_462),
.B(n_466),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_380),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_445),
.A2(n_405),
.B(n_433),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_423),
.A2(n_448),
.B1(n_421),
.B2(n_439),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_470),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_436),
.Y(n_470)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_472),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_429),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_473),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_448),
.A2(n_449),
.B1(n_446),
.B2(n_440),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_474),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_475),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_419),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_417),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_479),
.C(n_489),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_447),
.C(n_443),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_426),
.Y(n_481)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_471),
.B(n_430),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_460),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_454),
.A2(n_433),
.B(n_442),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_486),
.A2(n_462),
.B(n_464),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_474),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_424),
.C(n_422),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_424),
.C(n_422),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_499),
.C(n_500),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_417),
.Y(n_494)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_494),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_432),
.Y(n_498)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_498),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_435),
.C(n_450),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_450),
.C(n_465),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_480),
.B1(n_469),
.B2(n_491),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_502),
.A2(n_508),
.B1(n_495),
.B2(n_483),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_490),
.A2(n_453),
.B1(n_456),
.B2(n_470),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_503),
.A2(n_507),
.B1(n_483),
.B2(n_486),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_505),
.B(n_511),
.Y(n_533)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_506),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_490),
.A2(n_472),
.B1(n_459),
.B2(n_466),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_493),
.A2(n_455),
.B1(n_473),
.B2(n_458),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_452),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_496),
.Y(n_512)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_512),
.Y(n_526)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_496),
.Y(n_513)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_513),
.Y(n_519)
);

NOR2x1_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_458),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_514),
.A2(n_515),
.B(n_468),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_485),
.A2(n_451),
.B(n_464),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_487),
.Y(n_530)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_489),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_521),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g522 ( 
.A(n_501),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_522),
.B(n_523),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_510),
.B(n_500),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_525),
.B(n_527),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_492),
.C(n_479),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_529),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_488),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_511),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_508),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_531),
.B(n_532),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_478),
.C(n_487),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_525),
.A2(n_502),
.B1(n_515),
.B2(n_503),
.Y(n_535)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_535),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_533),
.Y(n_548)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_519),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_541),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_505),
.C(n_507),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_509),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_543),
.B(n_544),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_504),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_536),
.A2(n_527),
.B(n_514),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_545),
.A2(n_546),
.B(n_539),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_542),
.A2(n_519),
.B(n_526),
.Y(n_546)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_548),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_520),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_538),
.Y(n_552)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_552),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_554),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_550),
.B(n_534),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_555),
.B(n_549),
.C(n_547),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_557),
.A2(n_541),
.B(n_558),
.Y(n_560)
);

AOI21xp33_ASAP7_75t_L g559 ( 
.A1(n_556),
.A2(n_545),
.B(n_548),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_559),
.A2(n_560),
.B(n_537),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_561),
.B(n_535),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_468),
.B1(n_530),
.B2(n_533),
.Y(n_563)
);

BUFx24_ASAP7_75t_SL g564 ( 
.A(n_563),
.Y(n_564)
);


endmodule