module real_jpeg_11665_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_286, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_286;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_176;
wire n_215;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_244;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_0),
.A2(n_41),
.B1(n_59),
.B2(n_60),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_0),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_223)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B(n_282),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_4),
.B(n_283),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_27),
.B1(n_47),
.B2(n_48),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_27),
.B1(n_59),
.B2(n_60),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_9),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_11),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_12),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_12),
.A2(n_33),
.B(n_44),
.C(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_12),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_12),
.B(n_38),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_12),
.B(n_57),
.C(n_60),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_12),
.B(n_49),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_30),
.C(n_34),
.Y(n_167)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_76),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_74),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_71),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_71),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_65),
.C(n_68),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_19),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.C(n_52),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_20),
.A2(n_117),
.B1(n_119),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_20),
.B(n_117),
.C(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_20),
.A2(n_85),
.B1(n_86),
.B2(n_182),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_20),
.A2(n_182),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_36),
.B2(n_38),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_22),
.A2(n_32),
.B(n_70),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_24),
.B(n_167),
.Y(n_166)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_36),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_28),
.B(n_38),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_32),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_36),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_37),
.A2(n_45),
.B(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_37),
.B(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_37),
.B(n_63),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_39),
.A2(n_52),
.B1(n_257),
.B2(n_271),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_39),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_39)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_40),
.Y(n_259)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_42),
.A2(n_49),
.B1(n_89),
.B2(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_46),
.A2(n_67),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_46),
.A2(n_88),
.B(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_48),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_52),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_52),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_52),
.B(n_170),
.C(n_258),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_63),
.B(n_64),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_53),
.A2(n_63),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_94),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_54),
.A2(n_58),
.B1(n_92),
.B2(n_94),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_54),
.A2(n_58),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_59),
.B(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_91),
.B(n_93),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_63),
.A2(n_93),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_64),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_65),
.B(n_68),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_277),
.B(n_281),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_249),
.B(n_274),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_227),
.B(n_248),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_210),
.B(n_226),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_177),
.A3(n_205),
.B1(n_208),
.B2(n_209),
.C(n_286),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_159),
.B(n_176),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_125),
.B(n_158),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_106),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_84),
.B(n_106),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_95),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_142),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_85),
.A2(n_86),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_86),
.B(n_169),
.C(n_174),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_86),
.B(n_182),
.C(n_215),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_89),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_129),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_90),
.A2(n_142),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_95),
.A2(n_96),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_101),
.B(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_104),
.A2(n_105),
.B1(n_185),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_105),
.A2(n_115),
.B(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_120),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_122),
.C(n_123),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_117),
.B2(n_119),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_113),
.C(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_117),
.A2(n_243),
.B(n_246),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_117),
.B(n_243),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_124),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_134),
.C(n_136),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_122),
.A2(n_124),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_202),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_152),
.B(n_157),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_138),
.B(n_151),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_131),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_136),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_148),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_165),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_143),
.B(n_150),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_184),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_147),
.B(n_149),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_164),
.C(n_168),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_170),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_192),
.C(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_169),
.A2(n_170),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_169),
.A2(n_170),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_170),
.B(n_268),
.C(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_187),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_183),
.CI(n_187),
.CON(n_207),
.SN(n_207)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_184),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_204),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_199),
.B2(n_200),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_200),
.C(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_206),
.B(n_207),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_207),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_225),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_225),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_214),
.C(n_219),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_220),
.A2(n_224),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_233),
.B(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_229),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_247),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_241),
.B2(n_242),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_241),
.C(n_247),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_253),
.B1(n_254),
.B2(n_261),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_264),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_263),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_263),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_261),
.C(n_262),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_258),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_273),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_280),
.Y(n_281)
);


endmodule