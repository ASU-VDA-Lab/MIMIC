module fake_jpeg_12902_n_535 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_535);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_69),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g178 ( 
.A(n_71),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_18),
.B(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_77),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_0),
.CON(n_73),
.SN(n_73)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_73),
.B(n_75),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_54),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_29),
.B(n_7),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_89),
.Y(n_133)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx9p33_ASAP7_75t_R g171 ( 
.A(n_87),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_7),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_6),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_110),
.Y(n_139)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_6),
.C(n_1),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_39),
.C(n_28),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_35),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_100),
.A2(n_25),
.B1(n_58),
.B2(n_52),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

CKINVDCx9p33_ASAP7_75t_R g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_106),
.Y(n_192)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_10),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_11),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_122),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_40),
.Y(n_113)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_123),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_28),
.B(n_53),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_35),
.B1(n_57),
.B2(n_45),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_126),
.A2(n_146),
.B1(n_156),
.B2(n_179),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_49),
.B1(n_51),
.B2(n_35),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_135),
.A2(n_143),
.B(n_155),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_138),
.B(n_152),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_76),
.A2(n_49),
.B1(n_51),
.B2(n_57),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_90),
.A2(n_25),
.B1(n_45),
.B2(n_59),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_33),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_149),
.B(n_151),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_33),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_114),
.A2(n_51),
.B1(n_31),
.B2(n_36),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_39),
.B1(n_50),
.B2(n_56),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_93),
.A2(n_120),
.B1(n_97),
.B2(n_108),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_157),
.A2(n_193),
.B1(n_196),
.B2(n_34),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_50),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_159),
.B(n_165),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_78),
.B(n_53),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_60),
.B(n_55),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_173),
.B(n_183),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_73),
.A2(n_31),
.B1(n_58),
.B2(n_52),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_55),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_61),
.B(n_56),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_189),
.B(n_200),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_98),
.A2(n_26),
.B1(n_47),
.B2(n_42),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_63),
.A2(n_47),
.B1(n_42),
.B2(n_36),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_27),
.B1(n_80),
.B2(n_34),
.Y(n_221)
);

AOI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_71),
.A2(n_34),
.B(n_4),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_12),
.B(n_4),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_62),
.B(n_32),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_201),
.Y(n_317)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_203),
.Y(n_306)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

BUFx4f_ASAP7_75t_SL g283 ( 
.A(n_205),
.Y(n_283)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_207),
.B(n_229),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_59),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_235),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_87),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_210),
.B(n_212),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_32),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_213),
.Y(n_278)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_215),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_179),
.A2(n_122),
.B1(n_101),
.B2(n_85),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_216),
.A2(n_230),
.B1(n_253),
.B2(n_258),
.Y(n_280)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_232),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_192),
.A2(n_27),
.B1(n_67),
.B2(n_84),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_223),
.A2(n_242),
.B1(n_245),
.B2(n_251),
.Y(n_289)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_225),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_167),
.A2(n_83),
.B1(n_69),
.B2(n_68),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_226),
.A2(n_228),
.B1(n_233),
.B2(n_237),
.Y(n_272)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_227),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_126),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_231),
.B(n_249),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_139),
.B(n_5),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_234),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_133),
.B(n_5),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_157),
.A2(n_146),
.B1(n_177),
.B2(n_166),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_141),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_239),
.B(n_257),
.Y(n_282)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_130),
.A2(n_143),
.B1(n_135),
.B2(n_174),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_240),
.A2(n_243),
.B(n_210),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_134),
.B(n_13),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_261),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_150),
.A2(n_13),
.B1(n_15),
.B2(n_136),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_130),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_248),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_124),
.Y(n_245)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_176),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_246),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_129),
.A2(n_13),
.B1(n_160),
.B2(n_142),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_264),
.B1(n_172),
.B2(n_137),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_154),
.B(n_130),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_125),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_250),
.B(n_252),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_150),
.A2(n_128),
.B1(n_158),
.B2(n_145),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_155),
.A2(n_170),
.B1(n_180),
.B2(n_131),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_144),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_254),
.B(n_256),
.Y(n_298)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_164),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_129),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_161),
.A2(n_169),
.B1(n_163),
.B2(n_144),
.Y(n_258)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_162),
.A2(n_198),
.B1(n_195),
.B2(n_194),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_260),
.A2(n_265),
.B1(n_244),
.B2(n_266),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_161),
.B(n_169),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_163),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_263),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_162),
.A2(n_198),
.B1(n_195),
.B2(n_182),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_172),
.A2(n_186),
.B1(n_184),
.B2(n_127),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_266),
.B(n_268),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_137),
.B(n_127),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_267),
.B(n_207),
.Y(n_287)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_184),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_305),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_127),
.B(n_184),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_291),
.B(n_318),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_228),
.A2(n_243),
.B1(n_208),
.B2(n_262),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_292),
.B1(n_308),
.B2(n_311),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_287),
.B(n_320),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_241),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_307),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g302 ( 
.A1(n_220),
.A2(n_240),
.B1(n_229),
.B2(n_230),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_302),
.A2(n_311),
.B(n_246),
.C(n_268),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_261),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_212),
.B(n_235),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_312),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_213),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_271),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_240),
.B(n_222),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_236),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_262),
.A2(n_210),
.B1(n_218),
.B2(n_232),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_255),
.B1(n_263),
.B2(n_202),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_232),
.B(n_218),
.CI(n_224),
.CON(n_314),
.SN(n_314)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_314),
.B(n_209),
.CI(n_234),
.CON(n_338),
.SN(n_338)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_211),
.B(n_225),
.C(n_217),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_284),
.C(n_281),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_267),
.A2(n_250),
.B(n_257),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_214),
.B(n_238),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_301),
.B(n_204),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_323),
.B(n_344),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_316),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_326),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_316),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_327),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_215),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_357),
.C(n_358),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_316),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_329),
.B(n_336),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_307),
.A2(n_254),
.B1(n_245),
.B2(n_205),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_332),
.A2(n_350),
.B1(n_351),
.B2(n_303),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_297),
.B(n_259),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_333),
.B(n_352),
.Y(n_393)
);

OA22x2_ASAP7_75t_L g372 ( 
.A1(n_335),
.A2(n_300),
.B1(n_296),
.B2(n_306),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_298),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_312),
.B(n_206),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_337),
.B(n_338),
.Y(n_363)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_201),
.B1(n_203),
.B2(n_227),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_340),
.A2(n_343),
.B1(n_349),
.B2(n_359),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_252),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_300),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_285),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_346),
.B(n_347),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_295),
.B(n_269),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_282),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_348),
.B(n_354),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_287),
.A2(n_290),
.B1(n_275),
.B2(n_289),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_280),
.A2(n_302),
.B1(n_282),
.B2(n_311),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_280),
.A2(n_302),
.B1(n_311),
.B2(n_305),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_271),
.Y(n_353)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_353),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_273),
.B(n_270),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_304),
.A2(n_311),
.B(n_272),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_342),
.B(n_352),
.Y(n_370)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_269),
.C(n_313),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_284),
.C(n_294),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_284),
.A2(n_299),
.B1(n_279),
.B2(n_319),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_286),
.Y(n_360)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_275),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_361),
.A2(n_290),
.B(n_309),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_314),
.B(n_294),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_276),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_343),
.A2(n_288),
.B1(n_279),
.B2(n_299),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_365),
.A2(n_373),
.B1(n_374),
.B2(n_380),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_366),
.B(n_327),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_369),
.A2(n_375),
.B1(n_385),
.B2(n_386),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_372),
.B(n_342),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_371),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_344),
.A2(n_288),
.B1(n_319),
.B2(n_293),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_288),
.B1(n_293),
.B2(n_296),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_276),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_377),
.A2(n_324),
.B(n_326),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_378),
.B(n_379),
.Y(n_411)
);

NOR2x1_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_317),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_334),
.A2(n_336),
.B1(n_355),
.B2(n_331),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_277),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_381),
.B(n_382),
.C(n_390),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_333),
.B(n_277),
.C(n_306),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_328),
.B(n_321),
.C(n_303),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_355),
.A2(n_283),
.B1(n_317),
.B2(n_334),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_391),
.A2(n_341),
.B1(n_322),
.B2(n_335),
.Y(n_418)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_395),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_283),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_341),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_362),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_421),
.C(n_368),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_366),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_412),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_330),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_400),
.B(n_401),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_330),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_395),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_402),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_345),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_403),
.B(n_405),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_323),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_406),
.A2(n_397),
.B1(n_399),
.B2(n_423),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_407),
.A2(n_420),
.B(n_377),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_410),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_371),
.Y(n_440)
);

OAI32xp33_ASAP7_75t_L g410 ( 
.A1(n_363),
.A2(n_361),
.A3(n_331),
.B1(n_351),
.B2(n_354),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_384),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_414),
.Y(n_438)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_417),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_363),
.B(n_338),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_418),
.A2(n_422),
.B1(n_424),
.B2(n_335),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_339),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_423),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_370),
.A2(n_358),
.B(n_329),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_359),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_364),
.A2(n_322),
.B1(n_335),
.B2(n_325),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_377),
.A2(n_322),
.B1(n_335),
.B2(n_332),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_422),
.A2(n_369),
.B1(n_375),
.B2(n_389),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_432),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_427),
.A2(n_436),
.B(n_417),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_428),
.B(n_433),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_391),
.B1(n_365),
.B2(n_373),
.Y(n_429)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_381),
.C(n_393),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_434),
.C(n_441),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_404),
.A2(n_382),
.B1(n_372),
.B2(n_390),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_421),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_378),
.C(n_396),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_407),
.A2(n_372),
.B(n_371),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_440),
.B(n_434),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_338),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_443),
.A2(n_419),
.B1(n_415),
.B2(n_414),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_383),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_444),
.B(n_449),
.C(n_397),
.Y(n_452)
);

OAI21xp33_ASAP7_75t_L g446 ( 
.A1(n_411),
.A2(n_372),
.B(n_383),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_424),
.A2(n_394),
.B1(n_388),
.B2(n_376),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_406),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_388),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_466),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_401),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_453),
.B(n_437),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_435),
.A2(n_403),
.B(n_418),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_454),
.A2(n_465),
.B(n_445),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_404),
.B1(n_400),
.B2(n_408),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_456),
.A2(n_463),
.B1(n_437),
.B2(n_442),
.Y(n_479)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_438),
.Y(n_459)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_405),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_460),
.Y(n_486)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_426),
.B(n_448),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_416),
.C(n_411),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_431),
.C(n_440),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_417),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_416),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_468),
.A2(n_427),
.B(n_436),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_469),
.A2(n_447),
.B1(n_425),
.B2(n_430),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_356),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_472),
.B(n_479),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_473),
.A2(n_457),
.B1(n_450),
.B2(n_458),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_475),
.A2(n_484),
.B(n_468),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_477),
.C(n_478),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_432),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_449),
.C(n_435),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_441),
.Y(n_480)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_480),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_439),
.C(n_442),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_485),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_445),
.C(n_394),
.Y(n_485)
);

OAI21xp33_ASAP7_75t_L g495 ( 
.A1(n_487),
.A2(n_461),
.B(n_460),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_494),
.Y(n_507)
);

AO221x1_ASAP7_75t_L g491 ( 
.A1(n_474),
.A2(n_454),
.B1(n_462),
.B2(n_459),
.C(n_450),
.Y(n_491)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_481),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_496),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_360),
.Y(n_511)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_473),
.A2(n_456),
.B(n_457),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_497),
.A2(n_451),
.B1(n_476),
.B2(n_477),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_455),
.B1(n_463),
.B2(n_452),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_500),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_483),
.A2(n_455),
.B1(n_469),
.B2(n_465),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_497),
.A2(n_475),
.B1(n_478),
.B2(n_485),
.Y(n_501)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_501),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_471),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_503),
.B(n_508),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_505),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_471),
.C(n_487),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_488),
.C(n_490),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_493),
.B(n_466),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_353),
.C(n_376),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_502),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_502),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_493),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_513),
.C(n_500),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_498),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_519),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_518),
.A2(n_520),
.B1(n_509),
.B2(n_501),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_509),
.A2(n_504),
.B1(n_491),
.B2(n_494),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_521),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_517),
.A2(n_488),
.B(n_506),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_522),
.B(n_526),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_516),
.A2(n_511),
.B(n_499),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_524),
.A2(n_525),
.B1(n_518),
.B2(n_520),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_514),
.A2(n_492),
.B(n_496),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_523),
.B(n_515),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_529),
.B(n_519),
.C(n_489),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_530),
.Y(n_532)
);

AOI311xp33_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_527),
.A3(n_528),
.B(n_360),
.C(n_283),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_532),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_283),
.Y(n_535)
);


endmodule