module fake_netlist_1_8215_n_635 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_635);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_635;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g72 ( .A(n_57), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_60), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_41), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_37), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_68), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_11), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_15), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_40), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_64), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_49), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_12), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_55), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_71), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_8), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_50), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_25), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_16), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_31), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_11), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_33), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_26), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_51), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_48), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_52), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_9), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_27), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_3), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_36), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_19), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_46), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_14), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_17), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_54), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_56), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_30), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_42), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_100), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_100), .B(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_100), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_92), .Y(n_120) );
NAND2xp33_ASAP7_75t_R g121 ( .A(n_108), .B(n_34), .Y(n_121) );
NAND2x1p5_ASAP7_75t_L g122 ( .A(n_77), .B(n_29), .Y(n_122) );
NOR2xp33_ASAP7_75t_R g123 ( .A(n_98), .B(n_35), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_98), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_73), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_81), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_73), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_115), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_74), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_72), .Y(n_131) );
INVx5_ASAP7_75t_L g132 ( .A(n_92), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
NOR2xp67_ASAP7_75t_L g134 ( .A(n_95), .B(n_1), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_93), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_105), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_105), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_113), .B(n_28), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_113), .B(n_2), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_113), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_77), .B(n_2), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_114), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_74), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_84), .B(n_3), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_78), .B(n_4), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_75), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_99), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_75), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_76), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_76), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_99), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_79), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_79), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_78), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_103), .Y(n_156) );
NAND2xp33_ASAP7_75t_L g157 ( .A(n_80), .B(n_38), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_83), .B(n_4), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_137), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_138), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_126), .B(n_96), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_141), .B(n_116), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_132), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_131), .B(n_96), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_141), .A2(n_82), .B1(n_112), .B2(n_87), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_141), .A2(n_90), .B1(n_94), .B2(n_110), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
AOI22xp33_ASAP7_75t_SL g176 ( .A1(n_125), .A2(n_116), .B1(n_112), .B2(n_87), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
NAND2xp33_ASAP7_75t_SL g179 ( .A(n_123), .B(n_82), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_154), .B(n_102), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_136), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_141), .B(n_111), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_118), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_118), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_128), .B(n_97), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_147), .B(n_109), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_145), .B(n_109), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_145), .B(n_102), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_151), .B(n_104), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_135), .B(n_107), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_128), .B(n_107), .Y(n_200) );
NOR3xp33_ASAP7_75t_L g201 ( .A(n_144), .B(n_106), .C(n_104), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_138), .Y(n_202) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_130), .A2(n_88), .B(n_101), .Y(n_203) );
INVx8_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_140), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_138), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_130), .B(n_88), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_156), .B(n_101), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_140), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_132), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_152), .B(n_91), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_185), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_201), .B(n_145), .Y(n_217) );
BUFx10_ASAP7_75t_L g218 ( .A(n_208), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_185), .Y(n_219) );
BUFx12f_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_182), .B(n_164), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_164), .B(n_145), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_189), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
INVxp67_ASAP7_75t_SL g226 ( .A(n_186), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_164), .B(n_134), .Y(n_227) );
CKINVDCx14_ASAP7_75t_R g228 ( .A(n_179), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_167), .B(n_142), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_190), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_195), .B(n_153), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_193), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_186), .Y(n_235) );
NOR2xp33_ASAP7_75t_R g236 ( .A(n_204), .B(n_127), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_195), .B(n_152), .Y(n_237) );
OAI21xp33_ASAP7_75t_L g238 ( .A1(n_170), .A2(n_153), .B(n_118), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_205), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_163), .A2(n_158), .B(n_155), .C(n_150), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_184), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_165), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_195), .B(n_134), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_196), .B(n_143), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_196), .B(n_143), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_196), .B(n_143), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_194), .B(n_129), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_173), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_161), .B(n_122), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_196), .B(n_155), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_186), .B(n_150), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_194), .B(n_148), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_205), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_173), .A2(n_122), .B1(n_148), .B2(n_106), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_169), .B(n_122), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_209), .Y(n_256) );
NOR2xp33_ASAP7_75t_R g257 ( .A(n_204), .B(n_121), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_169), .B(n_132), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_169), .B(n_132), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_198), .B(n_139), .Y(n_260) );
BUFx6f_ASAP7_75t_SL g261 ( .A(n_209), .Y(n_261) );
NOR2xp33_ASAP7_75t_R g262 ( .A(n_204), .B(n_157), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_169), .B(n_132), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_165), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_171), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_198), .Y(n_266) );
INVx6_ASAP7_75t_L g267 ( .A(n_202), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_176), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_171), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_199), .B(n_117), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_212), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_172), .Y(n_272) );
BUFx5_ASAP7_75t_L g273 ( .A(n_206), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_187), .B(n_117), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_266), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_226), .A2(n_187), .B1(n_191), .B2(n_215), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_216), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_220), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_247), .B(n_192), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_220), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_240), .A2(n_187), .B(n_191), .C(n_207), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
INVx4_ASAP7_75t_L g284 ( .A(n_261), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_235), .A2(n_191), .B1(n_200), .B2(n_161), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_252), .Y(n_286) );
OR2x6_ASAP7_75t_L g287 ( .A(n_222), .B(n_204), .Y(n_287) );
OAI21x1_ASAP7_75t_SL g288 ( .A1(n_232), .A2(n_161), .B(n_211), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_221), .B(n_191), .Y(n_289) );
INVx5_ASAP7_75t_L g290 ( .A(n_267), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_227), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_219), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_261), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_217), .B(n_212), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_222), .A2(n_211), .B1(n_161), .B2(n_204), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_246), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_227), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_217), .A2(n_203), .B1(n_213), .B2(n_211), .Y(n_299) );
OAI21x1_ASAP7_75t_SL g300 ( .A1(n_237), .A2(n_211), .B(n_203), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_246), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_217), .B(n_213), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_267), .Y(n_303) );
OAI21xp33_ASAP7_75t_L g304 ( .A1(n_238), .A2(n_206), .B(n_166), .Y(n_304) );
OAI22xp33_ASAP7_75t_SL g305 ( .A1(n_268), .A2(n_85), .B1(n_86), .B2(n_89), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_274), .Y(n_306) );
INVx5_ASAP7_75t_L g307 ( .A(n_267), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_222), .A2(n_203), .B1(n_120), .B2(n_133), .Y(n_308) );
INVx3_ASAP7_75t_SL g309 ( .A(n_260), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g310 ( .A1(n_254), .A2(n_119), .B1(n_124), .B2(n_86), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_218), .B(n_188), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_251), .A2(n_197), .B1(n_210), .B2(n_202), .Y(n_312) );
INVx5_ASAP7_75t_L g313 ( .A(n_275), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_250), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_227), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_223), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_273), .B(n_210), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_255), .A2(n_210), .B(n_202), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_244), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_260), .A2(n_210), .B1(n_202), .B2(n_197), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_224), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_260), .B(n_197), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_249), .A2(n_210), .B(n_202), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_270), .B(n_166), .Y(n_324) );
BUFx8_ASAP7_75t_L g325 ( .A(n_243), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_236), .Y(n_326) );
BUFx12f_ASAP7_75t_L g327 ( .A(n_243), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_278), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_280), .A2(n_270), .B1(n_243), .B2(n_245), .Y(n_329) );
O2A1O1Ixp5_ASAP7_75t_SL g330 ( .A1(n_317), .A2(n_89), .B(n_91), .C(n_249), .Y(n_330) );
OA21x2_ASAP7_75t_L g331 ( .A1(n_300), .A2(n_282), .B(n_308), .Y(n_331) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_284), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_281), .B(n_270), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_281), .B(n_229), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_286), .B(n_248), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_306), .B(n_228), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_325), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_276), .A2(n_283), .B1(n_326), .B2(n_294), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_325), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_284), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_294), .B(n_236), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_325), .Y(n_342) );
INVx4_ASAP7_75t_SL g343 ( .A(n_287), .Y(n_343) );
CKINVDCx11_ASAP7_75t_R g344 ( .A(n_327), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_326), .Y(n_345) );
INVx6_ASAP7_75t_L g346 ( .A(n_327), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_291), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_314), .B(n_228), .Y(n_348) );
INVx4_ASAP7_75t_L g349 ( .A(n_287), .Y(n_349) );
AO31x2_ASAP7_75t_L g350 ( .A1(n_282), .A2(n_162), .A3(n_178), .B(n_159), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_313), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_287), .B(n_225), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_301), .B(n_230), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_311), .Y(n_354) );
INVx4_ASAP7_75t_SL g355 ( .A(n_309), .Y(n_355) );
INVx4_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_305), .A2(n_233), .B1(n_239), .B2(n_271), .C(n_253), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_278), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_293), .Y(n_359) );
CKINVDCx11_ASAP7_75t_R g360 ( .A(n_309), .Y(n_360) );
OAI222xp33_ASAP7_75t_L g361 ( .A1(n_310), .A2(n_234), .B1(n_256), .B2(n_259), .C1(n_258), .C2(n_263), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_361), .A2(n_299), .B(n_308), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_335), .B(n_279), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_338), .A2(n_289), .B1(n_319), .B2(n_302), .C(n_295), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_329), .A2(n_354), .B1(n_334), .B2(n_342), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_329), .A2(n_334), .B1(n_342), .B2(n_352), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_336), .A2(n_299), .B(n_315), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_328), .A2(n_359), .B1(n_358), .B2(n_313), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_328), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_343), .B(n_313), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g372 ( .A1(n_330), .A2(n_277), .B(n_285), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_352), .A2(n_316), .B1(n_293), .B2(n_321), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_352), .A2(n_321), .B1(n_316), .B2(n_297), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g375 ( .A1(n_357), .A2(n_304), .B(n_318), .C(n_292), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_334), .A2(n_298), .B1(n_322), .B2(n_218), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_333), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_356), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_337), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_349), .A2(n_322), .B1(n_297), .B2(n_279), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_331), .A2(n_323), .B(n_317), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_331), .B(n_348), .C(n_347), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_333), .A2(n_324), .B1(n_320), .B2(n_312), .C(n_296), .Y(n_384) );
AOI21xp33_ASAP7_75t_L g385 ( .A1(n_331), .A2(n_288), .B(n_322), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_353), .A2(n_210), .B(n_202), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_346), .A2(n_214), .B1(n_188), .B2(n_175), .C(n_177), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_349), .B(n_303), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_373), .A2(n_349), .B1(n_356), .B2(n_341), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_383), .B(n_351), .C(n_353), .Y(n_391) );
NAND2xp33_ASAP7_75t_R g392 ( .A(n_379), .B(n_341), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_370), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_370), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_362), .A2(n_353), .B(n_351), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_364), .B(n_351), .C(n_168), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_378), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_378), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_386), .Y(n_399) );
AOI33xp33_ASAP7_75t_L g400 ( .A1(n_365), .A2(n_340), .A3(n_180), .B1(n_174), .B2(n_175), .B3(n_177), .Y(n_400) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_374), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_363), .B(n_346), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_386), .B(n_350), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_371), .B(n_343), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_386), .B(n_350), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_389), .Y(n_407) );
OR2x6_ASAP7_75t_L g408 ( .A(n_371), .B(n_341), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_366), .A2(n_346), .B1(n_345), .B2(n_214), .C(n_174), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_377), .A2(n_345), .B1(n_332), .B2(n_343), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_389), .B(n_350), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_382), .B(n_350), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_367), .B(n_355), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_368), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_376), .B(n_355), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_369), .A2(n_181), .B1(n_183), .B2(n_257), .C(n_159), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_381), .A2(n_344), .B1(n_360), .B2(n_355), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_380), .Y(n_420) );
BUFx5_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_375), .B(n_360), .Y(n_422) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_396), .B(n_375), .Y(n_423) );
NAND2xp33_ASAP7_75t_L g424 ( .A(n_390), .B(n_344), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_410), .A2(n_388), .B1(n_372), .B2(n_387), .C(n_168), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_422), .A2(n_168), .B1(n_160), .B2(n_162), .C(n_178), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_404), .B(n_58), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_394), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_398), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_394), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_403), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_404), .B(n_59), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_411), .B(n_5), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_396), .B(n_332), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_411), .B(n_5), .Y(n_439) );
INVx5_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
AOI21xp33_ASAP7_75t_SL g441 ( .A1(n_392), .A2(n_408), .B(n_390), .Y(n_441) );
BUFx12f_ASAP7_75t_L g442 ( .A(n_420), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_406), .B(n_6), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_412), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_391), .B(n_168), .C(n_160), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_419), .A2(n_168), .B1(n_160), .B2(n_197), .C(n_307), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_393), .B(n_6), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_407), .B(n_7), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_407), .B(n_7), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_397), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_395), .A2(n_160), .B1(n_197), .B2(n_290), .C(n_307), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_399), .Y(n_455) );
OR2x6_ASAP7_75t_L g456 ( .A(n_395), .B(n_303), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_8), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_414), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_402), .B(n_265), .C(n_272), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_397), .B(n_9), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_399), .B(n_10), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_391), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_414), .B(n_10), .Y(n_465) );
NOR2x1p5_ASAP7_75t_L g466 ( .A(n_401), .B(n_12), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_405), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_414), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_437), .B(n_421), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_437), .B(n_418), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_424), .B(n_449), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_440), .B(n_408), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_439), .B(n_418), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_428), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_440), .B(n_408), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_439), .B(n_421), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_452), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_438), .A2(n_415), .B(n_413), .Y(n_479) );
AOI31xp33_ASAP7_75t_L g480 ( .A1(n_441), .A2(n_405), .A3(n_416), .B(n_408), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_443), .B(n_421), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_460), .B(n_409), .C(n_418), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_443), .B(n_415), .Y(n_483) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_466), .B(n_457), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_430), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_450), .B(n_414), .Y(n_486) );
NAND3xp33_ASAP7_75t_SL g487 ( .A(n_460), .B(n_400), .C(n_417), .Y(n_487) );
NAND2xp33_ASAP7_75t_L g488 ( .A(n_466), .B(n_421), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_450), .B(n_414), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_449), .B(n_421), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_442), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_440), .B(n_13), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_430), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_455), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_457), .B(n_421), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_432), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_442), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_429), .B(n_421), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_451), .B(n_421), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_457), .B(n_421), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_451), .B(n_15), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_433), .B(n_16), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_433), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_448), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_448), .B(n_18), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_442), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_436), .B(n_18), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_461), .B(n_19), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_432), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_461), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_436), .B(n_20), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_441), .B(n_20), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_453), .B(n_21), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_459), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_447), .B(n_21), .C(n_22), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_492), .Y(n_518) );
OAI32xp33_ASAP7_75t_L g519 ( .A1(n_508), .A2(n_434), .A3(n_467), .B1(n_447), .B2(n_465), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_502), .A2(n_464), .B1(n_465), .B2(n_463), .C(n_446), .Y(n_520) );
OAI31xp33_ASAP7_75t_L g521 ( .A1(n_514), .A2(n_453), .A3(n_467), .B(n_463), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g522 ( .A1(n_502), .A2(n_465), .B1(n_464), .B2(n_440), .C1(n_435), .C2(n_427), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_488), .A2(n_480), .B(n_517), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_477), .Y(n_524) );
OAI31xp33_ASAP7_75t_L g525 ( .A1(n_514), .A2(n_454), .A3(n_427), .B(n_435), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_478), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_511), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_482), .A2(n_440), .B1(n_427), .B2(n_435), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_507), .A2(n_444), .B1(n_446), .B2(n_458), .C(n_426), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_470), .B(n_444), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_517), .A2(n_445), .B(n_454), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_482), .A2(n_440), .B1(n_435), .B2(n_427), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_484), .B(n_468), .C(n_423), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_473), .B(n_444), .Y(n_534) );
AOI322xp5_ASAP7_75t_L g535 ( .A1(n_471), .A2(n_423), .A3(n_440), .B1(n_446), .B2(n_458), .C1(n_425), .C2(n_431), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_498), .B(n_22), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_471), .A2(n_458), .B1(n_425), .B2(n_468), .C1(n_431), .C2(n_459), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_511), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_510), .B(n_23), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_512), .B(n_23), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_506), .B(n_456), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_487), .B(n_445), .C(n_462), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_504), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_472), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_472), .B(n_462), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_485), .B(n_491), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_485), .B(n_456), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_494), .B(n_456), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_509), .A2(n_160), .B1(n_262), .B2(n_241), .C(n_231), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_513), .B(n_456), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_490), .A2(n_456), .B1(n_307), .B2(n_290), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_487), .A2(n_456), .B1(n_303), .B2(n_307), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_494), .A2(n_290), .B(n_303), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_479), .A2(n_290), .B1(n_241), .B2(n_272), .C(n_269), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_497), .B(n_39), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_491), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_497), .Y(n_559) );
OAI22xp33_ASAP7_75t_SL g560 ( .A1(n_503), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_526), .Y(n_563) );
XNOR2xp5_ASAP7_75t_L g564 ( .A(n_518), .B(n_475), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_523), .B(n_475), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_561), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_545), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_538), .Y(n_568) );
XNOR2xp5_ASAP7_75t_L g569 ( .A(n_528), .B(n_515), .Y(n_569) );
XOR2x2_ASAP7_75t_L g570 ( .A(n_536), .B(n_493), .Y(n_570) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_533), .B(n_483), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_532), .A2(n_469), .B1(n_476), .B2(n_481), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_547), .B(n_486), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_547), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_559), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_556), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_531), .A2(n_500), .B1(n_499), .B2(n_501), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_527), .B(n_489), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_525), .A2(n_496), .B(n_505), .C(n_516), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_544), .Y(n_580) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_539), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_530), .B(n_516), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_534), .B(n_505), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_545), .B(n_47), .Y(n_584) );
BUFx2_ASAP7_75t_L g585 ( .A(n_546), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_558), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_542), .B(n_53), .Y(n_587) );
INVx3_ASAP7_75t_SL g588 ( .A(n_546), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_549), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_548), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_579), .A2(n_535), .B(n_521), .Y(n_591) );
OAI321xp33_ASAP7_75t_L g592 ( .A1(n_565), .A2(n_553), .A3(n_520), .B1(n_541), .B2(n_552), .C(n_551), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_577), .A2(n_540), .B1(n_519), .B2(n_543), .C(n_529), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_579), .A2(n_560), .B(n_555), .C(n_537), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_574), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_588), .B(n_522), .Y(n_596) );
NAND2x1_ASAP7_75t_L g597 ( .A(n_585), .B(n_552), .Y(n_597) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_584), .B(n_554), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_570), .B(n_557), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_587), .B(n_550), .C(n_264), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_569), .A2(n_273), .B1(n_242), .B2(n_62), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_590), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_581), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_566), .A2(n_273), .B1(n_242), .B2(n_65), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_576), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g606 ( .A1(n_570), .A2(n_61), .B1(n_63), .B2(n_66), .C1(n_69), .C2(n_273), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_571), .A2(n_273), .B(n_578), .Y(n_607) );
INVxp33_ASAP7_75t_L g608 ( .A(n_597), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_599), .B(n_564), .Y(n_609) );
AO22x2_ASAP7_75t_L g610 ( .A1(n_603), .A2(n_567), .B1(n_575), .B2(n_562), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_595), .B(n_577), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_591), .A2(n_589), .B1(n_578), .B2(n_563), .C(n_580), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_591), .A2(n_573), .B1(n_583), .B2(n_572), .Y(n_613) );
NOR2xp33_ASAP7_75t_R g614 ( .A(n_596), .B(n_568), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_593), .A2(n_606), .B1(n_601), .B2(n_607), .Y(n_615) );
NAND3xp33_ASAP7_75t_SL g616 ( .A(n_606), .B(n_586), .C(n_576), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g617 ( .A(n_594), .B(n_582), .C(n_604), .D(n_600), .Y(n_617) );
OAI211xp5_ASAP7_75t_SL g618 ( .A1(n_602), .A2(n_582), .B(n_592), .C(n_605), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g619 ( .A1(n_598), .A2(n_508), .B1(n_597), .B2(n_599), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_598), .B(n_596), .Y(n_620) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_599), .B(n_570), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_597), .A2(n_565), .B(n_591), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_611), .B(n_616), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_620), .B(n_608), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_612), .B(n_613), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_621), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_626), .B(n_618), .C(n_619), .Y(n_627) );
XNOR2xp5_ASAP7_75t_L g628 ( .A(n_626), .B(n_615), .Y(n_628) );
OR5x1_ASAP7_75t_L g629 ( .A(n_623), .B(n_617), .C(n_622), .D(n_610), .E(n_614), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_628), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_629), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_630), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_631), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_632), .B(n_631), .C(n_627), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_634), .A2(n_633), .B1(n_625), .B2(n_624), .C(n_609), .Y(n_635) );
endmodule