module fake_ariane_3356_n_309 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_309);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_309;

wire n_295;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_180;
wire n_124;
wire n_119;
wire n_307;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_183;
wire n_299;
wire n_133;
wire n_66;
wire n_205;
wire n_71;
wire n_109;
wire n_245;
wire n_96;
wire n_283;
wire n_187;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_189;
wire n_72;
wire n_286;
wire n_57;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_214;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_52;
wire n_73;
wire n_77;
wire n_87;
wire n_279;
wire n_207;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_59;
wire n_239;
wire n_272;
wire n_54;
wire n_167;
wire n_90;
wire n_153;
wire n_269;
wire n_75;
wire n_158;
wire n_69;
wire n_259;
wire n_95;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_115;
wire n_267;
wire n_291;
wire n_62;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_79;
wire n_271;
wire n_247;
wire n_91;
wire n_240;
wire n_128;
wire n_224;
wire n_82;
wire n_222;
wire n_256;
wire n_227;
wire n_188;
wire n_129;
wire n_126;
wire n_282;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_276;
wire n_93;
wire n_108;
wire n_303;
wire n_168;
wire n_81;
wire n_206;
wire n_238;
wire n_136;
wire n_192;
wire n_300;
wire n_163;
wire n_88;
wire n_141;
wire n_104;
wire n_273;
wire n_305;
wire n_233;
wire n_56;
wire n_60;
wire n_221;
wire n_86;
wire n_89;
wire n_149;
wire n_237;
wire n_175;
wire n_74;
wire n_181;
wire n_53;
wire n_260;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_84;
wire n_199;
wire n_107;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_70;
wire n_287;
wire n_302;
wire n_94;
wire n_284;
wire n_249;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_61;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_55;
wire n_231;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_68;
wire n_78;
wire n_63;
wire n_99;
wire n_216;
wire n_223;
wire n_83;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_67;
wire n_306;
wire n_92;
wire n_203;
wire n_150;
wire n_98;
wire n_113;
wire n_114;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_76;
wire n_246;
wire n_159;
wire n_105;
wire n_131;
wire n_263;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_101;
wire n_243;
wire n_134;
wire n_185;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_258;
wire n_118;
wire n_121;
wire n_241;
wire n_191;
wire n_80;
wire n_211;
wire n_97;
wire n_251;
wire n_116;
wire n_155;
wire n_127;

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_51),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_3),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_3),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_71),
.B1(n_73),
.B2(n_83),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_63),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_58),
.B1(n_73),
.B2(n_55),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_68),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_55),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_7),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_85),
.B(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_11),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_88),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_112),
.Y(n_140)
);

AND3x1_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_84),
.C(n_89),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_103),
.Y(n_146)
);

NAND2x1p5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

AND2x6_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_92),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_84),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_110),
.B1(n_105),
.B2(n_104),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_104),
.Y(n_156)
);

OR2x6_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_110),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_125),
.B1(n_118),
.B2(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_125),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_129),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_134),
.B(n_133),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_135),
.B(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_143),
.Y(n_168)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_135),
.B(n_121),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_12),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_144),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_104),
.B(n_98),
.C(n_86),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_155),
.B(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_179),
.B1(n_176),
.B2(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_156),
.B(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_152),
.B(n_144),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_144),
.B(n_17),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_177),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_149),
.B1(n_104),
.B2(n_98),
.Y(n_197)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_13),
.B(n_22),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_158),
.B1(n_172),
.B2(n_173),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_187),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_170),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_188),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_158),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

AOI221xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_167),
.B1(n_161),
.B2(n_163),
.C(n_172),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_172),
.B1(n_175),
.B2(n_174),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_177),
.Y(n_216)
);

AO21x2_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_194),
.B(n_181),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_186),
.Y(n_223)
);

OAI31xp33_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_191),
.A3(n_193),
.B(n_187),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_211),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_232),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_243),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_227),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_223),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_242),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_217),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_211),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_221),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_221),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_215),
.B1(n_187),
.B2(n_193),
.Y(n_264)
);

AND2x4_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_193),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_245),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_198),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_217),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_224),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_254),
.Y(n_276)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_261),
.B(n_257),
.C(n_259),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_253),
.Y(n_278)
);

AOI211xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_264),
.B(n_259),
.C(n_262),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_264),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_277),
.B(n_281),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_273),
.C(n_270),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_271),
.B(n_284),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

AOI211xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_284),
.B(n_275),
.C(n_276),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_268),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_274),
.B1(n_266),
.B2(n_263),
.Y(n_292)
);

NAND2x1_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_190),
.Y(n_293)
);

OAI321xp33_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_192),
.A3(n_98),
.B1(n_181),
.B2(n_198),
.C(n_30),
.Y(n_294)
);

OR4x2_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_190),
.C(n_183),
.D(n_194),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

AOI211xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_98),
.B(n_193),
.C(n_26),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_293),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_190),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_298),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_295),
.B1(n_294),
.B2(n_190),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_183),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_183),
.Y(n_304)
);

AOI221xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_299),
.B1(n_302),
.B2(n_300),
.C(n_301),
.Y(n_305)
);

AO221x1_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_181),
.B1(n_25),
.B2(n_27),
.C(n_31),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

AOI221xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_305),
.B1(n_307),
.B2(n_41),
.C(n_44),
.Y(n_309)
);


endmodule