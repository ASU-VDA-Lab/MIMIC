module fake_netlist_5_168_n_4417 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_4417);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_4417;

wire n_924;
wire n_1263;
wire n_3304;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_977;
wire n_611;
wire n_2756;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_3241;
wire n_4129;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_667;
wire n_2955;
wire n_2899;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4138;
wire n_880;
wire n_4127;
wire n_3086;
wire n_3297;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_4217;
wire n_4395;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_956;
wire n_564;
wire n_4240;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_551;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_671;
wire n_4238;
wire n_819;
wire n_1451;
wire n_1022;
wire n_4038;
wire n_2302;
wire n_915;
wire n_4109;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_4412;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3599;
wire n_3571;
wire n_3785;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_516;
wire n_2244;
wire n_933;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_4013;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_1860;
wire n_2543;
wire n_4155;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_556;
wire n_3036;
wire n_2482;
wire n_3695;
wire n_3891;
wire n_4145;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3180;
wire n_3010;
wire n_3379;
wire n_3832;
wire n_4374;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_659;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_579;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_4315;
wire n_546;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_4311;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_4358;
wire n_3490;
wire n_3656;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_4369;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_4394;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_4350;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_3156;
wire n_550;
wire n_696;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_3876;
wire n_926;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_4135;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_1547;
wire n_1070;
wire n_777;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_521;
wire n_3744;
wire n_845;
wire n_663;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_673;
wire n_837;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_4255;
wire n_1587;
wire n_1473;
wire n_680;
wire n_2682;
wire n_553;
wire n_901;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_813;
wire n_4258;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_2506;
wire n_675;
wire n_2699;
wire n_4064;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3550;
wire n_637;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_3262;
wire n_1075;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3986;
wire n_4376;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_571;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3593;
wire n_3193;
wire n_3837;
wire n_3885;
wire n_1971;
wire n_1599;
wire n_3936;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2700;
wire n_2644;
wire n_4310;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_907;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_3915;
wire n_4414;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_4114;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3349;
wire n_3025;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_736;
wire n_892;
wire n_4385;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_593;
wire n_3487;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_3470;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_4327;
wire n_4405;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_953;
wire n_1014;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_4375;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_3781;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_4353;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_884;
wire n_3328;
wire n_944;
wire n_4130;
wire n_4234;
wire n_1754;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2674;
wire n_2606;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4161;
wire n_647;
wire n_3433;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_3392;
wire n_857;
wire n_832;
wire n_2305;
wire n_3430;
wire n_3975;
wire n_1072;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_561;
wire n_1319;
wire n_2379;
wire n_3447;
wire n_3331;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_4148;
wire n_4151;
wire n_1883;
wire n_1906;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_4415;
wire n_1387;
wire n_3649;
wire n_3528;
wire n_2262;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_4373;
wire n_1532;
wire n_4252;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3625;
wire n_3257;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_4331;
wire n_4160;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_3989;
wire n_2837;
wire n_847;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_558;
wire n_3655;
wire n_2808;
wire n_1276;
wire n_702;
wire n_3009;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_728;
wire n_4388;
wire n_2930;
wire n_1162;
wire n_1538;
wire n_4206;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_809;
wire n_3923;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_868;
wire n_2454;
wire n_4371;
wire n_639;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_2009;
wire n_1888;
wire n_759;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_3819;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_747;
wire n_2064;
wire n_784;
wire n_3978;
wire n_4325;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_4372;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_3747;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_3833;
wire n_865;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_678;
wire n_2671;
wire n_697;
wire n_4262;
wire n_4184;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_776;
wire n_2022;
wire n_1798;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_2592;
wire n_3416;
wire n_4379;
wire n_525;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_4340;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_4397;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_744;
wire n_629;
wire n_590;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_3317;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3220;
wire n_4391;
wire n_949;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_3855;
wire n_946;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_3452;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_3113;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_3205;
wire n_4156;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_4360;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_3866;
wire n_4404;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_524;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_4324;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_906;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4356;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_724;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_959;
wire n_2459;
wire n_3031;
wire n_4154;
wire n_535;
wire n_3396;
wire n_3701;
wire n_940;
wire n_4386;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_514;
wire n_1079;
wire n_2339;
wire n_2473;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_1045;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_4279;
wire n_4396;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_3820;
wire n_636;
wire n_4367;
wire n_3741;
wire n_660;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_2029;
wire n_750;
wire n_995;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_4232;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_4413;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_4387;
wire n_662;
wire n_2312;
wire n_3990;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_4365;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_974;
wire n_4152;
wire n_727;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_957;
wire n_3787;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_4392;
wire n_3149;
wire n_613;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_4285;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_3960;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_761;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3905;
wire n_4329;
wire n_1006;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_4271;
wire n_1486;
wire n_582;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_512;
wire n_1591;
wire n_2033;
wire n_4071;
wire n_4330;
wire n_4341;
wire n_4257;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_4361;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3838;
wire n_3077;
wire n_3929;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_765;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_3984;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_630;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_4326;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4305;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_860;
wire n_3229;
wire n_4213;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_628;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_4313;
wire n_970;
wire n_4037;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_513;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_560;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_602;
wire n_3525;
wire n_574;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_623;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_824;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4339;
wire n_4041;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_3751;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_589;
wire n_3961;
wire n_1630;
wire n_2122;
wire n_716;
wire n_2512;
wire n_3589;
wire n_4102;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_701;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_531;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2969;
wire n_2864;
wire n_3941;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_950;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_968;
wire n_912;
wire n_3548;
wire n_4348;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_4355;
wire n_3494;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_515;
wire n_2333;
wire n_3953;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_683;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_841;
wire n_1050;
wire n_1954;
wire n_802;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_4104;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_4377;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_3991;
wire n_3962;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_762;
wire n_1283;
wire n_1644;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_4384;
wire n_690;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_3816;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_4286;
wire n_3864;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3299;
wire n_3041;
wire n_3274;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_4362;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_3921;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_4400;
wire n_943;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_992;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_543;
wire n_842;
wire n_3734;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_4402;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_918;
wire n_3529;
wire n_3854;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_2533;
wire n_2364;
wire n_4338;
wire n_540;
wire n_3492;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_1511;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_3689;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_4416;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2751;
wire n_2707;
wire n_2793;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_1446;
wire n_2285;
wire n_4406;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_669;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_3869;
wire n_4307;
wire n_1149;
wire n_2618;
wire n_4359;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_555;
wire n_1848;
wire n_1928;
wire n_783;
wire n_2126;
wire n_4117;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_661;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_849;
wire n_2795;
wire n_4091;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_510;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_830;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3460;
wire n_3409;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_801;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_4247;
wire n_2638;
wire n_866;
wire n_1401;
wire n_969;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_3759;
wire n_1338;
wire n_577;
wire n_4409;
wire n_4411;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_4336;
wire n_3933;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_836;
wire n_990;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4253;
wire n_4290;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_711;
wire n_3061;
wire n_4398;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_3356;
wire n_3324;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_4304;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_601;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4115;
wire n_726;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1453;
wire n_2217;
wire n_1731;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_2745;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_774;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_3967;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_665;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_3839;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3972;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_3358;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_2224;
wire n_732;
wire n_1533;
wire n_791;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_2484;
wire n_808;
wire n_4111;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_766;
wire n_3928;
wire n_541;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_3534;
wire n_715;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_536;
wire n_3438;
wire n_4098;
wire n_872;
wire n_2012;
wire n_594;
wire n_3792;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_4269;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_4150;
wire n_827;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_676;
wire n_2103;
wire n_653;
wire n_3968;
wire n_2160;
wire n_642;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_4380;
wire n_980;
wire n_1115;
wire n_698;
wire n_703;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_998;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_823;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_725;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3172;
wire n_3292;
wire n_2773;
wire n_3139;
wire n_3239;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_4220;
wire n_4251;
wire n_1683;
wire n_1817;
wire n_1944;
wire n_909;
wire n_1497;
wire n_1530;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_4351;
wire n_2819;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_4368;
wire n_1718;
wire n_737;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_4136;
wire n_986;
wire n_2315;
wire n_509;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_4393;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_867;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_548;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_518;
wire n_505;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_760;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_4382;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_4178;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_751;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_704;
wire n_787;
wire n_4399;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_4401;
wire n_3904;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_3364;
wire n_1287;
wire n_4363;
wire n_1262;
wire n_2691;
wire n_930;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_622;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_682;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_4015;
wire n_591;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_631;
wire n_3627;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_839;
wire n_3551;
wire n_3903;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3859;
wire n_3722;
wire n_3865;
wire n_4171;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_598;
wire n_685;
wire n_608;
wire n_1367;
wire n_928;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_517;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2702;
wire n_2570;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_3115;
wire n_4287;
wire n_3509;
wire n_3352;
wire n_4390;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_3251;
wire n_1061;
wire n_1910;
wire n_3955;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2050;
wire n_2809;
wire n_4270;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_722;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1028;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_781;
wire n_2940;
wire n_542;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_595;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_4231;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3322;
wire n_3232;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2505;
wire n_2427;
wire n_2438;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_4061;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_3250;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_3125;
wire n_3114;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_648;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_4407;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_2823;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_4389;
wire n_3930;
wire n_730;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_695;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_805;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4319;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_657;
wire n_4320;
wire n_644;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_4245;
wire n_4288;
wire n_4364;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_4378;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1181;
wire n_1505;
wire n_4216;
wire n_4222;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_3225;
wire n_1558;
wire n_4241;
wire n_807;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_835;
wire n_666;
wire n_3319;
wire n_3594;
wire n_1433;
wire n_4309;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2920;
wire n_2689;
wire n_3259;
wire n_4265;
wire n_1004;
wire n_1186;
wire n_2614;
wire n_1032;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_4366;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

INVx1_ASAP7_75t_SL g503 ( 
.A(n_11),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_162),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_0),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_493),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_451),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_282),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_25),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_365),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_60),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_14),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_248),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_273),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_28),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_218),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_64),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_180),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_173),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_209),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_7),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_39),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_223),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_438),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_357),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_66),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_408),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_28),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_367),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_501),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_37),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_495),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_333),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_369),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_250),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_75),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_289),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_0),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_86),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_386),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_328),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_446),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_466),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_165),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_393),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_254),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_308),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_104),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_29),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_59),
.Y(n_552)
);

BUFx5_ASAP7_75t_L g553 ( 
.A(n_455),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_320),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_479),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_487),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_331),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_64),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_70),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_302),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_502),
.Y(n_561)
);

CKINVDCx16_ASAP7_75t_R g562 ( 
.A(n_236),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_365),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_245),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_152),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_40),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_465),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_293),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_207),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_412),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_404),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_100),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_29),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_191),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_23),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_88),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_204),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_330),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_58),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_474),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_79),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_198),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_106),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_428),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_227),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_57),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_197),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_264),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_489),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_39),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_323),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_239),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_176),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_70),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_145),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_5),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_317),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_439),
.Y(n_598)
);

CKINVDCx14_ASAP7_75t_R g599 ( 
.A(n_320),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_4),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_14),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_294),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_114),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_325),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_311),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_361),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_335),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_381),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_326),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_307),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_396),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_401),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_219),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_107),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_417),
.Y(n_615)
);

BUFx5_ASAP7_75t_L g616 ( 
.A(n_34),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_338),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_66),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_218),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_15),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_257),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_497),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_375),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_397),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_91),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_76),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_238),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_154),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_171),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_77),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_221),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_122),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_144),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_352),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_21),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_7),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_89),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_275),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_51),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_147),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_112),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_470),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_340),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_419),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_51),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_358),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_348),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_395),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_109),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_486),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_195),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_327),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_24),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_358),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_431),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_299),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_118),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_291),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_206),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_23),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_145),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_161),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_122),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_307),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_32),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_310),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_196),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_119),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_350),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_459),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_378),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_360),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_154),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_71),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_106),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_289),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_125),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_357),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_429),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_249),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_140),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_481),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_337),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_268),
.Y(n_684)
);

CKINVDCx14_ASAP7_75t_R g685 ( 
.A(n_322),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_380),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_104),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_98),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_113),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_420),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_209),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_338),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_424),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_137),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_298),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_212),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_468),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_173),
.Y(n_698)
);

CKINVDCx16_ASAP7_75t_R g699 ( 
.A(n_68),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_161),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_257),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_361),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_251),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_204),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_285),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_198),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_112),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_200),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_388),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_488),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_202),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_414),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_500),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_275),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_11),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_71),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_272),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_208),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_247),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_98),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_384),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_34),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_247),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_239),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_230),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_284),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_385),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_402),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_343),
.Y(n_729)
);

BUFx8_ASAP7_75t_SL g730 ( 
.A(n_187),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_391),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_194),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_321),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_233),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_339),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_329),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_242),
.Y(n_737)
);

CKINVDCx14_ASAP7_75t_R g738 ( 
.A(n_93),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_53),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_149),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_196),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_192),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_114),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_283),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_186),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_249),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_47),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_236),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_5),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_336),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_406),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_480),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_110),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_96),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_252),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_115),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_32),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_41),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_175),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_268),
.Y(n_760)
);

CKINVDCx16_ASAP7_75t_R g761 ( 
.A(n_158),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_379),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_356),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_228),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_272),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_136),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_108),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_360),
.Y(n_768)
);

BUFx10_ASAP7_75t_L g769 ( 
.A(n_405),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_83),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_25),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_387),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_344),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_169),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_418),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_376),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_180),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_171),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_4),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_146),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_142),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_67),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_208),
.Y(n_783)
);

BUFx10_ASAP7_75t_L g784 ( 
.A(n_471),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_227),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_118),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_24),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_162),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_484),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_43),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_85),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_288),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_62),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_62),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_354),
.Y(n_795)
);

CKINVDCx14_ASAP7_75t_R g796 ( 
.A(n_241),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_38),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_276),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_72),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_99),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_167),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_273),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_462),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_373),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_75),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_306),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_183),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_223),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_22),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_153),
.Y(n_810)
);

CKINVDCx14_ASAP7_75t_R g811 ( 
.A(n_143),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_292),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_163),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_46),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_237),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_342),
.Y(n_816)
);

CKINVDCx16_ASAP7_75t_R g817 ( 
.A(n_504),
.Y(n_817)
);

INVxp33_ASAP7_75t_SL g818 ( 
.A(n_627),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_616),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_616),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_730),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_556),
.Y(n_822)
);

INVxp33_ASAP7_75t_SL g823 ( 
.A(n_724),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_616),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_616),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_616),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_507),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_529),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_616),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_616),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_523),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_525),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_566),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_616),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_598),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_622),
.Y(n_836)
);

INVxp33_ASAP7_75t_SL g837 ( 
.A(n_745),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_616),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_679),
.Y(n_839)
);

INVxp33_ASAP7_75t_SL g840 ( 
.A(n_792),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_531),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_531),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_622),
.B(n_1),
.Y(n_843)
);

CKINVDCx14_ASAP7_75t_R g844 ( 
.A(n_599),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_534),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_531),
.Y(n_846)
);

INVxp33_ASAP7_75t_SL g847 ( 
.A(n_566),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_505),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_505),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_531),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_794),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_542),
.Y(n_852)
);

CKINVDCx14_ASAP7_75t_R g853 ( 
.A(n_685),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_522),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_531),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_531),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_533),
.Y(n_857)
);

CKINVDCx16_ASAP7_75t_R g858 ( 
.A(n_504),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_533),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_533),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_533),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_533),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_524),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_533),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_585),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_585),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_544),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_585),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_511),
.Y(n_869)
);

INVxp33_ASAP7_75t_L g870 ( 
.A(n_524),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_585),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_585),
.Y(n_872)
);

CKINVDCx16_ASAP7_75t_R g873 ( 
.A(n_511),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_547),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_794),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_585),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_629),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_629),
.Y(n_878)
);

CKINVDCx16_ASAP7_75t_R g879 ( 
.A(n_554),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_629),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_629),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_589),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_608),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_794),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_528),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_629),
.Y(n_886)
);

INVxp33_ASAP7_75t_L g887 ( 
.A(n_526),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_629),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_656),
.Y(n_889)
);

INVxp67_ASAP7_75t_SL g890 ( 
.A(n_794),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_656),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_656),
.Y(n_892)
);

CKINVDCx16_ASAP7_75t_R g893 ( 
.A(n_554),
.Y(n_893)
);

INVxp33_ASAP7_75t_SL g894 ( 
.A(n_508),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_656),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_656),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_656),
.Y(n_897)
);

CKINVDCx16_ASAP7_75t_R g898 ( 
.A(n_562),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_733),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_733),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_721),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_526),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_562),
.Y(n_903)
);

INVx4_ASAP7_75t_R g904 ( 
.A(n_529),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_733),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_789),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_733),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_733),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_733),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_788),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_788),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_788),
.Y(n_912)
);

INVxp67_ASAP7_75t_SL g913 ( 
.A(n_529),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_788),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_611),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_738),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_788),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_788),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_699),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_510),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_615),
.Y(n_921)
);

INVxp33_ASAP7_75t_L g922 ( 
.A(n_535),
.Y(n_922)
);

BUFx2_ASAP7_75t_SL g923 ( 
.A(n_509),
.Y(n_923)
);

INVxp33_ASAP7_75t_SL g924 ( 
.A(n_512),
.Y(n_924)
);

INVxp33_ASAP7_75t_SL g925 ( 
.A(n_513),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_510),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_520),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_520),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_623),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_535),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_624),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_553),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_691),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_796),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_626),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_691),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_811),
.Y(n_937)
);

INVxp33_ASAP7_75t_SL g938 ( 
.A(n_514),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_644),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_714),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_648),
.Y(n_941)
);

INVxp33_ASAP7_75t_SL g942 ( 
.A(n_515),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_714),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_726),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_650),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_626),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_682),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_726),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_626),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_758),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_758),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_773),
.Y(n_952)
);

INVxp33_ASAP7_75t_L g953 ( 
.A(n_541),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_773),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_766),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_655),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_686),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_766),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_766),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_553),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_806),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_806),
.Y(n_962)
);

INVxp33_ASAP7_75t_SL g963 ( 
.A(n_516),
.Y(n_963)
);

INVxp33_ASAP7_75t_SL g964 ( 
.A(n_517),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_806),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_699),
.Y(n_966)
);

INVxp33_ASAP7_75t_SL g967 ( 
.A(n_518),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_553),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_541),
.Y(n_969)
);

INVxp33_ASAP7_75t_L g970 ( 
.A(n_548),
.Y(n_970)
);

OAI22x1_ASAP7_75t_SL g971 ( 
.A1(n_847),
.A2(n_552),
.B1(n_593),
.B2(n_576),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_828),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_897),
.Y(n_973)
);

OAI22x1_ASAP7_75t_L g974 ( 
.A1(n_833),
.A2(n_509),
.B1(n_586),
.B2(n_573),
.Y(n_974)
);

OA21x2_ASAP7_75t_L g975 ( 
.A1(n_841),
.A2(n_545),
.B(n_528),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_897),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_891),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_891),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_897),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_894),
.B(n_545),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_875),
.B(n_506),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_828),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_895),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_895),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_896),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_841),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_896),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_818),
.A2(n_761),
.B1(n_617),
.B2(n_674),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_842),
.Y(n_989)
);

XNOR2x2_ASAP7_75t_L g990 ( 
.A(n_854),
.B(n_503),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_899),
.Y(n_991)
);

OAI22x1_ASAP7_75t_R g992 ( 
.A1(n_822),
.A2(n_675),
.B1(n_678),
.B2(n_604),
.Y(n_992)
);

OA21x2_ASAP7_75t_L g993 ( 
.A1(n_842),
.A2(n_561),
.B(n_555),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_899),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_910),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_910),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_884),
.B(n_506),
.Y(n_997)
);

AND2x6_ASAP7_75t_L g998 ( 
.A(n_819),
.B(n_532),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_846),
.Y(n_999)
);

OAI22x1_ASAP7_75t_L g1000 ( 
.A1(n_843),
.A2(n_586),
.B1(n_764),
.B2(n_573),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_827),
.B(n_642),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_846),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_850),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_850),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_823),
.A2(n_761),
.B1(n_840),
.B2(n_837),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_955),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_L g1007 ( 
.A(n_855),
.B(n_642),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_890),
.B(n_803),
.Y(n_1008)
);

CKINVDCx6p67_ASAP7_75t_R g1009 ( 
.A(n_916),
.Y(n_1009)
);

BUFx8_ASAP7_75t_L g1010 ( 
.A(n_949),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_851),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_855),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_955),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_851),
.B(n_885),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_935),
.B(n_590),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_946),
.B(n_590),
.Y(n_1016)
);

CKINVDCx8_ASAP7_75t_R g1017 ( 
.A(n_817),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_913),
.B(n_621),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_819),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_924),
.B(n_555),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_856),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_856),
.A2(n_570),
.B(n_561),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_857),
.Y(n_1023)
);

INVx6_ASAP7_75t_L g1024 ( 
.A(n_947),
.Y(n_1024)
);

BUFx8_ASAP7_75t_SL g1025 ( 
.A(n_821),
.Y(n_1025)
);

BUFx8_ASAP7_75t_SL g1026 ( 
.A(n_934),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_857),
.Y(n_1027)
);

OAI22x1_ASAP7_75t_SL g1028 ( 
.A1(n_835),
.A2(n_722),
.B1(n_729),
.B2(n_708),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_859),
.B(n_803),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_859),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_831),
.B(n_690),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_860),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_860),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_858),
.B(n_682),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_820),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_861),
.B(n_570),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_869),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_958),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_932),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_832),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_958),
.B(n_621),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_839),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_861),
.B(n_571),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_932),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_862),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_862),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_959),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_947),
.Y(n_1048)
);

BUFx8_ASAP7_75t_L g1049 ( 
.A(n_949),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_864),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_864),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_960),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_820),
.Y(n_1054)
);

INVx6_ASAP7_75t_L g1055 ( 
.A(n_904),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_865),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_959),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_845),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_903),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_866),
.A2(n_580),
.B(n_571),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_844),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_852),
.B(n_693),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_901),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_866),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_868),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_868),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_871),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_871),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_872),
.Y(n_1069)
);

BUFx8_ASAP7_75t_L g1070 ( 
.A(n_853),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_966),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_872),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_876),
.A2(n_584),
.B(n_580),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_867),
.B(n_710),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_876),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_877),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_874),
.B(n_882),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_883),
.B(n_713),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_877),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_878),
.Y(n_1080)
);

AND2x2_ASAP7_75t_SL g1081 ( 
.A(n_873),
.B(n_532),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_878),
.B(n_584),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_880),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_906),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_937),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_879),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_923),
.B(n_893),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_880),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_881),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_960),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_898),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_881),
.B(n_670),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_886),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_886),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_961),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_915),
.B(n_921),
.Y(n_1096)
);

AOI22x1_ASAP7_75t_SL g1097 ( 
.A1(n_836),
.A2(n_759),
.B1(n_779),
.B2(n_748),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_1081),
.B(n_929),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1026),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_984),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1042),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_976),
.A2(n_825),
.B(n_824),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1006),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_1063),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_1087),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1006),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1019),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1006),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_1039),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1084),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1009),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_984),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1013),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1018),
.B(n_923),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1009),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1017),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_991),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_R g1118 ( 
.A(n_1040),
.B(n_931),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1013),
.Y(n_1119)
);

AND2x6_ASAP7_75t_L g1120 ( 
.A(n_981),
.B(n_532),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_991),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1013),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1001),
.B(n_939),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_981),
.B(n_941),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_983),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_1058),
.B(n_945),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1087),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1037),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1070),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1038),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1038),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_981),
.B(n_956),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1019),
.A2(n_825),
.B(n_824),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1070),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_1017),
.B(n_957),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1039),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1070),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1070),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1038),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1047),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_978),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1047),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1047),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1010),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1086),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_972),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1091),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1010),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1010),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_983),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1057),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_978),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1010),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1049),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1049),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_972),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1057),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_983),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1057),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_981),
.B(n_925),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_994),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1049),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1019),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_994),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_997),
.B(n_938),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1049),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1019),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1035),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_978),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_997),
.B(n_942),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1035),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1061),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1081),
.B(n_963),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_994),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1061),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1031),
.B(n_964),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_978),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1025),
.Y(n_1178)
);

XOR2xp5_ASAP7_75t_L g1179 ( 
.A(n_1028),
.B(n_919),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_996),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_1085),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1018),
.B(n_961),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_972),
.B(n_962),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1085),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_978),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_982),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_997),
.B(n_967),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_978),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1035),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_996),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1035),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1028),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_976),
.A2(n_829),
.B(n_826),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1054),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_996),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1003),
.Y(n_1196)
);

INVx6_ASAP7_75t_L g1197 ( 
.A(n_973),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_982),
.B(n_962),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1054),
.Y(n_1199)
);

AND2x6_ASAP7_75t_L g1200 ( 
.A(n_997),
.B(n_532),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_982),
.B(n_965),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1081),
.A2(n_618),
.B1(n_645),
.B2(n_596),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1062),
.B(n_970),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1003),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1059),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1074),
.B(n_849),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_971),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1027),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_971),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_987),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1015),
.B(n_965),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1008),
.B(n_888),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1054),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1027),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_1071),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_992),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1054),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1077),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1050),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_990),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1078),
.B(n_870),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1041),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1048),
.B(n_682),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_990),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1015),
.B(n_920),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1050),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1039),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1016),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1097),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_980),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1095),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1048),
.B(n_682),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1008),
.B(n_1020),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1039),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1052),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1095),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1097),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1016),
.B(n_920),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1052),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1014),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1096),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1056),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1014),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_992),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1014),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1024),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1024),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1024),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1024),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1014),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1056),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_988),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_988),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_979),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1008),
.B(n_670),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1002),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_979),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1005),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1005),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1034),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1055),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1044),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_986),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1008),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_986),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_987),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1002),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_989),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1002),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1041),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1044),
.B(n_888),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_989),
.A2(n_1004),
.B(n_999),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1055),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1044),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1044),
.B(n_889),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1055),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1055),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_999),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_975),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1000),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1004),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1000),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1012),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1033),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1036),
.B(n_926),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1090),
.B(n_953),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1036),
.B(n_926),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1012),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_975),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_974),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_SL g1291 ( 
.A(n_974),
.B(n_764),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1023),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1036),
.Y(n_1293)
);

BUFx8_ASAP7_75t_L g1294 ( 
.A(n_1036),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1023),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_987),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1043),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_987),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1030),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1033),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1090),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1043),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1030),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_987),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1033),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_987),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1065),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1043),
.B(n_927),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1065),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1066),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1046),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1043),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1090),
.B(n_889),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1082),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1082),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1046),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1066),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1046),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1079),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1082),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1082),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1064),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1079),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1090),
.B(n_892),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1080),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1114),
.B(n_1203),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1109),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1206),
.B(n_1092),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1264),
.A2(n_993),
.B1(n_1022),
.B2(n_975),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1272),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1221),
.B(n_1092),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1272),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1272),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1272),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1107),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1114),
.B(n_727),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1107),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1163),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1102),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1264),
.A2(n_1289),
.B1(n_1279),
.B2(n_1255),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1163),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1274),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1127),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1102),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1102),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1274),
.Y(n_1346)
);

INVx5_ASAP7_75t_L g1347 ( 
.A(n_1197),
.Y(n_1347)
);

NOR3xp33_ASAP7_75t_L g1348 ( 
.A(n_1230),
.B(n_787),
.C(n_664),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1102),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1285),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1285),
.Y(n_1351)
);

AND3x2_ASAP7_75t_L g1352 ( 
.A(n_1127),
.B(n_550),
.C(n_548),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1193),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1287),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1109),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1287),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1183),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1241),
.B(n_751),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1286),
.B(n_1092),
.Y(n_1359)
);

XNOR2x2_ASAP7_75t_SL g1360 ( 
.A(n_1202),
.B(n_550),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1228),
.B(n_671),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1193),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1241),
.B(n_887),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1105),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1193),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1193),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1100),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1228),
.B(n_752),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1100),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1112),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1205),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1112),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1117),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1308),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1308),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1261),
.B(n_762),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1133),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1117),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1240),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1098),
.A2(n_612),
.B1(n_567),
.B2(n_1092),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1243),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1121),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1109),
.B(n_1029),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1245),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1176),
.B(n_922),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1121),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1099),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1136),
.B(n_1029),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1250),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1196),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1123),
.B(n_646),
.Y(n_1391)
);

XNOR2xp5_ASAP7_75t_L g1392 ( 
.A(n_1179),
.B(n_786),
.Y(n_1392)
);

BUFx10_ASAP7_75t_L g1393 ( 
.A(n_1178),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1233),
.B(n_1124),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1181),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1196),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1183),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1145),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1133),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1204),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1270),
.B(n_671),
.Y(n_1401)
);

INVxp33_ASAP7_75t_L g1402 ( 
.A(n_1147),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1186),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1182),
.B(n_975),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1320),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1183),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1132),
.B(n_736),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1270),
.B(n_763),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1261),
.B(n_776),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1160),
.B(n_697),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1182),
.B(n_993),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1204),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1173),
.A2(n_1029),
.B1(n_709),
.B2(n_712),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1211),
.B(n_993),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1165),
.B(n_519),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1255),
.A2(n_1321),
.B1(n_1211),
.B2(n_1200),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1208),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1136),
.B(n_1029),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1208),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1170),
.B(n_521),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1136),
.B(n_1080),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1214),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1214),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1187),
.B(n_527),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1219),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1219),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1227),
.B(n_1088),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1226),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1128),
.B(n_530),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1103),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1226),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1227),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1146),
.B(n_697),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1235),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1273),
.B(n_769),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1146),
.B(n_709),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1227),
.B(n_1088),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1234),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1235),
.Y(n_1439)
);

NOR2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1129),
.B(n_647),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_R g1441 ( 
.A(n_1135),
.B(n_993),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1239),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1186),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1234),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1239),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1242),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1242),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1251),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1255),
.A2(n_1060),
.B1(n_1073),
.B2(n_1022),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1215),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1251),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1212),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1254),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1222),
.B(n_1220),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1225),
.B(n_1073),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1248),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1225),
.B(n_1073),
.Y(n_1457)
);

INVxp67_ASAP7_75t_SL g1458 ( 
.A(n_1234),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1273),
.B(n_769),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1238),
.B(n_1073),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1248),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1120),
.A2(n_1060),
.B1(n_1022),
.B2(n_712),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1125),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1125),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1120),
.A2(n_1200),
.B1(n_1238),
.B2(n_1262),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1262),
.B(n_1089),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1120),
.A2(n_1060),
.B1(n_1022),
.B2(n_728),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1257),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1150),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1141),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1167),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1120),
.A2(n_1060),
.B1(n_728),
.B2(n_772),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1150),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1262),
.B(n_1089),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1158),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1301),
.B(n_1093),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_L g1477 ( 
.A(n_1120),
.B(n_553),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1156),
.B(n_536),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1168),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1158),
.Y(n_1480)
);

AND2x6_ASAP7_75t_L g1481 ( 
.A(n_1171),
.B(n_731),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1293),
.A2(n_772),
.B1(n_731),
.B2(n_998),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1161),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1161),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1276),
.B(n_769),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1189),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1198),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1164),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1198),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1106),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1301),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1301),
.B(n_1093),
.Y(n_1492)
);

BUFx8_ASAP7_75t_SL g1493 ( 
.A(n_1178),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1197),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1164),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1198),
.B(n_848),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1191),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1101),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1194),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1104),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1201),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1293),
.A2(n_774),
.B1(n_804),
.B2(n_799),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1199),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1213),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1108),
.B(n_1011),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1141),
.Y(n_1506)
);

BUFx4f_ASAP7_75t_L g1507 ( 
.A(n_1120),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1174),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1174),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1141),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1141),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1141),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1217),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1244),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1256),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1113),
.B(n_1011),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1119),
.B(n_1011),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1201),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_L g1519 ( 
.A(n_1120),
.B(n_553),
.Y(n_1519)
);

AND2x6_ASAP7_75t_L g1520 ( 
.A(n_1122),
.B(n_532),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1180),
.Y(n_1521)
);

INVxp33_ASAP7_75t_L g1522 ( 
.A(n_1118),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1256),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1297),
.A2(n_998),
.B1(n_1007),
.B2(n_829),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1130),
.B(n_1011),
.Y(n_1525)
);

NAND2xp33_ASAP7_75t_SL g1526 ( 
.A(n_1260),
.B(n_774),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1276),
.B(n_769),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1201),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1223),
.B(n_537),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1131),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1232),
.B(n_538),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1152),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1200),
.A2(n_998),
.B1(n_1007),
.B2(n_1011),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1297),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1139),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1231),
.B(n_539),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1302),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1180),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1190),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1152),
.Y(n_1540)
);

NAND2xp33_ASAP7_75t_L g1541 ( 
.A(n_1200),
.B(n_553),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1140),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1142),
.B(n_1011),
.Y(n_1543)
);

INVx4_ASAP7_75t_L g1544 ( 
.A(n_1152),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1190),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1195),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1236),
.B(n_540),
.Y(n_1547)
);

AND3x2_ASAP7_75t_L g1548 ( 
.A(n_1143),
.B(n_563),
.C(n_559),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1277),
.B(n_784),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1151),
.B(n_998),
.Y(n_1550)
);

BUFx4f_ASAP7_75t_L g1551 ( 
.A(n_1200),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1157),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1267),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1159),
.B(n_998),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1263),
.B(n_998),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1265),
.B(n_998),
.Y(n_1556)
);

AO21x2_ASAP7_75t_L g1557 ( 
.A1(n_1271),
.A2(n_900),
.B(n_892),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1267),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1302),
.B(n_543),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1152),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1200),
.A2(n_775),
.B1(n_532),
.B2(n_826),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1277),
.B(n_784),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1101),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1269),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1269),
.Y(n_1565)
);

NAND2xp33_ASAP7_75t_SL g1566 ( 
.A(n_1126),
.B(n_581),
.Y(n_1566)
);

AO21x2_ASAP7_75t_L g1567 ( 
.A1(n_1275),
.A2(n_905),
.B(n_900),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1284),
.Y(n_1568)
);

INVx6_ASAP7_75t_L g1569 ( 
.A(n_1294),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1312),
.B(n_863),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1110),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1195),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1363),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1570),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1454),
.B(n_1252),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1394),
.B(n_1312),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1470),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1328),
.B(n_1314),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1335),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1335),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1337),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1470),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1343),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1331),
.B(n_1314),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1385),
.B(n_1218),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1337),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1338),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1343),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1416),
.A2(n_1315),
.B1(n_1247),
.B2(n_1249),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1338),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1458),
.B(n_1327),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1341),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1487),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1570),
.B(n_1172),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1341),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1470),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1327),
.B(n_1315),
.Y(n_1597)
);

AO22x2_ASAP7_75t_L g1598 ( 
.A1(n_1360),
.A2(n_1220),
.B1(n_1224),
.B2(n_1179),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1398),
.Y(n_1599)
);

AO22x2_ASAP7_75t_L g1600 ( 
.A1(n_1454),
.A2(n_1224),
.B1(n_563),
.B2(n_568),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1371),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1371),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1367),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1327),
.B(n_1246),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1355),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1379),
.Y(n_1606)
);

AO22x1_ASAP7_75t_L g1607 ( 
.A1(n_1391),
.A2(n_1259),
.B1(n_1258),
.B2(n_1253),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1470),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1379),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1407),
.B(n_1172),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1367),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1381),
.Y(n_1612)
);

AND2x6_ASAP7_75t_L g1613 ( 
.A(n_1330),
.B(n_775),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1326),
.B(n_1280),
.Y(n_1614)
);

AO22x2_ASAP7_75t_L g1615 ( 
.A1(n_1334),
.A2(n_568),
.B1(n_574),
.B2(n_559),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1355),
.B(n_1246),
.Y(n_1616)
);

INVx4_ASAP7_75t_SL g1617 ( 
.A(n_1481),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1350),
.A2(n_1282),
.B1(n_1280),
.B2(n_1259),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1487),
.B(n_1268),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1398),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1369),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1381),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1355),
.B(n_1247),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1384),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1384),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1501),
.B(n_1278),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1491),
.B(n_1249),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1491),
.B(n_1281),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1491),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1369),
.Y(n_1630)
);

INVx4_ASAP7_75t_L g1631 ( 
.A(n_1470),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1501),
.B(n_1518),
.Y(n_1632)
);

AO22x2_ASAP7_75t_L g1633 ( 
.A1(n_1334),
.A2(n_575),
.B1(n_579),
.B2(n_574),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1452),
.B(n_1283),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1389),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1389),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1496),
.B(n_1175),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1496),
.B(n_1408),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1364),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1370),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1370),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1500),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1372),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1372),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1429),
.B(n_1253),
.C(n_1252),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1506),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1500),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1364),
.B(n_1522),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1471),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1350),
.A2(n_1282),
.B1(n_1258),
.B2(n_1290),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1373),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1373),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1450),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1518),
.B(n_1288),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1408),
.B(n_1290),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1514),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1471),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1403),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1432),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1479),
.Y(n_1660)
);

AO22x2_ASAP7_75t_L g1661 ( 
.A1(n_1405),
.A2(n_579),
.B1(n_588),
.B2(n_575),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1432),
.B(n_1292),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1506),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1403),
.B(n_1295),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1452),
.B(n_1299),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1378),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1432),
.Y(n_1667)
);

INVx4_ASAP7_75t_SL g1668 ( 
.A(n_1481),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1357),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1351),
.A2(n_1303),
.B1(n_1309),
.B2(n_1307),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1455),
.A2(n_1200),
.B1(n_588),
.B2(n_603),
.Y(n_1671)
);

NAND2x1p5_ASAP7_75t_L g1672 ( 
.A(n_1507),
.B(n_1317),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1357),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1438),
.B(n_1444),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1479),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1486),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1443),
.B(n_1310),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1486),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1443),
.B(n_1319),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1497),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1351),
.B(n_1354),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1354),
.B(n_1356),
.Y(n_1682)
);

AO22x2_ASAP7_75t_L g1683 ( 
.A1(n_1330),
.A2(n_603),
.B1(n_605),
.B2(n_591),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1497),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1450),
.B(n_1175),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1395),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1499),
.Y(n_1687)
);

OR2x2_ASAP7_75t_SL g1688 ( 
.A(n_1569),
.B(n_1216),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1499),
.Y(n_1689)
);

AO22x2_ASAP7_75t_L g1690 ( 
.A1(n_1332),
.A2(n_605),
.B1(n_609),
.B2(n_591),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1503),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1438),
.B(n_1323),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1503),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1378),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1456),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1559),
.B(n_1184),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1498),
.Y(n_1697)
);

NAND2x1p5_ASAP7_75t_L g1698 ( 
.A(n_1507),
.B(n_1325),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1356),
.B(n_1116),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1456),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1410),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1563),
.B(n_1110),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1438),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1374),
.B(n_1306),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1415),
.B(n_1184),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1382),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1506),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1433),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1420),
.B(n_1144),
.Y(n_1709)
);

AND2x6_ASAP7_75t_L g1710 ( 
.A(n_1332),
.B(n_775),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1382),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1433),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1504),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1444),
.B(n_1313),
.Y(n_1714)
);

BUFx4f_ASAP7_75t_L g1715 ( 
.A(n_1569),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1424),
.B(n_1144),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1504),
.Y(n_1717)
);

INVx8_ASAP7_75t_L g1718 ( 
.A(n_1433),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1513),
.Y(n_1719)
);

INVx8_ASAP7_75t_L g1720 ( 
.A(n_1433),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1571),
.B(n_1361),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1513),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1444),
.B(n_1324),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1374),
.B(n_1148),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1375),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1375),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1455),
.A2(n_609),
.B1(n_632),
.B2(n_610),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1390),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1461),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1348),
.B(n_1149),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1386),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1390),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1386),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1397),
.B(n_1148),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1534),
.B(n_1149),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1359),
.B(n_1294),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1402),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1400),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1506),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1400),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1534),
.B(n_1153),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1412),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1506),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1397),
.B(n_1153),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1396),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1412),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1453),
.B(n_1294),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1417),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1436),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1417),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1423),
.Y(n_1751)
);

AO22x2_ASAP7_75t_L g1752 ( 
.A1(n_1333),
.A2(n_632),
.B1(n_635),
.B2(n_610),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1423),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1396),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1507),
.B(n_1154),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1425),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1502),
.B(n_1537),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1419),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1425),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1419),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1461),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_SL g1762 ( 
.A(n_1387),
.B(n_1099),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1453),
.B(n_1284),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1410),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1426),
.Y(n_1765)
);

INVx4_ASAP7_75t_L g1766 ( 
.A(n_1512),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1406),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1426),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1468),
.B(n_1300),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1537),
.B(n_1166),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1428),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1457),
.A2(n_635),
.B1(n_649),
.B2(n_636),
.Y(n_1772)
);

BUFx4f_ASAP7_75t_L g1773 ( 
.A(n_1569),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1406),
.B(n_1154),
.Y(n_1774)
);

INVx4_ASAP7_75t_L g1775 ( 
.A(n_1512),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1489),
.B(n_1162),
.Y(n_1776)
);

OR2x6_ASAP7_75t_L g1777 ( 
.A(n_1569),
.B(n_647),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1422),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1551),
.B(n_1162),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1428),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1336),
.B(n_1361),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1468),
.B(n_1300),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1439),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1422),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1489),
.B(n_1166),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1439),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1342),
.B(n_1305),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1342),
.B(n_1305),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1410),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1442),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1526),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1431),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1346),
.B(n_1311),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1340),
.A2(n_1129),
.B1(n_1137),
.B2(n_1134),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1528),
.B(n_1134),
.Y(n_1795)
);

BUFx8_ASAP7_75t_SL g1796 ( 
.A(n_1493),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1478),
.B(n_1115),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1512),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1361),
.B(n_1115),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1361),
.B(n_1291),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1352),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1431),
.Y(n_1802)
);

AND3x1_ASAP7_75t_L g1803 ( 
.A(n_1529),
.B(n_649),
.C(n_636),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1442),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1346),
.B(n_1528),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1387),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1401),
.B(n_1137),
.Y(n_1807)
);

NAND2xp33_ASAP7_75t_L g1808 ( 
.A(n_1465),
.B(n_553),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1436),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1445),
.Y(n_1810)
);

NAND3x1_ASAP7_75t_L g1811 ( 
.A(n_1531),
.B(n_653),
.C(n_652),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1457),
.A2(n_1460),
.B1(n_1411),
.B2(n_1414),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1445),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1512),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1462),
.A2(n_1138),
.B1(n_1322),
.B2(n_1316),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1446),
.Y(n_1816)
);

INVx2_ASAP7_75t_SL g1817 ( 
.A(n_1548),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1430),
.B(n_1490),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1434),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1512),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1460),
.A2(n_1411),
.B1(n_1414),
.B2(n_1404),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1446),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1576),
.B(n_1410),
.Y(n_1823)
);

OAI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1812),
.A2(n_1404),
.B(n_1388),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1578),
.B(n_1584),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1715),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1634),
.B(n_1530),
.Y(n_1827)
);

INVx8_ASAP7_75t_L g1828 ( 
.A(n_1718),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1638),
.B(n_1401),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1579),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1631),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1579),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1605),
.A2(n_1551),
.B(n_1418),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1590),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1727),
.A2(n_1481),
.B1(n_1401),
.B2(n_1535),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1665),
.B(n_1542),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1602),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1727),
.A2(n_1481),
.B1(n_1401),
.B2(n_1552),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1590),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1573),
.B(n_1358),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1812),
.A2(n_1821),
.B(n_1808),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1681),
.B(n_1536),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1681),
.B(n_1547),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1772),
.A2(n_1481),
.B1(n_1519),
.B2(n_1477),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1603),
.Y(n_1845)
);

NAND2xp33_ASAP7_75t_L g1846 ( 
.A(n_1736),
.B(n_1481),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1602),
.Y(n_1847)
);

INVx5_ASAP7_75t_L g1848 ( 
.A(n_1577),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1639),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1603),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1580),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1614),
.A2(n_1441),
.B1(n_1459),
.B2(n_1435),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1695),
.B(n_1436),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1581),
.Y(n_1854)
);

NOR2x1p5_ASAP7_75t_L g1855 ( 
.A(n_1747),
.B(n_1138),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1599),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1586),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1681),
.B(n_1436),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1611),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1587),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1614),
.A2(n_1527),
.B1(n_1549),
.B2(n_1485),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1620),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1573),
.B(n_1562),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1583),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1682),
.B(n_1413),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1588),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1601),
.Y(n_1867)
);

BUFx5_ASAP7_75t_L g1868 ( 
.A(n_1613),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1610),
.B(n_1368),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1682),
.B(n_1339),
.Y(n_1870)
);

NOR2x1p5_ASAP7_75t_L g1871 ( 
.A(n_1575),
.B(n_1192),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1611),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1682),
.B(n_1339),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1725),
.B(n_1339),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1605),
.B(n_1551),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1592),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1594),
.B(n_1440),
.Y(n_1877)
);

NAND2xp33_ASAP7_75t_L g1878 ( 
.A(n_1577),
.B(n_1481),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1595),
.Y(n_1879)
);

BUFx6f_ASAP7_75t_L g1880 ( 
.A(n_1577),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1621),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1574),
.A2(n_1380),
.B1(n_1524),
.B2(n_1229),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1726),
.B(n_1349),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1574),
.B(n_1376),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1605),
.B(n_1377),
.Y(n_1885)
);

INVx5_ASAP7_75t_L g1886 ( 
.A(n_1577),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1715),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1606),
.B(n_1349),
.Y(n_1888)
);

NAND2xp33_ASAP7_75t_L g1889 ( 
.A(n_1582),
.B(n_1467),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1653),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1695),
.B(n_1448),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1609),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1781),
.A2(n_1705),
.B1(n_1585),
.B2(n_1645),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1781),
.A2(n_1566),
.B1(n_1409),
.B2(n_1155),
.Y(n_1894)
);

NAND3xp33_ASAP7_75t_SL g1895 ( 
.A(n_1696),
.B(n_1111),
.C(n_1229),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1796),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1612),
.Y(n_1897)
);

AO22x1_ASAP7_75t_L g1898 ( 
.A1(n_1655),
.A2(n_1207),
.B1(n_1209),
.B2(n_1192),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1622),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1621),
.Y(n_1900)
);

O2A1O1Ixp5_ASAP7_75t_L g1901 ( 
.A1(n_1627),
.A2(n_1516),
.B(n_1517),
.C(n_1505),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1629),
.A2(n_1383),
.B(n_1510),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1757),
.A2(n_1519),
.B(n_1541),
.C(n_1477),
.Y(n_1903)
);

OR2x6_ASAP7_75t_L g1904 ( 
.A(n_1718),
.B(n_1333),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1772),
.A2(n_1541),
.B1(n_1451),
.B2(n_1448),
.Y(n_1905)
);

O2A1O1Ixp5_ASAP7_75t_L g1906 ( 
.A1(n_1627),
.A2(n_1543),
.B(n_1525),
.C(n_1427),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1624),
.B(n_1349),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1625),
.B(n_1353),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1635),
.B(n_1353),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1808),
.A2(n_1451),
.B1(n_777),
.B2(n_805),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1796),
.Y(n_1911)
);

OR2x6_ASAP7_75t_SL g1912 ( 
.A(n_1794),
.B(n_1207),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1636),
.B(n_1353),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1649),
.B(n_1657),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1660),
.B(n_1366),
.Y(n_1915)
);

AO22x1_ASAP7_75t_L g1916 ( 
.A1(n_1655),
.A2(n_1209),
.B1(n_1237),
.B2(n_1392),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1615),
.A2(n_777),
.B1(n_805),
.B2(n_746),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1637),
.B(n_1393),
.Y(n_1918)
);

NOR2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1721),
.B(n_1237),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1589),
.A2(n_1556),
.B1(n_1555),
.B2(n_1550),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_SL g1921 ( 
.A1(n_1598),
.A2(n_1393),
.B1(n_784),
.B2(n_1392),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1685),
.B(n_1393),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1675),
.Y(n_1923)
);

NOR3xp33_ASAP7_75t_L g1924 ( 
.A(n_1607),
.B(n_930),
.C(n_902),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1676),
.Y(n_1925)
);

NOR2x2_ASAP7_75t_L g1926 ( 
.A(n_1777),
.B(n_1344),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1630),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1615),
.A2(n_746),
.B1(n_1472),
.B2(n_1557),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1630),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1757),
.A2(n_1554),
.B1(n_1482),
.B2(n_1447),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1615),
.A2(n_1567),
.B1(n_1557),
.B2(n_652),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1631),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1629),
.B(n_1377),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1800),
.A2(n_1447),
.B1(n_1434),
.B2(n_1515),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1640),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1629),
.B(n_1377),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1633),
.A2(n_1567),
.B1(n_1557),
.B2(n_653),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1773),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1678),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1686),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1633),
.A2(n_1567),
.B1(n_654),
.B2(n_668),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1656),
.A2(n_1514),
.B1(n_597),
.B2(n_619),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1680),
.B(n_1366),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1684),
.B(n_1366),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1633),
.A2(n_654),
.B1(n_668),
.B2(n_658),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1687),
.B(n_1421),
.Y(n_1946)
);

AND2x6_ASAP7_75t_L g1947 ( 
.A(n_1659),
.B(n_1344),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1597),
.B(n_1377),
.Y(n_1948)
);

INVx3_ASAP7_75t_L g1949 ( 
.A(n_1631),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1689),
.B(n_1437),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1640),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1691),
.B(n_1466),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1693),
.B(n_1474),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1641),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1713),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1704),
.B(n_1632),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1717),
.B(n_1476),
.Y(n_1957)
);

NAND3xp33_ASAP7_75t_SL g1958 ( 
.A(n_1797),
.B(n_549),
.C(n_546),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1719),
.B(n_1492),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1683),
.A2(n_669),
.B1(n_672),
.B2(n_658),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1582),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1722),
.B(n_1515),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1704),
.B(n_1523),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1639),
.B(n_1345),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1728),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1743),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1732),
.Y(n_1967)
);

INVx4_ASAP7_75t_L g1968 ( 
.A(n_1773),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1704),
.B(n_1523),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1738),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1740),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1683),
.A2(n_672),
.B1(n_673),
.B2(n_669),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1648),
.B(n_1345),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1641),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1742),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_SL g1976 ( 
.A(n_1762),
.B(n_784),
.Y(n_1976)
);

INVx8_ASAP7_75t_L g1977 ( 
.A(n_1718),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1821),
.B(n_1553),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1582),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1683),
.A2(n_677),
.B1(n_681),
.B2(n_673),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1737),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1690),
.A2(n_677),
.B1(n_687),
.B2(n_681),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1697),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1632),
.B(n_1377),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1648),
.B(n_1365),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1690),
.A2(n_687),
.B1(n_698),
.B2(n_694),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1709),
.B(n_1716),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1800),
.A2(n_1553),
.B1(n_1564),
.B2(n_1558),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1669),
.B(n_1673),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1746),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1643),
.Y(n_1991)
);

INVx5_ASAP7_75t_L g1992 ( 
.A(n_1582),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1690),
.A2(n_694),
.B1(n_700),
.B2(n_698),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1669),
.B(n_1558),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1632),
.B(n_1399),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1699),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1699),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1673),
.B(n_1564),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1748),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1735),
.B(n_676),
.Y(n_2000)
);

INVxp67_ASAP7_75t_SL g2001 ( 
.A(n_1596),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1700),
.B(n_1532),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1750),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1650),
.B(n_1362),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1741),
.B(n_676),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1618),
.B(n_1362),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1767),
.B(n_1565),
.Y(n_2007)
);

A2O1A1Ixp33_ASAP7_75t_L g2008 ( 
.A1(n_1671),
.A2(n_1561),
.B(n_1449),
.C(n_1329),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1767),
.B(n_1565),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1619),
.B(n_1568),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1751),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1753),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1643),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1596),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1752),
.A2(n_700),
.B1(n_704),
.B2(n_703),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1593),
.B(n_1399),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1619),
.B(n_1568),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1770),
.B(n_1799),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_SL g2019 ( 
.A1(n_1656),
.A2(n_582),
.B1(n_602),
.B2(n_558),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_1658),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1752),
.A2(n_703),
.B1(n_718),
.B2(n_704),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1619),
.B(n_1365),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1756),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1626),
.B(n_1463),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1759),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1593),
.B(n_1399),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1626),
.B(n_1463),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1644),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1626),
.B(n_1464),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1659),
.B(n_1399),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1644),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1765),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1667),
.B(n_1399),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1702),
.B(n_1464),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1699),
.B(n_676),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1701),
.A2(n_1540),
.B1(n_1560),
.B2(n_1532),
.Y(n_2036)
);

INVxp67_ASAP7_75t_SL g2037 ( 
.A(n_1596),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1853),
.B(n_1658),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1825),
.B(n_1664),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1940),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1845),
.Y(n_2041)
);

NAND3xp33_ASAP7_75t_SL g2042 ( 
.A(n_1976),
.B(n_1791),
.C(n_1806),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1892),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1897),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1848),
.Y(n_2045)
);

INVx1_ASAP7_75t_SL g2046 ( 
.A(n_1867),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1856),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1852),
.B(n_1805),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1890),
.B(n_1642),
.Y(n_2049)
);

INVx4_ASAP7_75t_L g2050 ( 
.A(n_1828),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1845),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_1848),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1899),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1827),
.B(n_1664),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1823),
.B(n_1701),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1850),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1837),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1850),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1872),
.Y(n_2059)
);

NOR3xp33_ASAP7_75t_SL g2060 ( 
.A(n_1958),
.B(n_1895),
.C(n_1882),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1853),
.B(n_1700),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1836),
.B(n_1664),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1987),
.B(n_1598),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1840),
.B(n_1677),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_R g2065 ( 
.A(n_1896),
.B(n_1911),
.Y(n_2065)
);

NOR3xp33_ASAP7_75t_SL g2066 ( 
.A(n_1882),
.B(n_557),
.C(n_551),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1840),
.B(n_1677),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1973),
.B(n_1677),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1872),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_2020),
.B(n_1729),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_1831),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1829),
.B(n_1598),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1900),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1923),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1981),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1925),
.Y(n_2076)
);

CKINVDCx20_ASAP7_75t_R g2077 ( 
.A(n_1856),
.Y(n_2077)
);

INVx4_ASAP7_75t_L g2078 ( 
.A(n_1828),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1939),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1955),
.Y(n_2080)
);

INVx1_ASAP7_75t_SL g2081 ( 
.A(n_1983),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1847),
.Y(n_2082)
);

OAI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1893),
.A2(n_1861),
.B1(n_1841),
.B2(n_1843),
.Y(n_2083)
);

INVx4_ASAP7_75t_L g2084 ( 
.A(n_1828),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_1864),
.Y(n_2085)
);

NOR3xp33_ASAP7_75t_SL g2086 ( 
.A(n_1863),
.B(n_564),
.C(n_560),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1900),
.Y(n_2087)
);

BUFx3_ASAP7_75t_L g2088 ( 
.A(n_1864),
.Y(n_2088)
);

OR2x6_ASAP7_75t_L g2089 ( 
.A(n_1977),
.B(n_1720),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1851),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1842),
.B(n_1604),
.Y(n_2091)
);

BUFx10_ASAP7_75t_L g2092 ( 
.A(n_1871),
.Y(n_2092)
);

NOR2xp67_ASAP7_75t_L g2093 ( 
.A(n_1894),
.B(n_1724),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1866),
.Y(n_2094)
);

NAND3xp33_ASAP7_75t_SL g2095 ( 
.A(n_1921),
.B(n_1789),
.C(n_1764),
.Y(n_2095)
);

INVxp33_ASAP7_75t_L g2096 ( 
.A(n_2034),
.Y(n_2096)
);

INVx8_ASAP7_75t_L g2097 ( 
.A(n_1977),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1884),
.B(n_1616),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1848),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1973),
.B(n_1679),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1985),
.B(n_1679),
.Y(n_2101)
);

AND2x4_ASAP7_75t_SL g2102 ( 
.A(n_1826),
.B(n_1777),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1854),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2020),
.B(n_1729),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_1884),
.B(n_1623),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1985),
.B(n_1679),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1857),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1860),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_SL g2109 ( 
.A(n_1866),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1876),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2018),
.B(n_1708),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1879),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2034),
.B(n_1818),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1965),
.Y(n_2114)
);

OR2x6_ASAP7_75t_L g2115 ( 
.A(n_1977),
.B(n_1720),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1863),
.B(n_1818),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1862),
.Y(n_2117)
);

INVx2_ASAP7_75t_SL g2118 ( 
.A(n_1919),
.Y(n_2118)
);

NOR3xp33_ASAP7_75t_SL g2119 ( 
.A(n_1942),
.B(n_569),
.C(n_565),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2004),
.B(n_1818),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_1849),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_2004),
.B(n_1764),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_1945),
.A2(n_1600),
.B1(n_1661),
.B2(n_1752),
.Y(n_2123)
);

INVx4_ASAP7_75t_L g2124 ( 
.A(n_1848),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2022),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1922),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_1996),
.B(n_1647),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_1886),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_L g2129 ( 
.A(n_1886),
.Y(n_2129)
);

CKINVDCx16_ASAP7_75t_R g2130 ( 
.A(n_1918),
.Y(n_2130)
);

NAND2xp33_ASAP7_75t_SL g2131 ( 
.A(n_1844),
.B(n_1826),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1967),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2006),
.B(n_1789),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2006),
.B(n_1761),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_1887),
.B(n_1724),
.Y(n_2135)
);

INVx5_ASAP7_75t_L g2136 ( 
.A(n_1947),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1970),
.Y(n_2137)
);

BUFx3_ASAP7_75t_L g2138 ( 
.A(n_1887),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1831),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1971),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1975),
.Y(n_2141)
);

INVx4_ASAP7_75t_L g2142 ( 
.A(n_1886),
.Y(n_2142)
);

NAND2xp33_ASAP7_75t_R g2143 ( 
.A(n_1877),
.B(n_1869),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_1945),
.A2(n_1600),
.B1(n_1661),
.B2(n_1768),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1964),
.B(n_1761),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1990),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_1938),
.B(n_1724),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_1858),
.B(n_1712),
.Y(n_2148)
);

NOR3xp33_ASAP7_75t_SL g2149 ( 
.A(n_2019),
.B(n_577),
.C(n_572),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1956),
.A2(n_1591),
.B1(n_1671),
.B2(n_1654),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1999),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_1938),
.B(n_1795),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_1997),
.B(n_1688),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1964),
.B(n_1654),
.Y(n_2154)
);

INVxp67_ASAP7_75t_SL g2155 ( 
.A(n_1889),
.Y(n_2155)
);

INVx1_ASAP7_75t_SL g2156 ( 
.A(n_2035),
.Y(n_2156)
);

NOR3xp33_ASAP7_75t_SL g2157 ( 
.A(n_1956),
.B(n_583),
.C(n_578),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_1886),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1914),
.B(n_1946),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_R g2160 ( 
.A(n_1968),
.B(n_1720),
.Y(n_2160)
);

NAND2x1p5_ASAP7_75t_L g2161 ( 
.A(n_1992),
.B(n_1743),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1912),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1968),
.B(n_1795),
.Y(n_2163)
);

BUFx2_ASAP7_75t_L g2164 ( 
.A(n_1891),
.Y(n_2164)
);

AND2x4_ASAP7_75t_SL g2165 ( 
.A(n_2002),
.B(n_1777),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1935),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_1992),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1950),
.B(n_1654),
.Y(n_2168)
);

NOR3xp33_ASAP7_75t_SL g2169 ( 
.A(n_1865),
.B(n_592),
.C(n_587),
.Y(n_2169)
);

AOI211xp5_ASAP7_75t_L g2170 ( 
.A1(n_1924),
.A2(n_1916),
.B(n_1898),
.C(n_1730),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1935),
.Y(n_2171)
);

BUFx2_ASAP7_75t_L g2172 ( 
.A(n_1891),
.Y(n_2172)
);

INVx4_ASAP7_75t_L g2173 ( 
.A(n_1992),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_1992),
.Y(n_2174)
);

BUFx4f_ASAP7_75t_L g2175 ( 
.A(n_1904),
.Y(n_2175)
);

BUFx8_ASAP7_75t_L g2176 ( 
.A(n_2000),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1954),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2003),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2011),
.Y(n_2179)
);

AOI221xp5_ASAP7_75t_L g2180 ( 
.A1(n_1917),
.A2(n_1803),
.B1(n_1600),
.B2(n_1661),
.C(n_1801),
.Y(n_2180)
);

INVx5_ASAP7_75t_L g2181 ( 
.A(n_1947),
.Y(n_2181)
);

BUFx2_ASAP7_75t_L g2182 ( 
.A(n_1926),
.Y(n_2182)
);

BUFx10_ASAP7_75t_L g2183 ( 
.A(n_1855),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2012),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1952),
.B(n_1628),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2023),
.Y(n_2186)
);

HB1xp67_ASAP7_75t_L g2187 ( 
.A(n_1870),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2002),
.B(n_1795),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2025),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_1873),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1953),
.B(n_1670),
.Y(n_2191)
);

INVx5_ASAP7_75t_L g2192 ( 
.A(n_1947),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1880),
.Y(n_2193)
);

BUFx2_ASAP7_75t_L g2194 ( 
.A(n_1904),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_1960),
.A2(n_1980),
.B1(n_1982),
.B2(n_1972),
.Y(n_2195)
);

BUFx3_ASAP7_75t_L g2196 ( 
.A(n_1904),
.Y(n_2196)
);

INVx3_ASAP7_75t_L g2197 ( 
.A(n_1932),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2032),
.Y(n_2198)
);

INVx6_ASAP7_75t_L g2199 ( 
.A(n_1880),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1830),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_1989),
.Y(n_2201)
);

INVx3_ASAP7_75t_L g2202 ( 
.A(n_1932),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1957),
.B(n_1749),
.Y(n_2203)
);

INVx3_ASAP7_75t_SL g2204 ( 
.A(n_2005),
.Y(n_2204)
);

NOR3xp33_ASAP7_75t_SL g2205 ( 
.A(n_1948),
.B(n_595),
.C(n_594),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1954),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_2010),
.B(n_1809),
.Y(n_2207)
);

BUFx12f_ASAP7_75t_L g2208 ( 
.A(n_1880),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1959),
.B(n_1785),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1991),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1832),
.Y(n_2211)
);

BUFx12f_ASAP7_75t_L g2212 ( 
.A(n_1880),
.Y(n_2212)
);

INVx5_ASAP7_75t_L g2213 ( 
.A(n_1947),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2017),
.B(n_1807),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_SL g2215 ( 
.A(n_1963),
.B(n_1734),
.Y(n_2215)
);

NAND2xp33_ASAP7_75t_SL g2216 ( 
.A(n_1844),
.B(n_1814),
.Y(n_2216)
);

HB1xp67_ASAP7_75t_L g2217 ( 
.A(n_1969),
.Y(n_2217)
);

BUFx2_ASAP7_75t_L g2218 ( 
.A(n_1961),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1834),
.Y(n_2219)
);

OR2x2_ASAP7_75t_SL g2220 ( 
.A(n_2024),
.B(n_1811),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_1949),
.B(n_1734),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1839),
.B(n_1785),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1824),
.B(n_1771),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1859),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1991),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1949),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2013),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2013),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_1988),
.B(n_1780),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2031),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2031),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_1835),
.A2(n_1838),
.B1(n_2008),
.B2(n_1905),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1881),
.Y(n_2233)
);

NOR3xp33_ASAP7_75t_SL g2234 ( 
.A(n_1948),
.B(n_601),
.C(n_600),
.Y(n_2234)
);

BUFx12f_ASAP7_75t_L g2235 ( 
.A(n_1961),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1961),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1927),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1929),
.Y(n_2238)
);

AND2x6_ASAP7_75t_SL g2239 ( 
.A(n_2027),
.B(n_1734),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1978),
.B(n_1744),
.Y(n_2240)
);

AOI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_2008),
.A2(n_1674),
.B(n_1714),
.Y(n_2241)
);

INVx3_ASAP7_75t_L g2242 ( 
.A(n_1966),
.Y(n_2242)
);

OR2x4_ASAP7_75t_L g2243 ( 
.A(n_1961),
.B(n_1707),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1951),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2029),
.B(n_1744),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1974),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2028),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1979),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1962),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1835),
.B(n_1744),
.Y(n_2250)
);

OAI22xp33_ASAP7_75t_L g2251 ( 
.A1(n_1994),
.A2(n_1786),
.B1(n_1790),
.B2(n_1783),
.Y(n_2251)
);

INVx4_ASAP7_75t_L g2252 ( 
.A(n_1979),
.Y(n_2252)
);

BUFx6f_ASAP7_75t_L g2253 ( 
.A(n_1979),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1998),
.Y(n_2254)
);

NAND2x1p5_ASAP7_75t_L g2255 ( 
.A(n_1966),
.B(n_1743),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1838),
.B(n_1774),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2007),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2009),
.Y(n_2258)
);

NAND2xp33_ASAP7_75t_SL g2259 ( 
.A(n_1979),
.B(n_1596),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1874),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_1903),
.A2(n_1723),
.B(n_1692),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_1960),
.A2(n_1810),
.B1(n_1813),
.B2(n_1804),
.Y(n_2262)
);

CKINVDCx6p67_ASAP7_75t_R g2263 ( 
.A(n_2014),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1883),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_R g2265 ( 
.A(n_1878),
.B(n_1667),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1888),
.B(n_1774),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1907),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_2014),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1908),
.Y(n_2269)
);

INVx4_ASAP7_75t_L g2270 ( 
.A(n_2014),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2075),
.Y(n_2271)
);

INVxp67_ASAP7_75t_SL g2272 ( 
.A(n_2057),
.Y(n_2272)
);

OAI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2195),
.A2(n_2232),
.B1(n_2123),
.B2(n_2159),
.Y(n_2273)
);

A2O1A1Ixp33_ASAP7_75t_L g2274 ( 
.A1(n_2060),
.A2(n_1846),
.B(n_1776),
.C(n_1785),
.Y(n_2274)
);

OAI21x1_ASAP7_75t_L g2275 ( 
.A1(n_2261),
.A2(n_1901),
.B(n_1906),
.Y(n_2275)
);

INVx1_ASAP7_75t_SL g2276 ( 
.A(n_2081),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2120),
.B(n_1972),
.Y(n_2277)
);

A2O1A1Ixp33_ASAP7_75t_L g2278 ( 
.A1(n_2060),
.A2(n_1776),
.B(n_1774),
.C(n_1986),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2249),
.B(n_1986),
.Y(n_2279)
);

AOI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2216),
.A2(n_1933),
.B(n_1885),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2039),
.B(n_1776),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2261),
.A2(n_1902),
.B(n_1833),
.Y(n_2282)
);

AOI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2216),
.A2(n_1933),
.B(n_1885),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2043),
.Y(n_2284)
);

AO31x2_ASAP7_75t_L g2285 ( 
.A1(n_2241),
.A2(n_1815),
.A3(n_1788),
.B(n_1793),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2044),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2195),
.A2(n_2123),
.B1(n_2144),
.B2(n_1982),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2125),
.B(n_1980),
.Y(n_2288)
);

OAI21x1_ASAP7_75t_L g2289 ( 
.A1(n_2241),
.A2(n_1936),
.B(n_2030),
.Y(n_2289)
);

HB1xp67_ASAP7_75t_L g2290 ( 
.A(n_2057),
.Y(n_2290)
);

OAI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2144),
.A2(n_2015),
.B1(n_2021),
.B2(n_1993),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_2045),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_SL g2293 ( 
.A1(n_2155),
.A2(n_1775),
.B(n_1766),
.Y(n_2293)
);

AOI21x1_ASAP7_75t_L g2294 ( 
.A1(n_2048),
.A2(n_1936),
.B(n_2033),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2125),
.B(n_2083),
.Y(n_2295)
);

NAND2x1p5_ASAP7_75t_L g2296 ( 
.A(n_2136),
.B(n_1984),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2083),
.B(n_1993),
.Y(n_2297)
);

AND3x4_ASAP7_75t_L g2298 ( 
.A(n_2119),
.B(n_1817),
.C(n_1811),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2155),
.A2(n_1930),
.B(n_1920),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2111),
.B(n_1917),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2113),
.A2(n_2015),
.B1(n_2021),
.B2(n_1905),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2041),
.Y(n_2302)
);

AOI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_2131),
.A2(n_1875),
.B(n_1995),
.Y(n_2303)
);

AOI21x1_ASAP7_75t_L g2304 ( 
.A1(n_2048),
.A2(n_2033),
.B(n_2030),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2122),
.B(n_1941),
.Y(n_2305)
);

OAI21x1_ASAP7_75t_L g2306 ( 
.A1(n_2223),
.A2(n_2026),
.B(n_2016),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_SL g2307 ( 
.A1(n_2150),
.A2(n_1775),
.B(n_1766),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2122),
.B(n_1941),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2051),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_2077),
.Y(n_2310)
);

OAI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2098),
.A2(n_1934),
.B(n_1984),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2063),
.B(n_2096),
.Y(n_2312)
);

OAI21x1_ASAP7_75t_L g2313 ( 
.A1(n_2223),
.A2(n_2026),
.B(n_2016),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2133),
.B(n_1931),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_SL g2315 ( 
.A(n_2136),
.B(n_1766),
.Y(n_2315)
);

OAI21x1_ASAP7_75t_L g2316 ( 
.A1(n_2091),
.A2(n_1995),
.B(n_1787),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2131),
.A2(n_2185),
.B(n_2105),
.Y(n_2317)
);

INVx3_ASAP7_75t_L g2318 ( 
.A(n_2045),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2180),
.A2(n_613),
.B1(n_614),
.B2(n_607),
.C(n_606),
.Y(n_2319)
);

AOI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2185),
.A2(n_1875),
.B(n_1909),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2053),
.Y(n_2321)
);

NAND3xp33_ASAP7_75t_L g2322 ( 
.A(n_2066),
.B(n_1910),
.C(n_625),
.Y(n_2322)
);

OAI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2096),
.A2(n_1928),
.B1(n_1937),
.B2(n_1931),
.Y(n_2323)
);

OAI21x1_ASAP7_75t_L g2324 ( 
.A1(n_2091),
.A2(n_1769),
.B(n_1763),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2049),
.B(n_2130),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2072),
.B(n_1910),
.Y(n_2326)
);

OAI21x1_ASAP7_75t_L g2327 ( 
.A1(n_2229),
.A2(n_1782),
.B(n_1662),
.Y(n_2327)
);

OAI21x1_ASAP7_75t_L g2328 ( 
.A1(n_2229),
.A2(n_2105),
.B(n_2098),
.Y(n_2328)
);

INVxp67_ASAP7_75t_L g2329 ( 
.A(n_2040),
.Y(n_2329)
);

AO22x1_ASAP7_75t_L g2330 ( 
.A1(n_2176),
.A2(n_628),
.B1(n_630),
.B2(n_620),
.Y(n_2330)
);

OAI21x1_ASAP7_75t_L g2331 ( 
.A1(n_2134),
.A2(n_1662),
.B(n_1672),
.Y(n_2331)
);

AOI221x1_ASAP7_75t_L g2332 ( 
.A1(n_2095),
.A2(n_1822),
.B1(n_1816),
.B2(n_740),
.C(n_743),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2116),
.B(n_1672),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2074),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2254),
.B(n_2257),
.Y(n_2335)
);

AOI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_2191),
.A2(n_1915),
.B(n_1913),
.Y(n_2336)
);

INVx3_ASAP7_75t_L g2337 ( 
.A(n_2045),
.Y(n_2337)
);

AOI21xp33_ASAP7_75t_L g2338 ( 
.A1(n_2143),
.A2(n_1937),
.B(n_1928),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2076),
.Y(n_2339)
);

OAI22x1_ASAP7_75t_L g2340 ( 
.A1(n_2204),
.A2(n_2036),
.B1(n_725),
.B2(n_740),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_2045),
.Y(n_2341)
);

NAND2x1p5_ASAP7_75t_L g2342 ( 
.A(n_2136),
.B(n_2014),
.Y(n_2342)
);

OAI21x1_ASAP7_75t_L g2343 ( 
.A1(n_2255),
.A2(n_2240),
.B(n_1698),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2258),
.B(n_1943),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2093),
.A2(n_1755),
.B1(n_1779),
.B2(n_1698),
.Y(n_2345)
);

AO21x1_ASAP7_75t_L g2346 ( 
.A1(n_2251),
.A2(n_1944),
.B(n_1779),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2217),
.B(n_2054),
.Y(n_2347)
);

OAI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2266),
.A2(n_1710),
.B(n_1613),
.Y(n_2348)
);

O2A1O1Ixp5_ASAP7_75t_L g2349 ( 
.A1(n_2251),
.A2(n_1755),
.B(n_2037),
.C(n_2001),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2136),
.A2(n_1775),
.B(n_1511),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2079),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2217),
.B(n_1754),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2214),
.B(n_969),
.Y(n_2353)
);

OAI21x1_ASAP7_75t_L g2354 ( 
.A1(n_2255),
.A2(n_1703),
.B(n_1652),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_2052),
.Y(n_2355)
);

AOI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_2181),
.A2(n_2213),
.B(n_2192),
.Y(n_2356)
);

BUFx2_ASAP7_75t_L g2357 ( 
.A(n_2088),
.Y(n_2357)
);

OAI21x1_ASAP7_75t_L g2358 ( 
.A1(n_2260),
.A2(n_1703),
.B(n_1652),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2080),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2090),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2181),
.A2(n_2213),
.B(n_2192),
.Y(n_2361)
);

OAI21x1_ASAP7_75t_SL g2362 ( 
.A1(n_2250),
.A2(n_1666),
.B(n_1651),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2070),
.B(n_1651),
.Y(n_2363)
);

NOR2x1p5_ASAP7_75t_L g2364 ( 
.A(n_2095),
.B(n_1666),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2064),
.B(n_1694),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2103),
.Y(n_2366)
);

AO31x2_ASAP7_75t_L g2367 ( 
.A1(n_2266),
.A2(n_1511),
.A3(n_1544),
.B(n_1510),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2214),
.B(n_969),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2181),
.A2(n_1511),
.B(n_1510),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2062),
.B(n_1802),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2067),
.B(n_1802),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2181),
.A2(n_1544),
.B(n_1814),
.Y(n_2372)
);

INVx4_ASAP7_75t_L g2373 ( 
.A(n_2052),
.Y(n_2373)
);

OAI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_2055),
.A2(n_1710),
.B(n_1613),
.Y(n_2374)
);

INVx3_ASAP7_75t_SL g2375 ( 
.A(n_2126),
.Y(n_2375)
);

OAI21x1_ASAP7_75t_L g2376 ( 
.A1(n_2269),
.A2(n_1706),
.B(n_1694),
.Y(n_2376)
);

OAI21x1_ASAP7_75t_L g2377 ( 
.A1(n_2056),
.A2(n_1711),
.B(n_1706),
.Y(n_2377)
);

OAI21x1_ASAP7_75t_L g2378 ( 
.A1(n_2058),
.A2(n_2069),
.B(n_2059),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2192),
.A2(n_1544),
.B(n_1820),
.Y(n_2379)
);

INVx3_ASAP7_75t_L g2380 ( 
.A(n_2052),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2192),
.A2(n_1646),
.B(n_1608),
.Y(n_2381)
);

INVx4_ASAP7_75t_L g2382 ( 
.A(n_2052),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2143),
.A2(n_631),
.B1(n_634),
.B2(n_633),
.Y(n_2383)
);

O2A1O1Ixp5_ASAP7_75t_L g2384 ( 
.A1(n_2055),
.A2(n_1731),
.B(n_1733),
.C(n_1711),
.Y(n_2384)
);

OAI22x1_ASAP7_75t_L g2385 ( 
.A1(n_2204),
.A2(n_725),
.B1(n_743),
.B2(n_718),
.Y(n_2385)
);

INVx4_ASAP7_75t_L g2386 ( 
.A(n_2099),
.Y(n_2386)
);

AO22x1_ASAP7_75t_L g2387 ( 
.A1(n_2176),
.A2(n_638),
.B1(n_639),
.B2(n_637),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2213),
.A2(n_1814),
.B(n_1798),
.Y(n_2388)
);

INVx5_ASAP7_75t_L g2389 ( 
.A(n_2099),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2068),
.B(n_1731),
.Y(n_2390)
);

AOI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2213),
.A2(n_2259),
.B(n_2209),
.Y(n_2391)
);

AO31x2_ASAP7_75t_L g2392 ( 
.A1(n_2256),
.A2(n_1745),
.A3(n_1754),
.B(n_1733),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2107),
.Y(n_2393)
);

O2A1O1Ixp5_ASAP7_75t_L g2394 ( 
.A1(n_2175),
.A2(n_2145),
.B(n_2259),
.C(n_2154),
.Y(n_2394)
);

AOI21x1_ASAP7_75t_L g2395 ( 
.A1(n_2194),
.A2(n_1819),
.B(n_1758),
.Y(n_2395)
);

AO31x2_ASAP7_75t_L g2396 ( 
.A1(n_2264),
.A2(n_1758),
.A3(n_1760),
.B(n_1745),
.Y(n_2396)
);

INVx1_ASAP7_75t_SL g2397 ( 
.A(n_2046),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2168),
.A2(n_1820),
.B(n_1646),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2203),
.B(n_2127),
.Y(n_2399)
);

A2O1A1Ixp33_ASAP7_75t_L g2400 ( 
.A1(n_2066),
.A2(n_753),
.B(n_754),
.C(n_744),
.Y(n_2400)
);

AOI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2215),
.A2(n_1820),
.B(n_1646),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2100),
.B(n_1760),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2101),
.B(n_1778),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2106),
.B(n_1778),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2156),
.A2(n_640),
.B1(n_643),
.B2(n_641),
.Y(n_2405)
);

A2O1A1Ixp33_ASAP7_75t_L g2406 ( 
.A1(n_2086),
.A2(n_753),
.B(n_754),
.C(n_744),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2187),
.B(n_2190),
.Y(n_2407)
);

A2O1A1Ixp33_ASAP7_75t_L g2408 ( 
.A1(n_2086),
.A2(n_757),
.B(n_765),
.C(n_756),
.Y(n_2408)
);

OAI21x1_ASAP7_75t_L g2409 ( 
.A1(n_2073),
.A2(n_1792),
.B(n_1784),
.Y(n_2409)
);

OAI21x1_ASAP7_75t_L g2410 ( 
.A1(n_2087),
.A2(n_1792),
.B(n_1784),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2187),
.B(n_1819),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2190),
.B(n_1947),
.Y(n_2412)
);

A2O1A1Ixp33_ASAP7_75t_L g2413 ( 
.A1(n_2205),
.A2(n_757),
.B(n_765),
.C(n_756),
.Y(n_2413)
);

AOI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2175),
.A2(n_2245),
.B(n_2267),
.Y(n_2414)
);

BUFx2_ASAP7_75t_L g2415 ( 
.A(n_2088),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2262),
.B(n_1868),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2262),
.B(n_1868),
.Y(n_2417)
);

AOI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2222),
.A2(n_1814),
.B(n_1798),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2161),
.A2(n_1820),
.B(n_1798),
.Y(n_2419)
);

OAI21x1_ASAP7_75t_L g2420 ( 
.A1(n_2166),
.A2(n_1540),
.B(n_1532),
.Y(n_2420)
);

OAI21x1_ASAP7_75t_L g2421 ( 
.A1(n_2171),
.A2(n_1560),
.B(n_1540),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2200),
.B(n_1868),
.Y(n_2422)
);

AOI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_2161),
.A2(n_1646),
.B(n_1608),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2201),
.B(n_2153),
.Y(n_2424)
);

OAI21x1_ASAP7_75t_L g2425 ( 
.A1(n_2177),
.A2(n_1560),
.B(n_1473),
.Y(n_2425)
);

INVx2_ASAP7_75t_SL g2426 ( 
.A(n_2117),
.Y(n_2426)
);

AOI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_2221),
.A2(n_1663),
.B(n_1608),
.Y(n_2427)
);

AOI221xp5_ASAP7_75t_L g2428 ( 
.A1(n_2042),
.A2(n_659),
.B1(n_660),
.B2(n_657),
.C(n_651),
.Y(n_2428)
);

OAI21x1_ASAP7_75t_L g2429 ( 
.A1(n_2206),
.A2(n_1473),
.B(n_1469),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2220),
.A2(n_1663),
.B1(n_1707),
.B2(n_1608),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2211),
.B(n_1868),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2108),
.Y(n_2432)
);

INVx6_ASAP7_75t_L g2433 ( 
.A(n_2183),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_2138),
.Y(n_2434)
);

OAI21x1_ASAP7_75t_L g2435 ( 
.A1(n_2210),
.A2(n_1475),
.B(n_1469),
.Y(n_2435)
);

AOI21xp33_ASAP7_75t_L g2436 ( 
.A1(n_2207),
.A2(n_771),
.B(n_768),
.Y(n_2436)
);

AOI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2221),
.A2(n_1707),
.B(n_1663),
.Y(n_2437)
);

A2O1A1Ixp33_ASAP7_75t_L g2438 ( 
.A1(n_2205),
.A2(n_771),
.B(n_783),
.C(n_768),
.Y(n_2438)
);

INVx1_ASAP7_75t_SL g2439 ( 
.A(n_2085),
.Y(n_2439)
);

AO31x2_ASAP7_75t_L g2440 ( 
.A1(n_2219),
.A2(n_1480),
.A3(n_1483),
.B(n_1475),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2110),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2207),
.B(n_1868),
.Y(n_2442)
);

AO21x2_ASAP7_75t_L g2443 ( 
.A1(n_2234),
.A2(n_1483),
.B(n_1480),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2138),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2070),
.B(n_1617),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2148),
.B(n_676),
.Y(n_2446)
);

OAI22xp5_ASAP7_75t_L g2447 ( 
.A1(n_2112),
.A2(n_1707),
.B1(n_1739),
.B2(n_1663),
.Y(n_2447)
);

INVx3_ASAP7_75t_L g2448 ( 
.A(n_2099),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2114),
.B(n_1868),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2132),
.Y(n_2450)
);

A2O1A1Ixp33_ASAP7_75t_L g2451 ( 
.A1(n_2234),
.A2(n_790),
.B(n_795),
.C(n_783),
.Y(n_2451)
);

AOI21x1_ASAP7_75t_L g2452 ( 
.A1(n_2128),
.A2(n_1488),
.B(n_1484),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_SL g2453 ( 
.A1(n_2182),
.A2(n_705),
.B1(n_795),
.B2(n_790),
.Y(n_2453)
);

BUFx4_ASAP7_75t_SL g2454 ( 
.A(n_2236),
.Y(n_2454)
);

OAI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2157),
.A2(n_1710),
.B(n_1613),
.Y(n_2455)
);

OAI21xp5_ASAP7_75t_L g2456 ( 
.A1(n_2157),
.A2(n_1710),
.B(n_1613),
.Y(n_2456)
);

AOI21x1_ASAP7_75t_L g2457 ( 
.A1(n_2128),
.A2(n_1488),
.B(n_1484),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2099),
.Y(n_2458)
);

OAI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2169),
.A2(n_1710),
.B(n_1508),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2137),
.Y(n_2460)
);

AOI21x1_ASAP7_75t_L g2461 ( 
.A1(n_2140),
.A2(n_1508),
.B(n_1495),
.Y(n_2461)
);

CKINVDCx8_ASAP7_75t_R g2462 ( 
.A(n_2104),
.Y(n_2462)
);

AOI21xp33_ASAP7_75t_L g2463 ( 
.A1(n_2148),
.A2(n_809),
.B(n_807),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2071),
.A2(n_1798),
.B(n_1739),
.Y(n_2464)
);

OAI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2169),
.A2(n_1509),
.B(n_1495),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2141),
.B(n_1509),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2146),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2071),
.A2(n_1739),
.B(n_1533),
.Y(n_2468)
);

OAI21xp5_ASAP7_75t_SL g2469 ( 
.A1(n_2042),
.A2(n_809),
.B(n_807),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2151),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2178),
.B(n_1521),
.Y(n_2471)
);

OAI21x1_ASAP7_75t_L g2472 ( 
.A1(n_2225),
.A2(n_2228),
.B(n_2227),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2129),
.Y(n_2473)
);

OAI21x1_ASAP7_75t_L g2474 ( 
.A1(n_2230),
.A2(n_1538),
.B(n_1521),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2231),
.Y(n_2475)
);

OAI21x1_ASAP7_75t_L g2476 ( 
.A1(n_2139),
.A2(n_1539),
.B(n_1538),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2179),
.B(n_1539),
.Y(n_2477)
);

OAI21x1_ASAP7_75t_L g2478 ( 
.A1(n_2139),
.A2(n_1546),
.B(n_1545),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2184),
.B(n_1545),
.Y(n_2479)
);

OAI21xp5_ASAP7_75t_L g2480 ( 
.A1(n_2224),
.A2(n_1572),
.B(n_1546),
.Y(n_2480)
);

OAI21x1_ASAP7_75t_L g2481 ( 
.A1(n_2197),
.A2(n_1572),
.B(n_1316),
.Y(n_2481)
);

OAI21x1_ASAP7_75t_L g2482 ( 
.A1(n_2197),
.A2(n_1318),
.B(n_1311),
.Y(n_2482)
);

NAND3xp33_ASAP7_75t_L g2483 ( 
.A(n_2149),
.B(n_662),
.C(n_661),
.Y(n_2483)
);

INVxp67_ASAP7_75t_L g2484 ( 
.A(n_2082),
.Y(n_2484)
);

NAND2x1_ASAP7_75t_L g2485 ( 
.A(n_2124),
.B(n_1739),
.Y(n_2485)
);

AOI21xp5_ASAP7_75t_SL g2486 ( 
.A1(n_2124),
.A2(n_1668),
.B(n_1617),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_L g2487 ( 
.A1(n_2202),
.A2(n_2242),
.B(n_2226),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2186),
.Y(n_2488)
);

OA22x2_ASAP7_75t_L g2489 ( 
.A1(n_2162),
.A2(n_2121),
.B1(n_2082),
.B2(n_2201),
.Y(n_2489)
);

NAND3xp33_ASAP7_75t_L g2490 ( 
.A(n_2149),
.B(n_2119),
.C(n_2170),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2164),
.B(n_663),
.Y(n_2491)
);

AND2x2_ASAP7_75t_SL g2492 ( 
.A(n_2102),
.B(n_810),
.Y(n_2492)
);

OA21x2_ASAP7_75t_L g2493 ( 
.A1(n_2233),
.A2(n_1322),
.B(n_1318),
.Y(n_2493)
);

OAI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2237),
.A2(n_1520),
.B(n_1067),
.Y(n_2494)
);

NAND2x1p5_ASAP7_75t_L g2495 ( 
.A(n_2142),
.B(n_2173),
.Y(n_2495)
);

AOI21x1_ASAP7_75t_SL g2496 ( 
.A1(n_2163),
.A2(n_1668),
.B(n_1617),
.Y(n_2496)
);

AOI21xp33_ASAP7_75t_L g2497 ( 
.A1(n_2189),
.A2(n_812),
.B(n_810),
.Y(n_2497)
);

NAND3xp33_ASAP7_75t_SL g2498 ( 
.A(n_2160),
.B(n_666),
.C(n_665),
.Y(n_2498)
);

INVx2_ASAP7_75t_SL g2499 ( 
.A(n_2047),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2202),
.A2(n_2242),
.B(n_2226),
.Y(n_2500)
);

OAI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2247),
.A2(n_1520),
.B(n_1067),
.Y(n_2501)
);

AOI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2118),
.A2(n_667),
.B1(n_683),
.B2(n_680),
.Y(n_2502)
);

NAND2x1p5_ASAP7_75t_L g2503 ( 
.A(n_2142),
.B(n_1152),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2172),
.B(n_684),
.Y(n_2504)
);

BUFx6f_ASAP7_75t_L g2505 ( 
.A(n_2129),
.Y(n_2505)
);

OAI21xp5_ASAP7_75t_L g2506 ( 
.A1(n_2238),
.A2(n_1520),
.B(n_1067),
.Y(n_2506)
);

INVx1_ASAP7_75t_SL g2507 ( 
.A(n_2121),
.Y(n_2507)
);

INVx3_ASAP7_75t_L g2508 ( 
.A(n_2129),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2198),
.Y(n_2509)
);

AO31x2_ASAP7_75t_L g2510 ( 
.A1(n_2244),
.A2(n_812),
.A3(n_816),
.B(n_905),
.Y(n_2510)
);

OAI21x1_ASAP7_75t_L g2511 ( 
.A1(n_2246),
.A2(n_1068),
.B(n_1064),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2163),
.B(n_1668),
.Y(n_2512)
);

OAI21x1_ASAP7_75t_L g2513 ( 
.A1(n_2265),
.A2(n_1068),
.B(n_1064),
.Y(n_2513)
);

AOI21xp5_ASAP7_75t_L g2514 ( 
.A1(n_2243),
.A2(n_1494),
.B(n_1347),
.Y(n_2514)
);

OAI21x1_ASAP7_75t_L g2515 ( 
.A1(n_2265),
.A2(n_1069),
.B(n_1068),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2243),
.A2(n_1494),
.B(n_1347),
.Y(n_2516)
);

OAI22x1_ASAP7_75t_L g2517 ( 
.A1(n_2152),
.A2(n_816),
.B1(n_689),
.B2(n_692),
.Y(n_2517)
);

AOI221xp5_ASAP7_75t_L g2518 ( 
.A1(n_2135),
.A2(n_696),
.B1(n_701),
.B2(n_695),
.C(n_688),
.Y(n_2518)
);

OAI21x1_ASAP7_75t_L g2519 ( 
.A1(n_2239),
.A2(n_1069),
.B(n_968),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2188),
.B(n_702),
.Y(n_2520)
);

AOI21x1_ASAP7_75t_L g2521 ( 
.A1(n_2218),
.A2(n_928),
.B(n_927),
.Y(n_2521)
);

OAI21x1_ASAP7_75t_L g2522 ( 
.A1(n_2196),
.A2(n_1069),
.B(n_968),
.Y(n_2522)
);

BUFx6f_ASAP7_75t_L g2523 ( 
.A(n_2129),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2268),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2152),
.B(n_705),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2268),
.Y(n_2526)
);

AOI21xp5_ASAP7_75t_L g2527 ( 
.A1(n_2173),
.A2(n_1494),
.B(n_1347),
.Y(n_2527)
);

AOI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_2089),
.A2(n_2115),
.B(n_2158),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2193),
.Y(n_2529)
);

AND2x6_ASAP7_75t_L g2530 ( 
.A(n_2158),
.B(n_775),
.Y(n_2530)
);

OAI21x1_ASAP7_75t_L g2531 ( 
.A1(n_2263),
.A2(n_834),
.B(n_830),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2193),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2094),
.Y(n_2533)
);

NAND2x1p5_ASAP7_75t_L g2534 ( 
.A(n_2158),
.B(n_1169),
.Y(n_2534)
);

AO21x2_ASAP7_75t_L g2535 ( 
.A1(n_2160),
.A2(n_933),
.B(n_928),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2193),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2188),
.B(n_907),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2505),
.Y(n_2538)
);

INVx3_ASAP7_75t_SL g2539 ( 
.A(n_2375),
.Y(n_2539)
);

OAI22xp33_ASAP7_75t_SL g2540 ( 
.A1(n_2287),
.A2(n_706),
.B1(n_711),
.B2(n_707),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2347),
.B(n_2038),
.Y(n_2541)
);

INVx2_ASAP7_75t_SL g2542 ( 
.A(n_2454),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2312),
.B(n_2038),
.Y(n_2543)
);

CKINVDCx8_ASAP7_75t_R g2544 ( 
.A(n_2271),
.Y(n_2544)
);

OAI22xp33_ASAP7_75t_L g2545 ( 
.A1(n_2291),
.A2(n_2115),
.B1(n_2089),
.B2(n_715),
.Y(n_2545)
);

INVx2_ASAP7_75t_SL g2546 ( 
.A(n_2433),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2302),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2310),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2444),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2335),
.B(n_2061),
.Y(n_2550)
);

INVx1_ASAP7_75t_SL g2551 ( 
.A(n_2397),
.Y(n_2551)
);

BUFx3_ASAP7_75t_L g2552 ( 
.A(n_2434),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2300),
.B(n_2061),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2407),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2357),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2353),
.B(n_2135),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2368),
.B(n_2147),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2309),
.Y(n_2558)
);

BUFx2_ASAP7_75t_L g2559 ( 
.A(n_2415),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2396),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2397),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2407),
.Y(n_2562)
);

INVx3_ASAP7_75t_L g2563 ( 
.A(n_2505),
.Y(n_2563)
);

AND2x4_ASAP7_75t_L g2564 ( 
.A(n_2528),
.B(n_2089),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2505),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2433),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2426),
.Y(n_2567)
);

INVx3_ASAP7_75t_SL g2568 ( 
.A(n_2492),
.Y(n_2568)
);

OR2x6_ASAP7_75t_L g2569 ( 
.A(n_2317),
.B(n_2097),
.Y(n_2569)
);

INVx3_ASAP7_75t_L g2570 ( 
.A(n_2523),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2523),
.Y(n_2571)
);

AOI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2299),
.A2(n_2167),
.B(n_2158),
.Y(n_2572)
);

AND2x4_ASAP7_75t_L g2573 ( 
.A(n_2507),
.B(n_2115),
.Y(n_2573)
);

INVxp67_ASAP7_75t_SL g2574 ( 
.A(n_2295),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2523),
.Y(n_2575)
);

AOI21x1_ASAP7_75t_L g2576 ( 
.A1(n_2395),
.A2(n_936),
.B(n_933),
.Y(n_2576)
);

AOI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2490),
.A2(n_2147),
.B1(n_2109),
.B2(n_2092),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_2389),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2299),
.A2(n_2174),
.B(n_2167),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2462),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2284),
.Y(n_2581)
);

BUFx4_ASAP7_75t_SL g2582 ( 
.A(n_2325),
.Y(n_2582)
);

BUFx3_ASAP7_75t_L g2583 ( 
.A(n_2363),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2286),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2475),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2321),
.Y(n_2586)
);

BUFx2_ASAP7_75t_L g2587 ( 
.A(n_2329),
.Y(n_2587)
);

OAI221xp5_ASAP7_75t_L g2588 ( 
.A1(n_2400),
.A2(n_2278),
.B1(n_2469),
.B2(n_2463),
.C(n_2436),
.Y(n_2588)
);

AOI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2307),
.A2(n_2174),
.B(n_2167),
.Y(n_2589)
);

HB1xp67_ASAP7_75t_L g2590 ( 
.A(n_2392),
.Y(n_2590)
);

CKINVDCx6p67_ASAP7_75t_R g2591 ( 
.A(n_2389),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2334),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2399),
.B(n_2104),
.Y(n_2593)
);

INVx5_ASAP7_75t_L g2594 ( 
.A(n_2530),
.Y(n_2594)
);

AND2x4_ASAP7_75t_L g2595 ( 
.A(n_2507),
.B(n_2292),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2339),
.Y(n_2596)
);

OAI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2298),
.A2(n_2109),
.B1(n_2165),
.B2(n_2248),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2396),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2351),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2389),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2363),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2499),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2281),
.B(n_2193),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2389),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_2392),
.Y(n_2605)
);

AOI21xp33_ASAP7_75t_L g2606 ( 
.A1(n_2297),
.A2(n_2253),
.B(n_2252),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2293),
.A2(n_2315),
.B(n_2336),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_2315),
.A2(n_2174),
.B(n_2167),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2359),
.Y(n_2609)
);

INVxp67_ASAP7_75t_L g2610 ( 
.A(n_2290),
.Y(n_2610)
);

AOI21xp33_ASAP7_75t_L g2611 ( 
.A1(n_2297),
.A2(n_2253),
.B(n_2252),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2396),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2292),
.B(n_2050),
.Y(n_2613)
);

O2A1O1Ixp33_ASAP7_75t_L g2614 ( 
.A1(n_2463),
.A2(n_940),
.B(n_943),
.C(n_936),
.Y(n_2614)
);

AND2x4_ASAP7_75t_L g2615 ( 
.A(n_2318),
.B(n_2050),
.Y(n_2615)
);

AO21x2_ASAP7_75t_L g2616 ( 
.A1(n_2374),
.A2(n_2275),
.B(n_2282),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2360),
.Y(n_2617)
);

HB1xp67_ASAP7_75t_L g2618 ( 
.A(n_2392),
.Y(n_2618)
);

HB1xp67_ASAP7_75t_L g2619 ( 
.A(n_2328),
.Y(n_2619)
);

CKINVDCx20_ASAP7_75t_R g2620 ( 
.A(n_2439),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2366),
.Y(n_2621)
);

BUFx3_ASAP7_75t_L g2622 ( 
.A(n_2533),
.Y(n_2622)
);

INVx5_ASAP7_75t_L g2623 ( 
.A(n_2530),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2318),
.B(n_2337),
.Y(n_2624)
);

BUFx3_ASAP7_75t_L g2625 ( 
.A(n_2445),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2373),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2393),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2432),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2441),
.Y(n_2629)
);

BUFx3_ASAP7_75t_L g2630 ( 
.A(n_2445),
.Y(n_2630)
);

BUFx6f_ASAP7_75t_L g2631 ( 
.A(n_2337),
.Y(n_2631)
);

OAI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2383),
.A2(n_2084),
.B1(n_2078),
.B2(n_2097),
.Y(n_2632)
);

INVx2_ASAP7_75t_SL g2633 ( 
.A(n_2276),
.Y(n_2633)
);

INVx1_ASAP7_75t_SL g2634 ( 
.A(n_2276),
.Y(n_2634)
);

AND2x4_ASAP7_75t_L g2635 ( 
.A(n_2341),
.B(n_2078),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2450),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_2373),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_2439),
.Y(n_2638)
);

INVx2_ASAP7_75t_SL g2639 ( 
.A(n_2424),
.Y(n_2639)
);

BUFx8_ASAP7_75t_SL g2640 ( 
.A(n_2520),
.Y(n_2640)
);

BUFx6f_ASAP7_75t_L g2641 ( 
.A(n_2341),
.Y(n_2641)
);

AOI21xp5_ASAP7_75t_L g2642 ( 
.A1(n_2280),
.A2(n_2174),
.B(n_2253),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2355),
.B(n_2084),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2355),
.B(n_2270),
.Y(n_2644)
);

INVx3_ASAP7_75t_L g2645 ( 
.A(n_2382),
.Y(n_2645)
);

INVx4_ASAP7_75t_L g2646 ( 
.A(n_2382),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2344),
.B(n_2253),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2440),
.Y(n_2648)
);

INVx5_ASAP7_75t_L g2649 ( 
.A(n_2530),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2326),
.B(n_2199),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2460),
.Y(n_2651)
);

INVx3_ASAP7_75t_L g2652 ( 
.A(n_2386),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_2380),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2484),
.B(n_2097),
.Y(n_2654)
);

OAI222xp33_ASAP7_75t_L g2655 ( 
.A1(n_2287),
.A2(n_719),
.B1(n_716),
.B2(n_723),
.C1(n_720),
.C2(n_717),
.Y(n_2655)
);

BUFx4f_ASAP7_75t_L g2656 ( 
.A(n_2530),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2380),
.B(n_2270),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2532),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2440),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2440),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2467),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2470),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2488),
.Y(n_2663)
);

BUFx3_ASAP7_75t_L g2664 ( 
.A(n_2448),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_2448),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2509),
.Y(n_2666)
);

INVx2_ASAP7_75t_SL g2667 ( 
.A(n_2458),
.Y(n_2667)
);

CKINVDCx20_ASAP7_75t_R g2668 ( 
.A(n_2502),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2272),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2411),
.Y(n_2670)
);

OAI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2291),
.A2(n_732),
.B1(n_735),
.B2(n_734),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2411),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2510),
.Y(n_2673)
);

OAI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2305),
.A2(n_2199),
.B1(n_2212),
.B2(n_2208),
.Y(n_2674)
);

NOR2x1_ASAP7_75t_L g2675 ( 
.A(n_2535),
.B(n_940),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2510),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2458),
.Y(n_2677)
);

CKINVDCx5p33_ASAP7_75t_R g2678 ( 
.A(n_2504),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_SL g2679 ( 
.A(n_2414),
.B(n_2183),
.Y(n_2679)
);

AND2x4_ASAP7_75t_L g2680 ( 
.A(n_2473),
.B(n_2235),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2436),
.A2(n_705),
.B1(n_739),
.B2(n_737),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_2489),
.Y(n_2682)
);

AND2x4_ASAP7_75t_L g2683 ( 
.A(n_2473),
.B(n_2199),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_SL g2684 ( 
.A1(n_2273),
.A2(n_705),
.B1(n_742),
.B2(n_741),
.Y(n_2684)
);

BUFx12f_ASAP7_75t_L g2685 ( 
.A(n_2386),
.Y(n_2685)
);

OR2x6_ASAP7_75t_L g2686 ( 
.A(n_2303),
.B(n_775),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2510),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2273),
.B(n_747),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2508),
.Y(n_2689)
);

OR2x2_ASAP7_75t_SL g2690 ( 
.A(n_2483),
.B(n_775),
.Y(n_2690)
);

HB1xp67_ASAP7_75t_L g2691 ( 
.A(n_2295),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2508),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2378),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2352),
.Y(n_2694)
);

OR2x6_ASAP7_75t_L g2695 ( 
.A(n_2391),
.B(n_2092),
.Y(n_2695)
);

OR2x2_ASAP7_75t_L g2696 ( 
.A(n_2314),
.B(n_943),
.Y(n_2696)
);

INVx3_ASAP7_75t_SL g2697 ( 
.A(n_2489),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2277),
.B(n_749),
.Y(n_2698)
);

INVx1_ASAP7_75t_SL g2699 ( 
.A(n_2491),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2449),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_2524),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2449),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2472),
.Y(n_2703)
);

INVx3_ASAP7_75t_L g2704 ( 
.A(n_2342),
.Y(n_2704)
);

INVx1_ASAP7_75t_SL g2705 ( 
.A(n_2526),
.Y(n_2705)
);

O2A1O1Ixp33_ASAP7_75t_L g2706 ( 
.A1(n_2406),
.A2(n_948),
.B(n_950),
.C(n_944),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2306),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2446),
.B(n_553),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2529),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2422),
.Y(n_2710)
);

BUFx6f_ASAP7_75t_L g2711 ( 
.A(n_2342),
.Y(n_2711)
);

BUFx12f_ASAP7_75t_L g2712 ( 
.A(n_2495),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2536),
.B(n_377),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2364),
.B(n_553),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2525),
.A2(n_755),
.B1(n_760),
.B2(n_750),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_2330),
.Y(n_2716)
);

BUFx2_ASAP7_75t_L g2717 ( 
.A(n_2495),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2277),
.B(n_767),
.Y(n_2718)
);

BUFx2_ASAP7_75t_L g2719 ( 
.A(n_2296),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2296),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2283),
.A2(n_1177),
.B(n_1169),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2422),
.Y(n_2722)
);

CKINVDCx11_ASAP7_75t_R g2723 ( 
.A(n_2387),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2314),
.B(n_770),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_2512),
.B(n_382),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2537),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_L g2727 ( 
.A(n_2485),
.Y(n_2727)
);

BUFx2_ASAP7_75t_L g2728 ( 
.A(n_2412),
.Y(n_2728)
);

AOI21xp5_ASAP7_75t_L g2729 ( 
.A1(n_2348),
.A2(n_1177),
.B(n_1169),
.Y(n_2729)
);

INVx5_ASAP7_75t_L g2730 ( 
.A(n_2332),
.Y(n_2730)
);

OR2x6_ASAP7_75t_L g2731 ( 
.A(n_2356),
.B(n_2361),
.Y(n_2731)
);

NAND2x1p5_ASAP7_75t_L g2732 ( 
.A(n_2343),
.B(n_1169),
.Y(n_2732)
);

BUFx12f_ASAP7_75t_L g2733 ( 
.A(n_2365),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2313),
.Y(n_2734)
);

CKINVDCx20_ASAP7_75t_R g2735 ( 
.A(n_2405),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2431),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2431),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2305),
.A2(n_780),
.B1(n_781),
.B2(n_778),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2308),
.B(n_2279),
.Y(n_2739)
);

BUFx2_ASAP7_75t_R g2740 ( 
.A(n_2308),
.Y(n_2740)
);

O2A1O1Ixp33_ASAP7_75t_SL g2741 ( 
.A1(n_2274),
.A2(n_948),
.B(n_950),
.C(n_944),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2376),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2493),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2493),
.Y(n_2744)
);

INVx3_ASAP7_75t_L g2745 ( 
.A(n_2487),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_SL g2746 ( 
.A(n_2279),
.B(n_2065),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2289),
.Y(n_2747)
);

AOI22xp33_ASAP7_75t_L g2748 ( 
.A1(n_2338),
.A2(n_785),
.B1(n_791),
.B2(n_782),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2385),
.Y(n_2749)
);

BUFx6f_ASAP7_75t_L g2750 ( 
.A(n_2534),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2338),
.A2(n_797),
.B1(n_798),
.B2(n_793),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_2319),
.A2(n_801),
.B1(n_802),
.B2(n_800),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2412),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2403),
.B(n_808),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2500),
.B(n_383),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2371),
.B(n_813),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2534),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2404),
.B(n_814),
.Y(n_2758)
);

BUFx6f_ASAP7_75t_L g2759 ( 
.A(n_2537),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2288),
.B(n_2370),
.Y(n_2760)
);

NOR2xp67_ASAP7_75t_L g2761 ( 
.A(n_2498),
.B(n_2065),
.Y(n_2761)
);

BUFx2_ASAP7_75t_L g2762 ( 
.A(n_2442),
.Y(n_2762)
);

BUFx12f_ASAP7_75t_L g2763 ( 
.A(n_2503),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2503),
.Y(n_2764)
);

INVx6_ASAP7_75t_L g2765 ( 
.A(n_2496),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2517),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2304),
.Y(n_2767)
);

CKINVDCx8_ASAP7_75t_R g2768 ( 
.A(n_2453),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2519),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2442),
.B(n_815),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2466),
.Y(n_2771)
);

AOI21xp5_ASAP7_75t_L g2772 ( 
.A1(n_2348),
.A2(n_1177),
.B(n_1169),
.Y(n_2772)
);

INVx2_ASAP7_75t_SL g2773 ( 
.A(n_2340),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2466),
.Y(n_2774)
);

INVx5_ASAP7_75t_L g2775 ( 
.A(n_2535),
.Y(n_2775)
);

AOI21xp5_ASAP7_75t_L g2776 ( 
.A1(n_2320),
.A2(n_1185),
.B(n_1177),
.Y(n_2776)
);

NAND2x1p5_ASAP7_75t_L g2777 ( 
.A(n_2333),
.B(n_1177),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2471),
.Y(n_2778)
);

NAND3xp33_ASAP7_75t_L g2779 ( 
.A(n_2408),
.B(n_952),
.C(n_951),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2358),
.Y(n_2780)
);

AND2x2_ASAP7_75t_SL g2781 ( 
.A(n_2288),
.B(n_951),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2294),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2531),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2471),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2390),
.B(n_952),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_SL g2786 ( 
.A(n_2394),
.B(n_954),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2377),
.Y(n_2787)
);

BUFx6f_ASAP7_75t_L g2788 ( 
.A(n_2354),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2390),
.B(n_954),
.Y(n_2789)
);

INVx2_ASAP7_75t_SL g2790 ( 
.A(n_2477),
.Y(n_2790)
);

INVx5_ASAP7_75t_L g2791 ( 
.A(n_2349),
.Y(n_2791)
);

AOI21x1_ASAP7_75t_L g2792 ( 
.A1(n_2461),
.A2(n_908),
.B(n_907),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2477),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2401),
.B(n_389),
.Y(n_2794)
);

BUFx3_ASAP7_75t_L g2795 ( 
.A(n_2362),
.Y(n_2795)
);

AND2x4_ASAP7_75t_L g2796 ( 
.A(n_2427),
.B(n_390),
.Y(n_2796)
);

OAI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2322),
.A2(n_1188),
.B1(n_1210),
.B2(n_1185),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2684),
.A2(n_2301),
.B1(n_2438),
.B2(n_2413),
.Y(n_2798)
);

OAI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_2688),
.A2(n_2684),
.B(n_2588),
.Y(n_2799)
);

AOI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2588),
.A2(n_2301),
.B1(n_2451),
.B2(n_2428),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2671),
.A2(n_2497),
.B1(n_2323),
.B2(n_2346),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2671),
.A2(n_2497),
.B1(n_2323),
.B2(n_2518),
.Y(n_2802)
);

AO31x2_ASAP7_75t_L g2803 ( 
.A1(n_2648),
.A2(n_2447),
.A3(n_2430),
.B(n_2416),
.Y(n_2803)
);

AND2x4_ASAP7_75t_L g2804 ( 
.A(n_2573),
.B(n_2367),
.Y(n_2804)
);

OAI21x1_ASAP7_75t_L g2805 ( 
.A1(n_2721),
.A2(n_2316),
.B(n_2452),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2607),
.A2(n_2374),
.B(n_2369),
.Y(n_2806)
);

NAND2x1p5_ASAP7_75t_L g2807 ( 
.A(n_2594),
.B(n_2331),
.Y(n_2807)
);

OAI21x1_ASAP7_75t_L g2808 ( 
.A1(n_2721),
.A2(n_2457),
.B(n_2327),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2554),
.B(n_2402),
.Y(n_2809)
);

INVx1_ASAP7_75t_SL g2810 ( 
.A(n_2620),
.Y(n_2810)
);

OAI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2655),
.A2(n_2465),
.B(n_2345),
.Y(n_2811)
);

AND2x4_ASAP7_75t_L g2812 ( 
.A(n_2573),
.B(n_2367),
.Y(n_2812)
);

AND2x4_ASAP7_75t_L g2813 ( 
.A(n_2552),
.B(n_2367),
.Y(n_2813)
);

OA21x2_ASAP7_75t_L g2814 ( 
.A1(n_2776),
.A2(n_2311),
.B(n_2416),
.Y(n_2814)
);

OA21x2_ASAP7_75t_L g2815 ( 
.A1(n_2776),
.A2(n_2772),
.B(n_2729),
.Y(n_2815)
);

OR2x6_ASAP7_75t_L g2816 ( 
.A(n_2607),
.B(n_2430),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2661),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2562),
.B(n_2402),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2553),
.B(n_2443),
.Y(n_2819)
);

OAI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2655),
.A2(n_2465),
.B(n_2311),
.Y(n_2820)
);

AO21x2_ASAP7_75t_L g2821 ( 
.A1(n_2673),
.A2(n_2443),
.B(n_2455),
.Y(n_2821)
);

OR2x2_ASAP7_75t_L g2822 ( 
.A(n_2762),
.B(n_2417),
.Y(n_2822)
);

INVx2_ASAP7_75t_SL g2823 ( 
.A(n_2549),
.Y(n_2823)
);

OAI21x1_ASAP7_75t_L g2824 ( 
.A1(n_2576),
.A2(n_2324),
.B(n_2522),
.Y(n_2824)
);

BUFx2_ASAP7_75t_SL g2825 ( 
.A(n_2620),
.Y(n_2825)
);

AO21x2_ASAP7_75t_L g2826 ( 
.A1(n_2676),
.A2(n_2456),
.B(n_2455),
.Y(n_2826)
);

OA21x2_ASAP7_75t_L g2827 ( 
.A1(n_2729),
.A2(n_2417),
.B(n_2456),
.Y(n_2827)
);

AND2x2_ASAP7_75t_SL g2828 ( 
.A(n_2656),
.B(n_2479),
.Y(n_2828)
);

INVx1_ASAP7_75t_SL g2829 ( 
.A(n_2561),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2661),
.Y(n_2830)
);

OR2x6_ASAP7_75t_L g2831 ( 
.A(n_2572),
.B(n_2486),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_L g2832 ( 
.A1(n_2681),
.A2(n_2540),
.B1(n_2781),
.B2(n_2751),
.Y(n_2832)
);

A2O1A1Ixp33_ASAP7_75t_L g2833 ( 
.A1(n_2656),
.A2(n_2468),
.B(n_2501),
.C(n_2494),
.Y(n_2833)
);

CKINVDCx8_ASAP7_75t_R g2834 ( 
.A(n_2678),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2662),
.Y(n_2835)
);

OA21x2_ASAP7_75t_L g2836 ( 
.A1(n_2772),
.A2(n_2421),
.B(n_2420),
.Y(n_2836)
);

AOI22x1_ASAP7_75t_L g2837 ( 
.A1(n_2568),
.A2(n_2459),
.B1(n_2418),
.B2(n_2398),
.Y(n_2837)
);

OAI21x1_ASAP7_75t_L g2838 ( 
.A1(n_2792),
.A2(n_2642),
.B(n_2732),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2760),
.B(n_2285),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2662),
.Y(n_2840)
);

A2O1A1Ixp33_ASAP7_75t_L g2841 ( 
.A1(n_2781),
.A2(n_2501),
.B(n_2494),
.C(n_2459),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2582),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_SL g2843 ( 
.A(n_2740),
.B(n_2437),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2663),
.Y(n_2844)
);

AOI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2746),
.A2(n_2447),
.B1(n_2479),
.B2(n_2372),
.Y(n_2845)
);

INVx3_ASAP7_75t_L g2846 ( 
.A(n_2709),
.Y(n_2846)
);

OAI21x1_ASAP7_75t_L g2847 ( 
.A1(n_2642),
.A2(n_2515),
.B(n_2513),
.Y(n_2847)
);

OAI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2732),
.A2(n_2425),
.B(n_2384),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2543),
.B(n_2285),
.Y(n_2849)
);

BUFx12f_ASAP7_75t_L g2850 ( 
.A(n_2723),
.Y(n_2850)
);

BUFx6f_ASAP7_75t_L g2851 ( 
.A(n_2578),
.Y(n_2851)
);

OAI21x1_ASAP7_75t_L g2852 ( 
.A1(n_2572),
.A2(n_2511),
.B(n_2482),
.Y(n_2852)
);

O2A1O1Ixp33_ASAP7_75t_SL g2853 ( 
.A1(n_2545),
.A2(n_2388),
.B(n_2381),
.C(n_2419),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_2723),
.Y(n_2854)
);

CKINVDCx6p67_ASAP7_75t_R g2855 ( 
.A(n_2539),
.Y(n_2855)
);

INVx4_ASAP7_75t_L g2856 ( 
.A(n_2578),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2663),
.Y(n_2857)
);

AND2x6_ASAP7_75t_L g2858 ( 
.A(n_2564),
.B(n_2423),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2739),
.B(n_2521),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2579),
.A2(n_2481),
.B(n_2480),
.Y(n_2860)
);

OAI21x1_ASAP7_75t_L g2861 ( 
.A1(n_2579),
.A2(n_2480),
.B(n_2478),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2581),
.Y(n_2862)
);

OAI21x1_ASAP7_75t_SL g2863 ( 
.A1(n_2589),
.A2(n_2464),
.B(n_2379),
.Y(n_2863)
);

OAI21x1_ASAP7_75t_L g2864 ( 
.A1(n_2648),
.A2(n_2476),
.B(n_2435),
.Y(n_2864)
);

BUFx6f_ASAP7_75t_L g2865 ( 
.A(n_2578),
.Y(n_2865)
);

NAND3xp33_ASAP7_75t_L g2866 ( 
.A(n_2748),
.B(n_909),
.C(n_908),
.Y(n_2866)
);

CKINVDCx20_ASAP7_75t_R g2867 ( 
.A(n_2640),
.Y(n_2867)
);

O2A1O1Ixp33_ASAP7_75t_SL g2868 ( 
.A1(n_2545),
.A2(n_2350),
.B(n_2506),
.C(n_2514),
.Y(n_2868)
);

AO21x2_ASAP7_75t_L g2869 ( 
.A1(n_2687),
.A2(n_2506),
.B(n_2474),
.Y(n_2869)
);

BUFx12f_ASAP7_75t_L g2870 ( 
.A(n_2542),
.Y(n_2870)
);

OAI21x1_ASAP7_75t_L g2871 ( 
.A1(n_2659),
.A2(n_2429),
.B(n_2410),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2584),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2586),
.Y(n_2873)
);

AOI22xp33_ASAP7_75t_L g2874 ( 
.A1(n_2681),
.A2(n_2409),
.B1(n_834),
.B2(n_838),
.Y(n_2874)
);

AOI222xp33_ASAP7_75t_L g2875 ( 
.A1(n_2748),
.A2(n_838),
.B1(n_830),
.B2(n_3),
.C1(n_8),
.C2(n_1),
.Y(n_2875)
);

INVx2_ASAP7_75t_SL g2876 ( 
.A(n_2549),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2694),
.B(n_2285),
.Y(n_2877)
);

OAI21x1_ASAP7_75t_L g2878 ( 
.A1(n_2659),
.A2(n_2527),
.B(n_2516),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2592),
.Y(n_2879)
);

AO31x2_ASAP7_75t_L g2880 ( 
.A1(n_2660),
.A2(n_911),
.A3(n_912),
.B(n_909),
.Y(n_2880)
);

OA21x2_ASAP7_75t_L g2881 ( 
.A1(n_2560),
.A2(n_912),
.B(n_911),
.Y(n_2881)
);

NOR2x1_ASAP7_75t_R g2882 ( 
.A(n_2716),
.B(n_914),
.Y(n_2882)
);

HB1xp67_ASAP7_75t_L g2883 ( 
.A(n_2619),
.Y(n_2883)
);

OAI21x1_ASAP7_75t_L g2884 ( 
.A1(n_2660),
.A2(n_917),
.B(n_914),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2759),
.B(n_917),
.Y(n_2885)
);

AOI22xp33_ASAP7_75t_L g2886 ( 
.A1(n_2751),
.A2(n_918),
.B1(n_6),
.B2(n_2),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2596),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2609),
.Y(n_2888)
);

AND2x4_ASAP7_75t_L g2889 ( 
.A(n_2552),
.B(n_392),
.Y(n_2889)
);

INVx2_ASAP7_75t_SL g2890 ( 
.A(n_2622),
.Y(n_2890)
);

OAI21x1_ASAP7_75t_L g2891 ( 
.A1(n_2560),
.A2(n_918),
.B(n_977),
.Y(n_2891)
);

AOI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2668),
.A2(n_1520),
.B1(n_985),
.B2(n_977),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2617),
.Y(n_2893)
);

BUFx3_ASAP7_75t_L g2894 ( 
.A(n_2685),
.Y(n_2894)
);

AOI22xp33_ASAP7_75t_SL g2895 ( 
.A1(n_2730),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_2895)
);

OAI21x1_ASAP7_75t_L g2896 ( 
.A1(n_2598),
.A2(n_985),
.B(n_977),
.Y(n_2896)
);

OAI21x1_ASAP7_75t_L g2897 ( 
.A1(n_2598),
.A2(n_985),
.B(n_977),
.Y(n_2897)
);

AOI22xp33_ASAP7_75t_L g2898 ( 
.A1(n_2668),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2898)
);

INVx1_ASAP7_75t_SL g2899 ( 
.A(n_2638),
.Y(n_2899)
);

BUFx2_ASAP7_75t_L g2900 ( 
.A(n_2733),
.Y(n_2900)
);

OAI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2679),
.A2(n_1520),
.B(n_985),
.Y(n_2901)
);

OAI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2679),
.A2(n_1520),
.B(n_398),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2621),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2650),
.B(n_9),
.Y(n_2904)
);

OAI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2738),
.A2(n_1520),
.B(n_399),
.Y(n_2905)
);

AO21x2_ASAP7_75t_L g2906 ( 
.A1(n_2612),
.A2(n_10),
.B(n_12),
.Y(n_2906)
);

OAI21x1_ASAP7_75t_L g2907 ( 
.A1(n_2612),
.A2(n_400),
.B(n_394),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2627),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_2582),
.Y(n_2909)
);

OAI21x1_ASAP7_75t_L g2910 ( 
.A1(n_2747),
.A2(n_407),
.B(n_403),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2628),
.Y(n_2911)
);

AO31x2_ASAP7_75t_L g2912 ( 
.A1(n_2743),
.A2(n_15),
.A3(n_12),
.B(n_13),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2768),
.A2(n_1188),
.B1(n_1210),
.B2(n_1185),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2741),
.A2(n_1188),
.B(n_1185),
.Y(n_2914)
);

AO31x2_ASAP7_75t_L g2915 ( 
.A1(n_2743),
.A2(n_17),
.A3(n_13),
.B(n_16),
.Y(n_2915)
);

OAI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2752),
.A2(n_410),
.B(n_409),
.Y(n_2916)
);

CKINVDCx5p33_ASAP7_75t_R g2917 ( 
.A(n_2539),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_L g2918 ( 
.A(n_2697),
.B(n_16),
.Y(n_2918)
);

AOI21x1_ASAP7_75t_L g2919 ( 
.A1(n_2786),
.A2(n_17),
.B(n_18),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2639),
.B(n_2670),
.Y(n_2920)
);

OAI22xp33_ASAP7_75t_SL g2921 ( 
.A1(n_2697),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2921)
);

AOI22xp33_ASAP7_75t_L g2922 ( 
.A1(n_2735),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2922)
);

OAI21x1_ASAP7_75t_L g2923 ( 
.A1(n_2747),
.A2(n_413),
.B(n_411),
.Y(n_2923)
);

AND2x4_ASAP7_75t_L g2924 ( 
.A(n_2555),
.B(n_2728),
.Y(n_2924)
);

AND2x4_ASAP7_75t_L g2925 ( 
.A(n_2555),
.B(n_415),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2629),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2636),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2651),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2753),
.B(n_22),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2568),
.A2(n_1188),
.B1(n_1210),
.B2(n_1185),
.Y(n_2930)
);

AOI21xp33_ASAP7_75t_L g2931 ( 
.A1(n_2724),
.A2(n_26),
.B(n_27),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2666),
.Y(n_2932)
);

OAI21x1_ASAP7_75t_L g2933 ( 
.A1(n_2767),
.A2(n_422),
.B(n_416),
.Y(n_2933)
);

OAI21x1_ASAP7_75t_L g2934 ( 
.A1(n_2767),
.A2(n_425),
.B(n_423),
.Y(n_2934)
);

AND2x4_ASAP7_75t_L g2935 ( 
.A(n_2564),
.B(n_426),
.Y(n_2935)
);

NAND2x1p5_ASAP7_75t_L g2936 ( 
.A(n_2594),
.B(n_995),
.Y(n_2936)
);

INVx3_ASAP7_75t_L g2937 ( 
.A(n_2709),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2595),
.B(n_2556),
.Y(n_2938)
);

AO21x2_ASAP7_75t_L g2939 ( 
.A1(n_2786),
.A2(n_2605),
.B(n_2590),
.Y(n_2939)
);

INVx3_ASAP7_75t_SL g2940 ( 
.A(n_2548),
.Y(n_2940)
);

AO21x2_ASAP7_75t_L g2941 ( 
.A1(n_2590),
.A2(n_26),
.B(n_27),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2595),
.B(n_2557),
.Y(n_2942)
);

OAI21x1_ASAP7_75t_L g2943 ( 
.A1(n_2782),
.A2(n_430),
.B(n_427),
.Y(n_2943)
);

OA21x2_ASAP7_75t_L g2944 ( 
.A1(n_2744),
.A2(n_30),
.B(n_31),
.Y(n_2944)
);

OAI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_2682),
.A2(n_1210),
.B1(n_1266),
.B2(n_1188),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2672),
.B(n_30),
.Y(n_2946)
);

OAI21x1_ASAP7_75t_L g2947 ( 
.A1(n_2782),
.A2(n_433),
.B(n_432),
.Y(n_2947)
);

AOI221xp5_ASAP7_75t_L g2948 ( 
.A1(n_2752),
.A2(n_35),
.B1(n_31),
.B2(n_33),
.C(n_36),
.Y(n_2948)
);

OAI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_2770),
.A2(n_435),
.B(n_434),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2669),
.Y(n_2950)
);

OAI21x1_ASAP7_75t_L g2951 ( 
.A1(n_2589),
.A2(n_437),
.B(n_436),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2599),
.Y(n_2952)
);

AOI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2735),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2700),
.Y(n_2954)
);

AO22x2_ASAP7_75t_L g2955 ( 
.A1(n_2574),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2702),
.Y(n_2956)
);

OAI21x1_ASAP7_75t_L g2957 ( 
.A1(n_2744),
.A2(n_441),
.B(n_440),
.Y(n_2957)
);

OAI21x1_ASAP7_75t_L g2958 ( 
.A1(n_2707),
.A2(n_443),
.B(n_442),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2710),
.Y(n_2959)
);

AO32x2_ASAP7_75t_L g2960 ( 
.A1(n_2790),
.A2(n_43),
.A3(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_2960)
);

OA21x2_ASAP7_75t_L g2961 ( 
.A1(n_2707),
.A2(n_2734),
.B(n_2618),
.Y(n_2961)
);

OAI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2770),
.A2(n_445),
.B(n_444),
.Y(n_2962)
);

AND2x4_ASAP7_75t_L g2963 ( 
.A(n_2610),
.B(n_2559),
.Y(n_2963)
);

OAI21x1_ASAP7_75t_L g2964 ( 
.A1(n_2734),
.A2(n_448),
.B(n_447),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2578),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2745),
.A2(n_450),
.B(n_449),
.Y(n_2966)
);

OAI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2698),
.A2(n_453),
.B(n_452),
.Y(n_2967)
);

AO21x1_ASAP7_75t_L g2968 ( 
.A1(n_2714),
.A2(n_42),
.B(n_44),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2722),
.Y(n_2969)
);

AOI22xp33_ASAP7_75t_L g2970 ( 
.A1(n_2766),
.A2(n_2773),
.B1(n_2749),
.B2(n_2730),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2736),
.Y(n_2971)
);

AOI21x1_ASAP7_75t_L g2972 ( 
.A1(n_2608),
.A2(n_45),
.B(n_46),
.Y(n_2972)
);

BUFx2_ASAP7_75t_L g2973 ( 
.A(n_2712),
.Y(n_2973)
);

HB1xp67_ASAP7_75t_L g2974 ( 
.A(n_2619),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2737),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2691),
.Y(n_2976)
);

CKINVDCx5p33_ASAP7_75t_R g2977 ( 
.A(n_2640),
.Y(n_2977)
);

OAI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2730),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_2978)
);

OAI21x1_ASAP7_75t_L g2979 ( 
.A1(n_2745),
.A2(n_456),
.B(n_454),
.Y(n_2979)
);

OAI21x1_ASAP7_75t_L g2980 ( 
.A1(n_2769),
.A2(n_458),
.B(n_457),
.Y(n_2980)
);

OAI22xp5_ASAP7_75t_L g2981 ( 
.A1(n_2577),
.A2(n_1266),
.B1(n_1296),
.B2(n_1210),
.Y(n_2981)
);

NAND2x1p5_ASAP7_75t_L g2982 ( 
.A(n_2594),
.B(n_995),
.Y(n_2982)
);

AOI22xp33_ASAP7_75t_SL g2983 ( 
.A1(n_2730),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2983)
);

OAI21x1_ASAP7_75t_L g2984 ( 
.A1(n_2769),
.A2(n_461),
.B(n_460),
.Y(n_2984)
);

OR2x2_ASAP7_75t_L g2985 ( 
.A(n_2691),
.B(n_49),
.Y(n_2985)
);

OAI21x1_ASAP7_75t_L g2986 ( 
.A1(n_2742),
.A2(n_464),
.B(n_463),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2541),
.B(n_50),
.Y(n_2987)
);

INVx2_ASAP7_75t_SL g2988 ( 
.A(n_2622),
.Y(n_2988)
);

AOI21xp33_ASAP7_75t_SL g2989 ( 
.A1(n_2718),
.A2(n_52),
.B(n_53),
.Y(n_2989)
);

OAI21x1_ASAP7_75t_L g2990 ( 
.A1(n_2742),
.A2(n_2780),
.B(n_2787),
.Y(n_2990)
);

OAI21x1_ASAP7_75t_SL g2991 ( 
.A1(n_2608),
.A2(n_52),
.B(n_54),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2574),
.B(n_54),
.Y(n_2992)
);

BUFx6f_ASAP7_75t_L g2993 ( 
.A(n_2600),
.Y(n_2993)
);

O2A1O1Ixp33_ASAP7_75t_SL g2994 ( 
.A1(n_2597),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2610),
.B(n_55),
.Y(n_2995)
);

AO21x2_ASAP7_75t_L g2996 ( 
.A1(n_2605),
.A2(n_2618),
.B(n_2616),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2696),
.B(n_56),
.Y(n_2997)
);

INVxp67_ASAP7_75t_L g2998 ( 
.A(n_2701),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2703),
.Y(n_2999)
);

AO21x1_ASAP7_75t_L g3000 ( 
.A1(n_2674),
.A2(n_58),
.B(n_59),
.Y(n_3000)
);

INVxp67_ASAP7_75t_SL g3001 ( 
.A(n_2693),
.Y(n_3001)
);

INVx3_ASAP7_75t_L g3002 ( 
.A(n_2653),
.Y(n_3002)
);

BUFx12f_ASAP7_75t_L g3003 ( 
.A(n_2546),
.Y(n_3003)
);

BUFx2_ASAP7_75t_L g3004 ( 
.A(n_2633),
.Y(n_3004)
);

AO32x2_ASAP7_75t_L g3005 ( 
.A1(n_2658),
.A2(n_63),
.A3(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_3005)
);

BUFx2_ASAP7_75t_L g3006 ( 
.A(n_2653),
.Y(n_3006)
);

AOI22xp5_ASAP7_75t_L g3007 ( 
.A1(n_2761),
.A2(n_2699),
.B1(n_2695),
.B2(n_2725),
.Y(n_3007)
);

OAI21x1_ASAP7_75t_L g3008 ( 
.A1(n_2780),
.A2(n_469),
.B(n_467),
.Y(n_3008)
);

NAND2x1p5_ASAP7_75t_L g3009 ( 
.A(n_2594),
.B(n_995),
.Y(n_3009)
);

OA21x2_ASAP7_75t_L g3010 ( 
.A1(n_2606),
.A2(n_61),
.B(n_63),
.Y(n_3010)
);

OAI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2777),
.A2(n_473),
.B(n_472),
.Y(n_3011)
);

OAI21x1_ASAP7_75t_L g3012 ( 
.A1(n_2777),
.A2(n_476),
.B(n_475),
.Y(n_3012)
);

OAI21x1_ASAP7_75t_SL g3013 ( 
.A1(n_2785),
.A2(n_65),
.B(n_67),
.Y(n_3013)
);

AO21x2_ASAP7_75t_L g3014 ( 
.A1(n_2616),
.A2(n_2611),
.B(n_2741),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2547),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2719),
.B(n_477),
.Y(n_3016)
);

BUFx4f_ASAP7_75t_SL g3017 ( 
.A(n_2580),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2558),
.Y(n_3018)
);

OAI21x1_ASAP7_75t_L g3019 ( 
.A1(n_2797),
.A2(n_482),
.B(n_478),
.Y(n_3019)
);

OAI21x1_ASAP7_75t_L g3020 ( 
.A1(n_2675),
.A2(n_485),
.B(n_483),
.Y(n_3020)
);

A2O1A1Ixp33_ASAP7_75t_L g3021 ( 
.A1(n_2623),
.A2(n_72),
.B(n_68),
.C(n_69),
.Y(n_3021)
);

O2A1O1Ixp33_ASAP7_75t_L g3022 ( 
.A1(n_2686),
.A2(n_74),
.B(n_69),
.C(n_73),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2585),
.Y(n_3023)
);

INVxp67_ASAP7_75t_L g3024 ( 
.A(n_2705),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_2799),
.A2(n_2686),
.B1(n_2708),
.B2(n_2779),
.Y(n_3025)
);

HB1xp67_ASAP7_75t_L g3026 ( 
.A(n_2883),
.Y(n_3026)
);

OAI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2798),
.A2(n_2800),
.B1(n_2820),
.B2(n_2811),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_2832),
.A2(n_2686),
.B1(n_2759),
.B2(n_2726),
.Y(n_3028)
);

OA21x2_ASAP7_75t_L g3029 ( 
.A1(n_2990),
.A2(n_2720),
.B(n_2717),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_3024),
.B(n_2551),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2872),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_2832),
.A2(n_2759),
.B1(n_2587),
.B2(n_2791),
.Y(n_3032)
);

AO31x2_ASAP7_75t_L g3033 ( 
.A1(n_2806),
.A2(n_2774),
.A3(n_2778),
.B(n_2771),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2872),
.Y(n_3034)
);

OAI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2802),
.A2(n_2690),
.B1(n_2649),
.B2(n_2623),
.Y(n_3035)
);

BUFx2_ASAP7_75t_L g3036 ( 
.A(n_2924),
.Y(n_3036)
);

AND2x4_ASAP7_75t_L g3037 ( 
.A(n_2813),
.B(n_2569),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2873),
.Y(n_3038)
);

AOI22xp33_ASAP7_75t_L g3039 ( 
.A1(n_2802),
.A2(n_2759),
.B1(n_2791),
.B2(n_2593),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2886),
.A2(n_2649),
.B1(n_2623),
.B2(n_2580),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_3024),
.B(n_2634),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2873),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2903),
.Y(n_3043)
);

AND2x4_ASAP7_75t_L g3044 ( 
.A(n_2813),
.B(n_2569),
.Y(n_3044)
);

OR2x2_ASAP7_75t_L g3045 ( 
.A(n_2822),
.B(n_2603),
.Y(n_3045)
);

O2A1O1Ixp33_ASAP7_75t_L g3046 ( 
.A1(n_3021),
.A2(n_2706),
.B(n_2758),
.C(n_2756),
.Y(n_3046)
);

AOI222xp33_ASAP7_75t_L g3047 ( 
.A1(n_2948),
.A2(n_2754),
.B1(n_2550),
.B2(n_2789),
.C1(n_2791),
.C2(n_2725),
.Y(n_3047)
);

BUFx2_ASAP7_75t_L g3048 ( 
.A(n_2924),
.Y(n_3048)
);

OAI22xp5_ASAP7_75t_L g3049 ( 
.A1(n_2886),
.A2(n_2623),
.B1(n_2649),
.B2(n_2569),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2903),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2908),
.Y(n_3051)
);

OAI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2898),
.A2(n_2649),
.B1(n_2544),
.B2(n_2695),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2908),
.Y(n_3053)
);

BUFx2_ASAP7_75t_L g3054 ( 
.A(n_3006),
.Y(n_3054)
);

AOI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2875),
.A2(n_2791),
.B1(n_2695),
.B2(n_2794),
.Y(n_3055)
);

OAI221xp5_ASAP7_75t_L g3056 ( 
.A1(n_2898),
.A2(n_2715),
.B1(n_2654),
.B2(n_2566),
.C(n_2567),
.Y(n_3056)
);

HB1xp67_ASAP7_75t_L g3057 ( 
.A(n_2883),
.Y(n_3057)
);

HB1xp67_ASAP7_75t_L g3058 ( 
.A(n_2974),
.Y(n_3058)
);

AO21x1_ASAP7_75t_L g3059 ( 
.A1(n_2918),
.A2(n_2647),
.B(n_2784),
.Y(n_3059)
);

AOI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_2948),
.A2(n_2794),
.B1(n_2796),
.B2(n_2583),
.Y(n_3060)
);

INVx1_ASAP7_75t_SL g3061 ( 
.A(n_2825),
.Y(n_3061)
);

HB1xp67_ASAP7_75t_L g3062 ( 
.A(n_2974),
.Y(n_3062)
);

INVx4_ASAP7_75t_L g3063 ( 
.A(n_2917),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_3007),
.A2(n_2796),
.B1(n_2632),
.B2(n_2755),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2922),
.A2(n_2583),
.B1(n_2795),
.B2(n_2755),
.Y(n_3065)
);

AOI21xp33_ASAP7_75t_L g3066 ( 
.A1(n_2978),
.A2(n_2916),
.B(n_2949),
.Y(n_3066)
);

AOI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_2801),
.A2(n_2601),
.B1(n_2795),
.B2(n_2731),
.Y(n_3067)
);

INVx4_ASAP7_75t_L g3068 ( 
.A(n_2917),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_2834),
.Y(n_3069)
);

OR2x2_ASAP7_75t_L g3070 ( 
.A(n_2976),
.B(n_2731),
.Y(n_3070)
);

INVx3_ASAP7_75t_L g3071 ( 
.A(n_2846),
.Y(n_3071)
);

OAI221xp5_ASAP7_75t_L g3072 ( 
.A1(n_2922),
.A2(n_2602),
.B1(n_2601),
.B2(n_2706),
.C(n_2731),
.Y(n_3072)
);

OAI222xp33_ASAP7_75t_L g3073 ( 
.A1(n_2895),
.A2(n_2793),
.B1(n_2775),
.B2(n_2704),
.C1(n_2630),
.C2(n_2625),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2926),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2926),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2851),
.Y(n_3076)
);

CKINVDCx6p67_ASAP7_75t_R g3077 ( 
.A(n_2940),
.Y(n_3077)
);

OAI21x1_ASAP7_75t_L g3078 ( 
.A1(n_2838),
.A2(n_2764),
.B(n_2704),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2932),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2932),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_SL g3081 ( 
.A1(n_2955),
.A2(n_2775),
.B1(n_2600),
.B2(n_2604),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2920),
.B(n_2624),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2950),
.B(n_2624),
.Y(n_3083)
);

INVx3_ASAP7_75t_L g3084 ( 
.A(n_2846),
.Y(n_3084)
);

AOI211xp5_ASAP7_75t_L g3085 ( 
.A1(n_2978),
.A2(n_2614),
.B(n_2713),
.C(n_2683),
.Y(n_3085)
);

OAI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_2843),
.A2(n_2816),
.B1(n_2918),
.B2(n_2962),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_2963),
.B(n_2625),
.Y(n_3087)
);

AO31x2_ASAP7_75t_L g3088 ( 
.A1(n_2806),
.A2(n_2775),
.A3(n_2646),
.B(n_2788),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2963),
.B(n_2630),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2862),
.Y(n_3090)
);

AOI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2953),
.A2(n_2801),
.B1(n_2931),
.B2(n_2895),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_L g3092 ( 
.A1(n_2953),
.A2(n_2713),
.B1(n_2775),
.B2(n_2783),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_2938),
.B(n_2664),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2879),
.Y(n_3094)
);

CKINVDCx11_ASAP7_75t_R g3095 ( 
.A(n_2867),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_SL g3096 ( 
.A(n_2828),
.B(n_2711),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2851),
.Y(n_3097)
);

BUFx2_ASAP7_75t_SL g3098 ( 
.A(n_2867),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2849),
.B(n_2692),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2942),
.B(n_2664),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2887),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2840),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2840),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_L g3104 ( 
.A(n_2992),
.B(n_2692),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2952),
.B(n_2631),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2857),
.Y(n_3106)
);

OAI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_2983),
.A2(n_2591),
.B1(n_2765),
.B2(n_2680),
.Y(n_3107)
);

NOR2x1_ASAP7_75t_SL g3108 ( 
.A(n_2816),
.B(n_2600),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2857),
.Y(n_3109)
);

OAI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_2983),
.A2(n_3021),
.B1(n_2970),
.B2(n_2842),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2954),
.B(n_2631),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_3000),
.A2(n_2783),
.B1(n_2680),
.B2(n_2765),
.Y(n_3112)
);

CKINVDCx5p33_ASAP7_75t_R g3113 ( 
.A(n_2842),
.Y(n_3113)
);

AOI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_2828),
.A2(n_2765),
.B1(n_2615),
.B2(n_2635),
.Y(n_3114)
);

AOI22xp33_ASAP7_75t_SL g3115 ( 
.A1(n_2955),
.A2(n_2600),
.B1(n_2604),
.B2(n_2711),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_SL g3116 ( 
.A1(n_2955),
.A2(n_2604),
.B1(n_2711),
.B2(n_2783),
.Y(n_3116)
);

AOI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_2997),
.A2(n_2783),
.B1(n_2683),
.B2(n_2641),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2975),
.B(n_2631),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_2909),
.B(n_2711),
.Y(n_3119)
);

NOR2x1_ASAP7_75t_SL g3120 ( 
.A(n_2816),
.B(n_2604),
.Y(n_3120)
);

AOI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_2997),
.A2(n_2641),
.B1(n_2665),
.B2(n_2631),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2888),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_2968),
.A2(n_2665),
.B1(n_2677),
.B2(n_2641),
.Y(n_3123)
);

INVx3_ASAP7_75t_L g3124 ( 
.A(n_2937),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2893),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_2866),
.A2(n_2665),
.B1(n_2677),
.B2(n_2641),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2911),
.Y(n_3127)
);

AND2x4_ASAP7_75t_L g3128 ( 
.A(n_2804),
.B(n_2788),
.Y(n_3128)
);

OAI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_2909),
.A2(n_2763),
.B1(n_2689),
.B2(n_2667),
.Y(n_3129)
);

INVx4_ASAP7_75t_L g3130 ( 
.A(n_2855),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2927),
.Y(n_3131)
);

OR2x2_ASAP7_75t_L g3132 ( 
.A(n_2877),
.B(n_2788),
.Y(n_3132)
);

OR2x2_ASAP7_75t_L g3133 ( 
.A(n_2839),
.B(n_2788),
.Y(n_3133)
);

INVx2_ASAP7_75t_SL g3134 ( 
.A(n_2823),
.Y(n_3134)
);

NAND2x1_ASAP7_75t_L g3135 ( 
.A(n_2831),
.B(n_2626),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2928),
.Y(n_3136)
);

OAI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2970),
.A2(n_2646),
.B1(n_2637),
.B2(n_2645),
.Y(n_3137)
);

OA21x2_ASAP7_75t_L g3138 ( 
.A1(n_3001),
.A2(n_2657),
.B(n_2644),
.Y(n_3138)
);

A2O1A1Ixp33_ASAP7_75t_L g3139 ( 
.A1(n_3022),
.A2(n_2614),
.B(n_2615),
.C(n_2613),
.Y(n_3139)
);

AOI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_2935),
.A2(n_2635),
.B1(n_2643),
.B2(n_2613),
.Y(n_3140)
);

OAI22xp33_ASAP7_75t_L g3141 ( 
.A1(n_2989),
.A2(n_2677),
.B1(n_2665),
.B2(n_2727),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_3013),
.A2(n_2677),
.B1(n_2643),
.B2(n_2657),
.Y(n_3142)
);

AOI22xp33_ASAP7_75t_L g3143 ( 
.A1(n_2921),
.A2(n_2644),
.B1(n_2727),
.B2(n_2563),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_3004),
.B(n_2538),
.Y(n_3144)
);

AND2x4_ASAP7_75t_L g3145 ( 
.A(n_2804),
.B(n_2538),
.Y(n_3145)
);

NOR2x1p5_ASAP7_75t_L g3146 ( 
.A(n_2850),
.B(n_2626),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2817),
.Y(n_3147)
);

AO21x2_ASAP7_75t_L g3148 ( 
.A1(n_2996),
.A2(n_2757),
.B(n_2750),
.Y(n_3148)
);

OAI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_3022),
.A2(n_3017),
.B1(n_2854),
.B2(n_2845),
.Y(n_3149)
);

AO21x2_ASAP7_75t_L g3150 ( 
.A1(n_2996),
.A2(n_2757),
.B(n_2750),
.Y(n_3150)
);

AOI22xp33_ASAP7_75t_L g3151 ( 
.A1(n_2967),
.A2(n_2727),
.B1(n_2565),
.B2(n_2570),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_2819),
.B(n_2563),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2956),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_2900),
.B(n_2565),
.Y(n_3154)
);

BUFx3_ASAP7_75t_L g3155 ( 
.A(n_2870),
.Y(n_3155)
);

INVx2_ASAP7_75t_SL g3156 ( 
.A(n_2876),
.Y(n_3156)
);

INVx3_ASAP7_75t_L g3157 ( 
.A(n_2937),
.Y(n_3157)
);

OAI21x1_ASAP7_75t_L g3158 ( 
.A1(n_2808),
.A2(n_2764),
.B(n_2645),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2810),
.B(n_2570),
.Y(n_3159)
);

INVx1_ASAP7_75t_SL g3160 ( 
.A(n_3017),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2941),
.A2(n_2727),
.B1(n_2571),
.B2(n_2652),
.Y(n_3161)
);

OAI21xp33_ASAP7_75t_SL g3162 ( 
.A1(n_2985),
.A2(n_2652),
.B(n_2637),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2830),
.Y(n_3163)
);

AOI21xp33_ASAP7_75t_L g3164 ( 
.A1(n_2859),
.A2(n_2571),
.B(n_2575),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2835),
.Y(n_3165)
);

NAND2xp33_ASAP7_75t_R g3166 ( 
.A(n_2977),
.B(n_73),
.Y(n_3166)
);

NAND4xp25_ASAP7_75t_L g3167 ( 
.A(n_2995),
.B(n_77),
.C(n_74),
.D(n_76),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2956),
.B(n_2575),
.Y(n_3168)
);

OAI222xp33_ASAP7_75t_L g3169 ( 
.A1(n_2972),
.A2(n_2919),
.B1(n_2913),
.B2(n_2929),
.C1(n_2854),
.C2(n_2831),
.Y(n_3169)
);

CKINVDCx6p67_ASAP7_75t_R g3170 ( 
.A(n_2940),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2844),
.Y(n_3171)
);

A2O1A1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_2902),
.A2(n_2750),
.B(n_2757),
.C(n_2575),
.Y(n_3172)
);

AND2x4_ASAP7_75t_L g3173 ( 
.A(n_2812),
.B(n_2575),
.Y(n_3173)
);

OA21x2_ASAP7_75t_L g3174 ( 
.A1(n_3001),
.A2(n_2878),
.B(n_2999),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_R g3175 ( 
.A(n_2977),
.B(n_2750),
.Y(n_3175)
);

OAI221xp5_ASAP7_75t_L g3176 ( 
.A1(n_2994),
.A2(n_2757),
.B1(n_80),
.B2(n_78),
.C(n_79),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2935),
.B(n_1021),
.Y(n_3177)
);

AO31x2_ASAP7_75t_L g3178 ( 
.A1(n_2914),
.A2(n_81),
.A3(n_78),
.B(n_80),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_2941),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_2812),
.B(n_2959),
.Y(n_3180)
);

AOI22xp33_ASAP7_75t_L g3181 ( 
.A1(n_2850),
.A2(n_85),
.B1(n_82),
.B2(n_84),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_2959),
.B(n_84),
.Y(n_3182)
);

OAI21x1_ASAP7_75t_L g3183 ( 
.A1(n_2805),
.A2(n_491),
.B(n_490),
.Y(n_3183)
);

OAI22xp5_ASAP7_75t_L g3184 ( 
.A1(n_2841),
.A2(n_2833),
.B1(n_2988),
.B2(n_2890),
.Y(n_3184)
);

AOI22xp33_ASAP7_75t_L g3185 ( 
.A1(n_2905),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_3185)
);

CKINVDCx11_ASAP7_75t_R g3186 ( 
.A(n_2870),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2969),
.B(n_87),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2969),
.Y(n_3188)
);

AOI22xp33_ASAP7_75t_L g3189 ( 
.A1(n_2987),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2971),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2914),
.A2(n_2853),
.B(n_2841),
.Y(n_3191)
);

INVx6_ASAP7_75t_L g3192 ( 
.A(n_3003),
.Y(n_3192)
);

CKINVDCx11_ASAP7_75t_R g3193 ( 
.A(n_2829),
.Y(n_3193)
);

AOI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_2853),
.A2(n_1296),
.B(n_1266),
.Y(n_3194)
);

NAND2xp33_ASAP7_75t_SL g3195 ( 
.A(n_2889),
.B(n_90),
.Y(n_3195)
);

HB1xp67_ASAP7_75t_L g3196 ( 
.A(n_2961),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_2998),
.B(n_92),
.Y(n_3197)
);

INVx3_ASAP7_75t_L g3198 ( 
.A(n_3002),
.Y(n_3198)
);

AOI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_2859),
.A2(n_1021),
.B1(n_1045),
.B2(n_1032),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2971),
.Y(n_3200)
);

CKINVDCx6p67_ASAP7_75t_R g3201 ( 
.A(n_3003),
.Y(n_3201)
);

A2O1A1Ixp33_ASAP7_75t_L g3202 ( 
.A1(n_2951),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_3202)
);

OAI21x1_ASAP7_75t_L g3203 ( 
.A1(n_2847),
.A2(n_494),
.B(n_492),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3015),
.B(n_94),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3018),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_SL g3206 ( 
.A(n_2894),
.B(n_1021),
.Y(n_3206)
);

AO22x1_ASAP7_75t_L g3207 ( 
.A1(n_2973),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2998),
.B(n_95),
.Y(n_3208)
);

OAI21x1_ASAP7_75t_L g3209 ( 
.A1(n_2824),
.A2(n_498),
.B(n_496),
.Y(n_3209)
);

AND2x4_ASAP7_75t_L g3210 ( 
.A(n_3002),
.B(n_97),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2946),
.B(n_99),
.Y(n_3211)
);

INVx6_ASAP7_75t_L g3212 ( 
.A(n_2851),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3023),
.B(n_2809),
.Y(n_3213)
);

BUFx2_ASAP7_75t_L g3214 ( 
.A(n_2851),
.Y(n_3214)
);

INVx4_ASAP7_75t_L g3215 ( 
.A(n_2865),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2865),
.Y(n_3216)
);

CKINVDCx20_ASAP7_75t_R g3217 ( 
.A(n_2899),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2961),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_L g3219 ( 
.A(n_3026),
.Y(n_3219)
);

OA21x2_ASAP7_75t_L g3220 ( 
.A1(n_3218),
.A2(n_2848),
.B(n_2896),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3026),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3045),
.B(n_2818),
.Y(n_3222)
);

BUFx2_ASAP7_75t_L g3223 ( 
.A(n_3162),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3057),
.Y(n_3224)
);

INVx3_ASAP7_75t_L g3225 ( 
.A(n_3180),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3057),
.Y(n_3226)
);

BUFx2_ASAP7_75t_SL g3227 ( 
.A(n_3130),
.Y(n_3227)
);

BUFx2_ASAP7_75t_L g3228 ( 
.A(n_3138),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3196),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_3196),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3058),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_3138),
.Y(n_3232)
);

OAI21x1_ASAP7_75t_L g3233 ( 
.A1(n_3191),
.A2(n_3194),
.B(n_3135),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3058),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3062),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_3031),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3034),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3043),
.Y(n_3238)
);

OAI21x1_ASAP7_75t_SL g3239 ( 
.A1(n_3108),
.A2(n_2991),
.B(n_2944),
.Y(n_3239)
);

HB1xp67_ASAP7_75t_L g3240 ( 
.A(n_3062),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3050),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3079),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3188),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_3038),
.Y(n_3244)
);

HB1xp67_ASAP7_75t_L g3245 ( 
.A(n_3133),
.Y(n_3245)
);

AND2x4_ASAP7_75t_L g3246 ( 
.A(n_3128),
.B(n_2831),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_3042),
.Y(n_3247)
);

HB1xp67_ASAP7_75t_L g3248 ( 
.A(n_3054),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3200),
.Y(n_3249)
);

OA21x2_ASAP7_75t_L g3250 ( 
.A1(n_3191),
.A2(n_2897),
.B(n_2871),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3051),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3053),
.Y(n_3252)
);

OA21x2_ASAP7_75t_L g3253 ( 
.A1(n_3194),
.A2(n_2864),
.B(n_2884),
.Y(n_3253)
);

AO31x2_ASAP7_75t_L g3254 ( 
.A1(n_3120),
.A2(n_2945),
.A3(n_2833),
.B(n_2981),
.Y(n_3254)
);

AND2x4_ASAP7_75t_SL g3255 ( 
.A(n_3077),
.B(n_2865),
.Y(n_3255)
);

BUFx2_ASAP7_75t_L g3256 ( 
.A(n_3148),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3074),
.Y(n_3257)
);

AO21x2_ASAP7_75t_L g3258 ( 
.A1(n_3027),
.A2(n_3150),
.B(n_3148),
.Y(n_3258)
);

AO21x2_ASAP7_75t_L g3259 ( 
.A1(n_3027),
.A2(n_2863),
.B(n_2906),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3075),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_3180),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3213),
.B(n_2858),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3080),
.Y(n_3263)
);

OAI21x1_ASAP7_75t_L g3264 ( 
.A1(n_3158),
.A2(n_2807),
.B(n_2881),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_3102),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3103),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3090),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3094),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3106),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_3212),
.Y(n_3270)
);

HB1xp67_ASAP7_75t_L g3271 ( 
.A(n_3132),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3101),
.Y(n_3272)
);

INVxp33_ASAP7_75t_L g3273 ( 
.A(n_3095),
.Y(n_3273)
);

OAI21x1_ASAP7_75t_L g3274 ( 
.A1(n_3174),
.A2(n_2807),
.B(n_2881),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_3036),
.B(n_2827),
.Y(n_3275)
);

BUFx4f_ASAP7_75t_SL g3276 ( 
.A(n_3217),
.Y(n_3276)
);

AO31x2_ASAP7_75t_L g3277 ( 
.A1(n_3184),
.A2(n_2856),
.A3(n_2930),
.B(n_3005),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_3109),
.Y(n_3278)
);

INVx2_ASAP7_75t_SL g3279 ( 
.A(n_3212),
.Y(n_3279)
);

OR2x2_ASAP7_75t_L g3280 ( 
.A(n_3033),
.B(n_2814),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_3153),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3122),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3125),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_SL g3284 ( 
.A1(n_3172),
.A2(n_2944),
.B(n_3010),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3190),
.Y(n_3285)
);

OAI21x1_ASAP7_75t_L g3286 ( 
.A1(n_3174),
.A2(n_2881),
.B(n_2861),
.Y(n_3286)
);

AND2x4_ASAP7_75t_L g3287 ( 
.A(n_3128),
.B(n_2858),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3127),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3131),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3136),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_3048),
.B(n_2827),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3147),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3163),
.Y(n_3293)
);

BUFx2_ASAP7_75t_L g3294 ( 
.A(n_3150),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3104),
.B(n_3030),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_3165),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_3152),
.B(n_2827),
.Y(n_3297)
);

BUFx3_ASAP7_75t_L g3298 ( 
.A(n_3170),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3171),
.Y(n_3299)
);

AOI22xp33_ASAP7_75t_L g3300 ( 
.A1(n_3066),
.A2(n_2837),
.B1(n_2858),
.B2(n_2904),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_3205),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3033),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_3029),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3029),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3070),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3033),
.Y(n_3306)
);

BUFx3_ASAP7_75t_L g3307 ( 
.A(n_3186),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_3063),
.B(n_2894),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3033),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_3168),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3071),
.B(n_2939),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3071),
.B(n_2939),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3104),
.B(n_2858),
.Y(n_3313)
);

HB1xp67_ASAP7_75t_L g3314 ( 
.A(n_3111),
.Y(n_3314)
);

HB1xp67_ASAP7_75t_L g3315 ( 
.A(n_3118),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3105),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3083),
.Y(n_3317)
);

OAI21x1_ASAP7_75t_L g3318 ( 
.A1(n_3078),
.A2(n_2961),
.B(n_2860),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3214),
.Y(n_3319)
);

AO21x1_ASAP7_75t_SL g3320 ( 
.A1(n_3073),
.A2(n_3005),
.B(n_2960),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3198),
.Y(n_3321)
);

BUFx3_ASAP7_75t_L g3322 ( 
.A(n_3192),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3198),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3084),
.B(n_2821),
.Y(n_3324)
);

BUFx2_ASAP7_75t_R g3325 ( 
.A(n_3098),
.Y(n_3325)
);

INVx3_ASAP7_75t_L g3326 ( 
.A(n_3173),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3084),
.Y(n_3327)
);

NAND2xp33_ASAP7_75t_R g3328 ( 
.A(n_3175),
.B(n_3010),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3124),
.Y(n_3329)
);

HB1xp67_ASAP7_75t_L g3330 ( 
.A(n_3099),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_3124),
.B(n_2821),
.Y(n_3331)
);

OR2x2_ASAP7_75t_L g3332 ( 
.A(n_3041),
.B(n_3157),
.Y(n_3332)
);

OR2x6_ASAP7_75t_L g3333 ( 
.A(n_3037),
.B(n_2936),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3157),
.Y(n_3334)
);

INVx4_ASAP7_75t_L g3335 ( 
.A(n_3130),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3216),
.Y(n_3336)
);

INVx4_ASAP7_75t_L g3337 ( 
.A(n_3192),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3037),
.B(n_2826),
.Y(n_3338)
);

OA21x2_ASAP7_75t_L g3339 ( 
.A1(n_3161),
.A2(n_2891),
.B(n_2852),
.Y(n_3339)
);

HB1xp67_ASAP7_75t_L g3340 ( 
.A(n_3059),
.Y(n_3340)
);

HB1xp67_ASAP7_75t_L g3341 ( 
.A(n_3082),
.Y(n_3341)
);

OAI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_3086),
.A2(n_2994),
.B(n_3019),
.Y(n_3342)
);

INVx3_ASAP7_75t_L g3343 ( 
.A(n_3173),
.Y(n_3343)
);

HB1xp67_ASAP7_75t_L g3344 ( 
.A(n_3144),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3216),
.Y(n_3345)
);

HB1xp67_ASAP7_75t_L g3346 ( 
.A(n_3145),
.Y(n_3346)
);

BUFx6f_ASAP7_75t_L g3347 ( 
.A(n_3076),
.Y(n_3347)
);

HB1xp67_ASAP7_75t_L g3348 ( 
.A(n_3145),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3187),
.Y(n_3349)
);

AOI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_3091),
.A2(n_2858),
.B1(n_2826),
.B2(n_3016),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3076),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3164),
.B(n_2814),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3076),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3178),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3178),
.Y(n_3355)
);

OR2x2_ASAP7_75t_L g3356 ( 
.A(n_3088),
.B(n_2814),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3178),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3178),
.Y(n_3358)
);

OAI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3086),
.A2(n_3010),
.B(n_2925),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3076),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3032),
.B(n_2803),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3088),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3097),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3097),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3088),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3088),
.Y(n_3366)
);

INVx3_ASAP7_75t_L g3367 ( 
.A(n_3044),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3044),
.B(n_2803),
.Y(n_3368)
);

INVx3_ASAP7_75t_L g3369 ( 
.A(n_3097),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3097),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3116),
.Y(n_3371)
);

HB1xp67_ASAP7_75t_L g3372 ( 
.A(n_3134),
.Y(n_3372)
);

OR2x2_ASAP7_75t_L g3373 ( 
.A(n_3156),
.B(n_2815),
.Y(n_3373)
);

NOR2x1_ASAP7_75t_SL g3374 ( 
.A(n_3096),
.B(n_2906),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3182),
.Y(n_3375)
);

INVx3_ASAP7_75t_L g3376 ( 
.A(n_3215),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3116),
.Y(n_3377)
);

AOI222xp33_ASAP7_75t_L g3378 ( 
.A1(n_3342),
.A2(n_3091),
.B1(n_3181),
.B2(n_3110),
.C1(n_3189),
.C2(n_3176),
.Y(n_3378)
);

BUFx12f_ASAP7_75t_L g3379 ( 
.A(n_3307),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3369),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3292),
.Y(n_3381)
);

OAI22xp5_ASAP7_75t_L g3382 ( 
.A1(n_3300),
.A2(n_3055),
.B1(n_3112),
.B2(n_3179),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3320),
.A2(n_3185),
.B1(n_3167),
.B2(n_3181),
.Y(n_3383)
);

AOI21xp33_ASAP7_75t_L g3384 ( 
.A1(n_3340),
.A2(n_3149),
.B(n_3166),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_L g3385 ( 
.A(n_3273),
.B(n_3063),
.Y(n_3385)
);

OAI21xp33_ASAP7_75t_SL g3386 ( 
.A1(n_3377),
.A2(n_3179),
.B(n_3032),
.Y(n_3386)
);

OR2x2_ASAP7_75t_L g3387 ( 
.A(n_3330),
.B(n_3087),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3367),
.B(n_3089),
.Y(n_3388)
);

HB1xp67_ASAP7_75t_L g3389 ( 
.A(n_3219),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3317),
.B(n_3093),
.Y(n_3390)
);

OAI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3350),
.A2(n_3055),
.B1(n_3112),
.B2(n_3060),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3292),
.Y(n_3392)
);

AOI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_3359),
.A2(n_3046),
.B(n_3073),
.Y(n_3393)
);

OAI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3371),
.A2(n_3067),
.B1(n_3052),
.B2(n_3107),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3369),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_L g3396 ( 
.A1(n_3320),
.A2(n_3185),
.B1(n_3047),
.B2(n_3060),
.Y(n_3396)
);

HB1xp67_ASAP7_75t_L g3397 ( 
.A(n_3240),
.Y(n_3397)
);

INVxp67_ASAP7_75t_L g3398 ( 
.A(n_3248),
.Y(n_3398)
);

BUFx2_ASAP7_75t_SL g3399 ( 
.A(n_3307),
.Y(n_3399)
);

OAI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3325),
.A2(n_3028),
.B1(n_3143),
.B2(n_3065),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3317),
.B(n_3100),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3367),
.B(n_3154),
.Y(n_3402)
);

AOI221xp5_ASAP7_75t_L g3403 ( 
.A1(n_3377),
.A2(n_3211),
.B1(n_3207),
.B2(n_3189),
.C(n_3169),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_3367),
.B(n_3061),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3367),
.B(n_3068),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3293),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3349),
.B(n_3115),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3346),
.B(n_3068),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_L g3409 ( 
.A1(n_3371),
.A2(n_3065),
.B1(n_3211),
.B2(n_3028),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3293),
.Y(n_3410)
);

AOI211xp5_ASAP7_75t_L g3411 ( 
.A1(n_3284),
.A2(n_3169),
.B(n_3141),
.C(n_3049),
.Y(n_3411)
);

BUFx3_ASAP7_75t_L g3412 ( 
.A(n_3307),
.Y(n_3412)
);

INVx3_ASAP7_75t_L g3413 ( 
.A(n_3335),
.Y(n_3413)
);

OAI211xp5_ASAP7_75t_L g3414 ( 
.A1(n_3284),
.A2(n_3115),
.B(n_3081),
.C(n_3143),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3349),
.B(n_3081),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3316),
.B(n_3039),
.Y(n_3416)
);

AO221x1_ASAP7_75t_L g3417 ( 
.A1(n_3223),
.A2(n_3141),
.B1(n_3129),
.B2(n_3137),
.C(n_3035),
.Y(n_3417)
);

AOI22xp33_ASAP7_75t_L g3418 ( 
.A1(n_3259),
.A2(n_3025),
.B1(n_3195),
.B2(n_3040),
.Y(n_3418)
);

OAI22xp33_ASAP7_75t_L g3419 ( 
.A1(n_3328),
.A2(n_3064),
.B1(n_3072),
.B2(n_3114),
.Y(n_3419)
);

AOI21x1_ASAP7_75t_L g3420 ( 
.A1(n_3256),
.A2(n_3204),
.B(n_3119),
.Y(n_3420)
);

OR2x2_ASAP7_75t_L g3421 ( 
.A(n_3245),
.B(n_3039),
.Y(n_3421)
);

NAND3xp33_ASAP7_75t_L g3422 ( 
.A(n_3352),
.B(n_3123),
.C(n_3202),
.Y(n_3422)
);

AOI22xp33_ASAP7_75t_L g3423 ( 
.A1(n_3259),
.A2(n_3025),
.B1(n_3092),
.B2(n_3123),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3348),
.B(n_3159),
.Y(n_3424)
);

OR2x2_ASAP7_75t_L g3425 ( 
.A(n_3271),
.B(n_3332),
.Y(n_3425)
);

AOI22xp5_ASAP7_75t_L g3426 ( 
.A1(n_3313),
.A2(n_3085),
.B1(n_3092),
.B2(n_3177),
.Y(n_3426)
);

OAI211xp5_ASAP7_75t_L g3427 ( 
.A1(n_3361),
.A2(n_3161),
.B(n_3121),
.C(n_3046),
.Y(n_3427)
);

INVx2_ASAP7_75t_SL g3428 ( 
.A(n_3298),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3259),
.A2(n_3151),
.B1(n_3117),
.B2(n_3142),
.Y(n_3429)
);

CKINVDCx20_ASAP7_75t_R g3430 ( 
.A(n_3276),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3299),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3262),
.A2(n_3151),
.B1(n_3117),
.B2(n_3142),
.Y(n_3432)
);

OAI22xp33_ASAP7_75t_SL g3433 ( 
.A1(n_3223),
.A2(n_3337),
.B1(n_3335),
.B2(n_3228),
.Y(n_3433)
);

OR2x2_ASAP7_75t_L g3434 ( 
.A(n_3332),
.B(n_3121),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3299),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3369),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_3295),
.A2(n_3375),
.B1(n_3298),
.B2(n_3258),
.Y(n_3437)
);

OAI221xp5_ASAP7_75t_L g3438 ( 
.A1(n_3227),
.A2(n_3056),
.B1(n_3140),
.B2(n_3160),
.C(n_3139),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3267),
.Y(n_3439)
);

OAI22xp5_ASAP7_75t_SL g3440 ( 
.A1(n_3298),
.A2(n_3192),
.B1(n_3113),
.B2(n_3155),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3344),
.B(n_3146),
.Y(n_3441)
);

OR2x2_ASAP7_75t_L g3442 ( 
.A(n_3341),
.B(n_2803),
.Y(n_3442)
);

OAI211xp5_ASAP7_75t_SL g3443 ( 
.A1(n_3375),
.A2(n_3193),
.B(n_3199),
.C(n_3126),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3267),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3268),
.Y(n_3445)
);

AOI22xp33_ASAP7_75t_L g3446 ( 
.A1(n_3375),
.A2(n_3258),
.B1(n_3355),
.B2(n_3354),
.Y(n_3446)
);

AO31x2_ASAP7_75t_L g3447 ( 
.A1(n_3354),
.A2(n_3215),
.A3(n_2856),
.B(n_3005),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3258),
.A2(n_3182),
.B1(n_3210),
.B2(n_2944),
.Y(n_3448)
);

AOI222xp33_ASAP7_75t_L g3449 ( 
.A1(n_3355),
.A2(n_2882),
.B1(n_3208),
.B2(n_3197),
.C1(n_3210),
.C2(n_2925),
.Y(n_3449)
);

OAI21x1_ASAP7_75t_L g3450 ( 
.A1(n_3233),
.A2(n_3183),
.B(n_3209),
.Y(n_3450)
);

OAI221xp5_ASAP7_75t_L g3451 ( 
.A1(n_3227),
.A2(n_3126),
.B1(n_3069),
.B2(n_3206),
.C(n_3212),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3357),
.A2(n_2815),
.B1(n_3201),
.B2(n_2889),
.Y(n_3452)
);

OAI21x1_ASAP7_75t_L g3453 ( 
.A1(n_3233),
.A2(n_3203),
.B(n_2815),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3357),
.A2(n_3016),
.B1(n_3014),
.B2(n_2874),
.Y(n_3454)
);

CKINVDCx20_ASAP7_75t_R g3455 ( 
.A(n_3255),
.Y(n_3455)
);

AOI22xp33_ASAP7_75t_L g3456 ( 
.A1(n_3287),
.A2(n_3129),
.B1(n_3014),
.B2(n_2885),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_SL g3457 ( 
.A1(n_3374),
.A2(n_3005),
.B1(n_2960),
.B2(n_2965),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3335),
.B(n_2865),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3369),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3268),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3272),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_3337),
.B(n_3335),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3272),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3282),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_SL g3465 ( 
.A1(n_3374),
.A2(n_2960),
.B1(n_2993),
.B2(n_2965),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3347),
.Y(n_3466)
);

AOI221xp5_ASAP7_75t_L g3467 ( 
.A1(n_3358),
.A2(n_3228),
.B1(n_3316),
.B2(n_3222),
.C(n_3239),
.Y(n_3467)
);

INVx11_ASAP7_75t_L g3468 ( 
.A(n_3308),
.Y(n_3468)
);

AOI21xp33_ASAP7_75t_L g3469 ( 
.A1(n_3239),
.A2(n_2993),
.B(n_2965),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3347),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_SL g3471 ( 
.A1(n_3322),
.A2(n_3337),
.B1(n_3287),
.B2(n_3255),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3282),
.Y(n_3472)
);

BUFx6f_ASAP7_75t_L g3473 ( 
.A(n_3347),
.Y(n_3473)
);

OAI22xp33_ASAP7_75t_L g3474 ( 
.A1(n_3322),
.A2(n_2960),
.B1(n_2993),
.B2(n_2965),
.Y(n_3474)
);

NAND3xp33_ASAP7_75t_L g3475 ( 
.A(n_3358),
.B(n_2892),
.C(n_2885),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3314),
.B(n_2803),
.Y(n_3476)
);

NOR2xp67_ASAP7_75t_L g3477 ( 
.A(n_3337),
.B(n_2993),
.Y(n_3477)
);

AOI22xp33_ASAP7_75t_L g3478 ( 
.A1(n_3322),
.A2(n_2874),
.B1(n_2979),
.B2(n_2966),
.Y(n_3478)
);

OAI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3333),
.A2(n_2982),
.B1(n_3009),
.B2(n_2936),
.Y(n_3479)
);

AOI22xp33_ASAP7_75t_L g3480 ( 
.A1(n_3287),
.A2(n_3020),
.B1(n_2984),
.B2(n_2980),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3315),
.B(n_2912),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_L g3482 ( 
.A1(n_3287),
.A2(n_2901),
.B1(n_3012),
.B2(n_3011),
.Y(n_3482)
);

HB1xp67_ASAP7_75t_L g3483 ( 
.A(n_3229),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3310),
.B(n_2912),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3305),
.A2(n_2907),
.B1(n_2957),
.B2(n_2934),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3347),
.Y(n_3486)
);

AO21x2_ASAP7_75t_L g3487 ( 
.A1(n_3303),
.A2(n_2943),
.B(n_2933),
.Y(n_3487)
);

HB1xp67_ASAP7_75t_L g3488 ( 
.A(n_3229),
.Y(n_3488)
);

BUFx4f_ASAP7_75t_SL g3489 ( 
.A(n_3347),
.Y(n_3489)
);

AOI22xp33_ASAP7_75t_SL g3490 ( 
.A1(n_3255),
.A2(n_2947),
.B1(n_2964),
.B2(n_2958),
.Y(n_3490)
);

AOI22xp33_ASAP7_75t_SL g3491 ( 
.A1(n_3246),
.A2(n_3009),
.B1(n_2982),
.B2(n_2923),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3283),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3283),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_SL g3494 ( 
.A1(n_3246),
.A2(n_3338),
.B1(n_3368),
.B2(n_3291),
.Y(n_3494)
);

AOI22xp33_ASAP7_75t_L g3495 ( 
.A1(n_3305),
.A2(n_2910),
.B1(n_3008),
.B2(n_2986),
.Y(n_3495)
);

NOR2x1_ASAP7_75t_L g3496 ( 
.A(n_3376),
.B(n_2869),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3301),
.Y(n_3497)
);

OAI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_3333),
.A2(n_2836),
.B1(n_2915),
.B2(n_2912),
.Y(n_3498)
);

AOI221xp5_ASAP7_75t_L g3499 ( 
.A1(n_3275),
.A2(n_2868),
.B1(n_102),
.B2(n_100),
.C(n_101),
.Y(n_3499)
);

AOI211xp5_ASAP7_75t_L g3500 ( 
.A1(n_3356),
.A2(n_3338),
.B(n_3280),
.C(n_3373),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3327),
.Y(n_3501)
);

OAI211xp5_ASAP7_75t_SL g3502 ( 
.A1(n_3373),
.A2(n_3232),
.B(n_3304),
.C(n_3303),
.Y(n_3502)
);

AOI22xp33_ASAP7_75t_L g3503 ( 
.A1(n_3372),
.A2(n_2836),
.B1(n_2869),
.B2(n_2868),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3310),
.B(n_2912),
.Y(n_3504)
);

HB1xp67_ASAP7_75t_L g3505 ( 
.A(n_3230),
.Y(n_3505)
);

OAI21xp5_ASAP7_75t_SL g3506 ( 
.A1(n_3246),
.A2(n_2915),
.B(n_101),
.Y(n_3506)
);

AOI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_3246),
.A2(n_2836),
.B1(n_2915),
.B2(n_105),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_L g3508 ( 
.A1(n_3319),
.A2(n_3291),
.B1(n_3275),
.B2(n_3224),
.Y(n_3508)
);

OAI21x1_ASAP7_75t_L g3509 ( 
.A1(n_3318),
.A2(n_2880),
.B(n_2915),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3501),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3381),
.Y(n_3511)
);

HB1xp67_ASAP7_75t_L g3512 ( 
.A(n_3389),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3392),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3406),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3422),
.B(n_3297),
.Y(n_3515)
);

INVx1_ASAP7_75t_SL g3516 ( 
.A(n_3399),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3380),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3410),
.Y(n_3518)
);

NOR2x1_ASAP7_75t_SL g3519 ( 
.A(n_3414),
.B(n_3333),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3494),
.B(n_3326),
.Y(n_3520)
);

AND2x4_ASAP7_75t_L g3521 ( 
.A(n_3413),
.B(n_3232),
.Y(n_3521)
);

BUFx2_ASAP7_75t_L g3522 ( 
.A(n_3379),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3395),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3405),
.B(n_3326),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3398),
.B(n_3297),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3471),
.B(n_3326),
.Y(n_3526)
);

NOR2x1_ASAP7_75t_L g3527 ( 
.A(n_3412),
.B(n_3413),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3436),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3431),
.Y(n_3529)
);

INVx3_ASAP7_75t_L g3530 ( 
.A(n_3473),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3383),
.A2(n_3333),
.B1(n_3343),
.B2(n_3326),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3435),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3459),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3473),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3439),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3444),
.Y(n_3536)
);

INVx3_ASAP7_75t_L g3537 ( 
.A(n_3473),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3445),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3416),
.B(n_3301),
.Y(n_3539)
);

AND2x4_ASAP7_75t_L g3540 ( 
.A(n_3462),
.B(n_3362),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_3473),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3388),
.B(n_3343),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3483),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3402),
.B(n_3343),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3508),
.B(n_3343),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3460),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3508),
.B(n_3225),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3466),
.B(n_3225),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3461),
.Y(n_3549)
);

OR2x2_ASAP7_75t_L g3550 ( 
.A(n_3476),
.B(n_3221),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3463),
.Y(n_3551)
);

INVx2_ASAP7_75t_SL g3552 ( 
.A(n_3489),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3407),
.B(n_3319),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_SL g3554 ( 
.A1(n_3417),
.A2(n_3368),
.B1(n_3261),
.B2(n_3225),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3464),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3470),
.B(n_3225),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_3486),
.B(n_3261),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3404),
.B(n_3261),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3472),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3492),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3483),
.Y(n_3561)
);

HB1xp67_ASAP7_75t_L g3562 ( 
.A(n_3389),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3493),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_3440),
.B(n_3270),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3441),
.B(n_3261),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3488),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3408),
.B(n_3270),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3437),
.B(n_3279),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3497),
.Y(n_3569)
);

OR2x2_ASAP7_75t_L g3570 ( 
.A(n_3481),
.B(n_3221),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3437),
.B(n_3279),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3397),
.Y(n_3572)
);

AND2x2_ASAP7_75t_L g3573 ( 
.A(n_3397),
.B(n_3428),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3425),
.B(n_3351),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3415),
.B(n_3296),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3409),
.B(n_3296),
.Y(n_3576)
);

AND2x4_ASAP7_75t_L g3577 ( 
.A(n_3477),
.B(n_3362),
.Y(n_3577)
);

OR2x2_ASAP7_75t_L g3578 ( 
.A(n_3442),
.B(n_3224),
.Y(n_3578)
);

AND2x4_ASAP7_75t_L g3579 ( 
.A(n_3455),
.B(n_3496),
.Y(n_3579)
);

HB1xp67_ASAP7_75t_L g3580 ( 
.A(n_3434),
.Y(n_3580)
);

OR2x2_ASAP7_75t_L g3581 ( 
.A(n_3484),
.B(n_3226),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3488),
.Y(n_3582)
);

AND2x4_ASAP7_75t_L g3583 ( 
.A(n_3393),
.B(n_3365),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3424),
.B(n_3351),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3500),
.B(n_3353),
.Y(n_3585)
);

BUFx3_ASAP7_75t_L g3586 ( 
.A(n_3430),
.Y(n_3586)
);

INVx2_ASAP7_75t_L g3587 ( 
.A(n_3505),
.Y(n_3587)
);

HB1xp67_ASAP7_75t_L g3588 ( 
.A(n_3421),
.Y(n_3588)
);

BUFx6f_ASAP7_75t_L g3589 ( 
.A(n_3450),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3505),
.Y(n_3590)
);

AOI22xp33_ASAP7_75t_L g3591 ( 
.A1(n_3378),
.A2(n_3333),
.B1(n_3339),
.B2(n_3376),
.Y(n_3591)
);

NAND2x1p5_ASAP7_75t_L g3592 ( 
.A(n_3420),
.B(n_3274),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3409),
.B(n_3288),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3403),
.B(n_3288),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3504),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3447),
.Y(n_3596)
);

OR2x2_ASAP7_75t_L g3597 ( 
.A(n_3446),
.B(n_3226),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_3411),
.B(n_3467),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3427),
.B(n_3289),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3446),
.B(n_3353),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3465),
.B(n_3360),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3387),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3447),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3458),
.B(n_3360),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3509),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3429),
.B(n_3363),
.Y(n_3606)
);

NOR2x1_ASAP7_75t_L g3607 ( 
.A(n_3385),
.B(n_3376),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3489),
.Y(n_3608)
);

BUFx2_ASAP7_75t_L g3609 ( 
.A(n_3447),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3487),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3448),
.B(n_3363),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3390),
.Y(n_3612)
);

NOR2x1p5_ASAP7_75t_L g3613 ( 
.A(n_3401),
.B(n_3376),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3386),
.B(n_3289),
.Y(n_3614)
);

OR2x2_ASAP7_75t_L g3615 ( 
.A(n_3447),
.B(n_3231),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_3448),
.B(n_3364),
.Y(n_3616)
);

AOI22xp33_ASAP7_75t_SL g3617 ( 
.A1(n_3382),
.A2(n_3256),
.B1(n_3294),
.B2(n_3356),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3433),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3506),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3475),
.Y(n_3620)
);

AOI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3396),
.A2(n_3339),
.B1(n_3331),
.B2(n_3324),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3457),
.Y(n_3622)
);

OR2x2_ASAP7_75t_L g3623 ( 
.A(n_3474),
.B(n_3231),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3419),
.B(n_3290),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3474),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3423),
.B(n_3364),
.Y(n_3626)
);

AOI22xp33_ASAP7_75t_L g3627 ( 
.A1(n_3396),
.A2(n_3339),
.B1(n_3331),
.B2(n_3324),
.Y(n_3627)
);

HB1xp67_ASAP7_75t_L g3628 ( 
.A(n_3487),
.Y(n_3628)
);

HB1xp67_ASAP7_75t_L g3629 ( 
.A(n_3498),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_3419),
.B(n_3311),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3453),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3384),
.B(n_3290),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3426),
.B(n_3234),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3432),
.B(n_3234),
.Y(n_3634)
);

BUFx2_ASAP7_75t_L g3635 ( 
.A(n_3394),
.Y(n_3635)
);

NOR2xp67_ASAP7_75t_L g3636 ( 
.A(n_3579),
.B(n_3451),
.Y(n_3636)
);

OAI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3622),
.A2(n_3391),
.B1(n_3394),
.B2(n_3400),
.Y(n_3637)
);

BUFx6f_ASAP7_75t_L g3638 ( 
.A(n_3522),
.Y(n_3638)
);

AOI22xp33_ASAP7_75t_SL g3639 ( 
.A1(n_3635),
.A2(n_3438),
.B1(n_3383),
.B2(n_3418),
.Y(n_3639)
);

INVx3_ASAP7_75t_L g3640 ( 
.A(n_3521),
.Y(n_3640)
);

AOI22xp33_ASAP7_75t_SL g3641 ( 
.A1(n_3635),
.A2(n_3418),
.B1(n_3294),
.B2(n_3479),
.Y(n_3641)
);

OR2x6_ASAP7_75t_L g3642 ( 
.A(n_3527),
.B(n_3264),
.Y(n_3642)
);

HB1xp67_ASAP7_75t_L g3643 ( 
.A(n_3512),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3522),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3511),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3530),
.Y(n_3646)
);

AOI22xp33_ASAP7_75t_L g3647 ( 
.A1(n_3598),
.A2(n_3499),
.B1(n_3423),
.B2(n_3443),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3530),
.Y(n_3648)
);

OAI31xp33_ASAP7_75t_SL g3649 ( 
.A1(n_3598),
.A2(n_3502),
.A3(n_3491),
.B(n_3490),
.Y(n_3649)
);

HB1xp67_ASAP7_75t_L g3650 ( 
.A(n_3562),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3530),
.Y(n_3651)
);

OAI221xp5_ASAP7_75t_L g3652 ( 
.A1(n_3619),
.A2(n_3456),
.B1(n_3507),
.B2(n_3452),
.C(n_3454),
.Y(n_3652)
);

OAI21x1_ASAP7_75t_L g3653 ( 
.A1(n_3592),
.A2(n_3230),
.B(n_3304),
.Y(n_3653)
);

OAI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_3554),
.A2(n_3507),
.B(n_3449),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3537),
.Y(n_3655)
);

AOI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_3622),
.A2(n_3454),
.B1(n_3452),
.B2(n_3503),
.Y(n_3656)
);

INVx1_ASAP7_75t_SL g3657 ( 
.A(n_3516),
.Y(n_3657)
);

INVx3_ASAP7_75t_L g3658 ( 
.A(n_3521),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3511),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_SL g3660 ( 
.A1(n_3617),
.A2(n_3503),
.B(n_3478),
.Y(n_3660)
);

INVx2_ASAP7_75t_SL g3661 ( 
.A(n_3586),
.Y(n_3661)
);

AND2x2_ASAP7_75t_L g3662 ( 
.A(n_3567),
.B(n_3370),
.Y(n_3662)
);

OAI211xp5_ASAP7_75t_L g3663 ( 
.A1(n_3621),
.A2(n_3469),
.B(n_3478),
.C(n_3482),
.Y(n_3663)
);

OAI31xp33_ASAP7_75t_L g3664 ( 
.A1(n_3531),
.A2(n_3630),
.A3(n_3618),
.B(n_3591),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3513),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3513),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3567),
.B(n_3370),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3537),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3604),
.B(n_3327),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3588),
.B(n_3277),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3580),
.B(n_3277),
.Y(n_3671)
);

OAI211xp5_ASAP7_75t_L g3672 ( 
.A1(n_3627),
.A2(n_3485),
.B(n_3495),
.C(n_3480),
.Y(n_3672)
);

INVx1_ASAP7_75t_SL g3673 ( 
.A(n_3573),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3537),
.Y(n_3674)
);

AOI221xp5_ASAP7_75t_L g3675 ( 
.A1(n_3620),
.A2(n_3302),
.B1(n_3306),
.B2(n_3280),
.C(n_3309),
.Y(n_3675)
);

OAI21x1_ASAP7_75t_L g3676 ( 
.A1(n_3592),
.A2(n_3607),
.B(n_3623),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3521),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3565),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3565),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3577),
.Y(n_3680)
);

AND2x4_ASAP7_75t_L g3681 ( 
.A(n_3552),
.B(n_3311),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3576),
.B(n_3235),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3518),
.Y(n_3683)
);

OAI221xp5_ASAP7_75t_L g3684 ( 
.A1(n_3594),
.A2(n_3485),
.B1(n_3495),
.B2(n_3366),
.C(n_3365),
.Y(n_3684)
);

AOI221xp5_ASAP7_75t_L g3685 ( 
.A1(n_3625),
.A2(n_3306),
.B1(n_3302),
.B2(n_3309),
.C(n_3235),
.Y(n_3685)
);

NOR5xp2_ASAP7_75t_SL g3686 ( 
.A(n_3519),
.B(n_3468),
.C(n_3277),
.D(n_3366),
.E(n_3254),
.Y(n_3686)
);

OR2x6_ASAP7_75t_L g3687 ( 
.A(n_3552),
.B(n_3264),
.Y(n_3687)
);

AO21x2_ASAP7_75t_L g3688 ( 
.A1(n_3519),
.A2(n_3312),
.B(n_3321),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3604),
.B(n_3334),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_SL g3690 ( 
.A1(n_3515),
.A2(n_3312),
.B1(n_3274),
.B2(n_3339),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3518),
.Y(n_3691)
);

AOI22xp33_ASAP7_75t_L g3692 ( 
.A1(n_3606),
.A2(n_3634),
.B1(n_3625),
.B2(n_3626),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3584),
.B(n_3334),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_R g3694 ( 
.A(n_3586),
.B(n_102),
.Y(n_3694)
);

AOI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3606),
.A2(n_3323),
.B1(n_3329),
.B2(n_3321),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3577),
.Y(n_3696)
);

AOI22xp33_ASAP7_75t_L g3697 ( 
.A1(n_3626),
.A2(n_3602),
.B1(n_3633),
.B2(n_3593),
.Y(n_3697)
);

OR2x2_ASAP7_75t_L g3698 ( 
.A(n_3575),
.B(n_3277),
.Y(n_3698)
);

HB1xp67_ASAP7_75t_L g3699 ( 
.A(n_3573),
.Y(n_3699)
);

OAI221xp5_ASAP7_75t_L g3700 ( 
.A1(n_3614),
.A2(n_3329),
.B1(n_3323),
.B2(n_3345),
.C(n_3336),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3599),
.B(n_3242),
.Y(n_3701)
);

AOI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3609),
.A2(n_3345),
.B(n_3336),
.Y(n_3702)
);

AOI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3602),
.A2(n_3624),
.B1(n_3612),
.B2(n_3629),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3577),
.Y(n_3704)
);

NOR2x1_ASAP7_75t_SL g3705 ( 
.A(n_3526),
.B(n_3242),
.Y(n_3705)
);

CKINVDCx5p33_ASAP7_75t_R g3706 ( 
.A(n_3608),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3536),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3524),
.Y(n_3708)
);

OAI322xp33_ASAP7_75t_L g3709 ( 
.A1(n_3623),
.A2(n_3243),
.A3(n_3249),
.B1(n_3285),
.B2(n_3251),
.C1(n_3257),
.C2(n_3260),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_L g3710 ( 
.A(n_3572),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3536),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3539),
.B(n_3243),
.Y(n_3712)
);

INVxp67_ASAP7_75t_L g3713 ( 
.A(n_3564),
.Y(n_3713)
);

OAI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3608),
.A2(n_3249),
.B1(n_3277),
.B2(n_3237),
.Y(n_3714)
);

OAI221xp5_ASAP7_75t_L g3715 ( 
.A1(n_3632),
.A2(n_3260),
.B1(n_3263),
.B2(n_3257),
.C(n_3251),
.Y(n_3715)
);

AND2x4_ASAP7_75t_L g3716 ( 
.A(n_3526),
.B(n_3236),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3579),
.A2(n_3250),
.B1(n_3220),
.B2(n_3237),
.Y(n_3717)
);

NAND4xp25_ASAP7_75t_L g3718 ( 
.A(n_3568),
.B(n_3285),
.C(n_3263),
.D(n_3238),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3538),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_L g3720 ( 
.A(n_3553),
.B(n_3236),
.Y(n_3720)
);

AOI222xp33_ASAP7_75t_L g3721 ( 
.A1(n_3611),
.A2(n_3616),
.B1(n_3571),
.B2(n_3568),
.C1(n_3601),
.C2(n_3585),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3584),
.B(n_3238),
.Y(n_3722)
);

HB1xp67_ASAP7_75t_L g3723 ( 
.A(n_3543),
.Y(n_3723)
);

AOI221xp5_ASAP7_75t_L g3724 ( 
.A1(n_3611),
.A2(n_3241),
.B1(n_3247),
.B2(n_3252),
.C(n_3244),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3514),
.B(n_3241),
.Y(n_3725)
);

INVxp67_ASAP7_75t_L g3726 ( 
.A(n_3571),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3524),
.Y(n_3727)
);

NOR2x2_ASAP7_75t_L g3728 ( 
.A(n_3534),
.B(n_3244),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3538),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3529),
.B(n_3247),
.Y(n_3730)
);

OAI221xp5_ASAP7_75t_L g3731 ( 
.A1(n_3597),
.A2(n_3277),
.B1(n_3250),
.B2(n_3281),
.C(n_3252),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3579),
.A2(n_3281),
.B1(n_3266),
.B2(n_3269),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_3543),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3534),
.B(n_3265),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3549),
.Y(n_3735)
);

NAND3xp33_ASAP7_75t_L g3736 ( 
.A(n_3600),
.B(n_3220),
.C(n_3250),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3541),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3549),
.Y(n_3738)
);

NOR4xp25_ASAP7_75t_SL g3739 ( 
.A(n_3609),
.B(n_3254),
.C(n_3318),
.D(n_3286),
.Y(n_3739)
);

AND2x4_ASAP7_75t_L g3740 ( 
.A(n_3541),
.B(n_3265),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3551),
.Y(n_3741)
);

AOI221x1_ASAP7_75t_L g3742 ( 
.A1(n_3583),
.A2(n_3269),
.B1(n_3278),
.B2(n_3266),
.C(n_3254),
.Y(n_3742)
);

AOI221xp5_ASAP7_75t_L g3743 ( 
.A1(n_3616),
.A2(n_3278),
.B1(n_107),
.B2(n_103),
.C(n_105),
.Y(n_3743)
);

A2O1A1Ixp33_ASAP7_75t_L g3744 ( 
.A1(n_3583),
.A2(n_3601),
.B(n_3585),
.C(n_3545),
.Y(n_3744)
);

INVx5_ASAP7_75t_SL g3745 ( 
.A(n_3583),
.Y(n_3745)
);

AOI221xp5_ASAP7_75t_L g3746 ( 
.A1(n_3545),
.A2(n_109),
.B1(n_103),
.B2(n_108),
.C(n_110),
.Y(n_3746)
);

NAND2xp33_ASAP7_75t_SL g3747 ( 
.A(n_3613),
.B(n_3254),
.Y(n_3747)
);

NAND3xp33_ASAP7_75t_L g3748 ( 
.A(n_3600),
.B(n_3220),
.C(n_3250),
.Y(n_3748)
);

OAI222xp33_ASAP7_75t_L g3749 ( 
.A1(n_3520),
.A2(n_3254),
.B1(n_3286),
.B2(n_3220),
.C1(n_3253),
.C2(n_117),
.Y(n_3749)
);

NAND4xp75_ASAP7_75t_L g3750 ( 
.A(n_3664),
.B(n_3520),
.C(n_3547),
.D(n_3596),
.Y(n_3750)
);

NAND4xp75_ASAP7_75t_L g3751 ( 
.A(n_3636),
.B(n_3743),
.C(n_3654),
.D(n_3746),
.Y(n_3751)
);

OAI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3654),
.A2(n_3597),
.B(n_3592),
.Y(n_3752)
);

NOR3xp33_ASAP7_75t_SL g3753 ( 
.A(n_3706),
.B(n_3590),
.C(n_3525),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3657),
.B(n_3574),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3657),
.B(n_3574),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3644),
.B(n_3542),
.Y(n_3756)
);

BUFx2_ASAP7_75t_L g3757 ( 
.A(n_3638),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3639),
.B(n_3547),
.Y(n_3758)
);

OR2x2_ASAP7_75t_L g3759 ( 
.A(n_3726),
.B(n_3532),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3661),
.B(n_3535),
.Y(n_3760)
);

AOI211xp5_ASAP7_75t_L g3761 ( 
.A1(n_3637),
.A2(n_3589),
.B(n_3615),
.C(n_3603),
.Y(n_3761)
);

NAND3xp33_ASAP7_75t_L g3762 ( 
.A(n_3746),
.B(n_3589),
.C(n_3628),
.Y(n_3762)
);

NAND4xp75_ASAP7_75t_L g3763 ( 
.A(n_3743),
.B(n_3603),
.C(n_3596),
.D(n_3566),
.Y(n_3763)
);

OA211x2_ASAP7_75t_L g3764 ( 
.A1(n_3713),
.A2(n_3540),
.B(n_3589),
.C(n_3566),
.Y(n_3764)
);

NOR3xp33_ASAP7_75t_L g3765 ( 
.A(n_3660),
.B(n_3631),
.C(n_3595),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3697),
.B(n_3546),
.Y(n_3766)
);

OA21x2_ASAP7_75t_L g3767 ( 
.A1(n_3676),
.A2(n_3582),
.B(n_3561),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3643),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3638),
.B(n_3542),
.Y(n_3769)
);

AO21x2_ASAP7_75t_L g3770 ( 
.A1(n_3744),
.A2(n_3582),
.B(n_3561),
.Y(n_3770)
);

AOI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3647),
.A2(n_3558),
.B1(n_3544),
.B2(n_3556),
.Y(n_3771)
);

AND2x4_ASAP7_75t_L g3772 ( 
.A(n_3638),
.B(n_3544),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3662),
.B(n_3558),
.Y(n_3773)
);

INVx2_ASAP7_75t_SL g3774 ( 
.A(n_3699),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3692),
.B(n_3551),
.Y(n_3775)
);

NAND2x1p5_ASAP7_75t_L g3776 ( 
.A(n_3673),
.B(n_3589),
.Y(n_3776)
);

AND2x2_ASAP7_75t_L g3777 ( 
.A(n_3667),
.B(n_3548),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3721),
.B(n_3555),
.Y(n_3778)
);

NOR3xp33_ASAP7_75t_L g3779 ( 
.A(n_3684),
.B(n_3631),
.C(n_3587),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3652),
.A2(n_3589),
.B1(n_3540),
.B2(n_3569),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3650),
.Y(n_3781)
);

AND2x2_ASAP7_75t_SL g3782 ( 
.A(n_3649),
.B(n_3540),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3678),
.B(n_3679),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3723),
.Y(n_3784)
);

OR2x2_ASAP7_75t_L g3785 ( 
.A(n_3673),
.B(n_3682),
.Y(n_3785)
);

OR2x6_ASAP7_75t_L g3786 ( 
.A(n_3737),
.B(n_3587),
.Y(n_3786)
);

OR2x2_ASAP7_75t_L g3787 ( 
.A(n_3682),
.B(n_3570),
.Y(n_3787)
);

NAND4xp75_ASAP7_75t_L g3788 ( 
.A(n_3742),
.B(n_3610),
.C(n_3605),
.D(n_3556),
.Y(n_3788)
);

NAND3xp33_ASAP7_75t_L g3789 ( 
.A(n_3649),
.B(n_3615),
.C(n_3610),
.Y(n_3789)
);

AOI22xp33_ASAP7_75t_L g3790 ( 
.A1(n_3652),
.A2(n_3641),
.B1(n_3684),
.B2(n_3656),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_3721),
.A2(n_3557),
.B1(n_3548),
.B2(n_3510),
.Y(n_3791)
);

NAND3xp33_ASAP7_75t_L g3792 ( 
.A(n_3703),
.B(n_3605),
.C(n_3570),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3710),
.B(n_3555),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3640),
.Y(n_3794)
);

OR2x2_ASAP7_75t_L g3795 ( 
.A(n_3718),
.B(n_3701),
.Y(n_3795)
);

NOR2xp33_ASAP7_75t_L g3796 ( 
.A(n_3672),
.B(n_3663),
.Y(n_3796)
);

NOR3xp33_ASAP7_75t_L g3797 ( 
.A(n_3749),
.B(n_3560),
.C(n_3559),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3733),
.Y(n_3798)
);

OAI211xp5_ASAP7_75t_SL g3799 ( 
.A1(n_3690),
.A2(n_3560),
.B(n_3563),
.C(n_3559),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_3701),
.B(n_3563),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3708),
.B(n_3510),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3727),
.B(n_3745),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3745),
.B(n_3557),
.Y(n_3803)
);

HB1xp67_ASAP7_75t_L g3804 ( 
.A(n_3640),
.Y(n_3804)
);

OR2x2_ASAP7_75t_L g3805 ( 
.A(n_3712),
.B(n_3550),
.Y(n_3805)
);

NAND3xp33_ASAP7_75t_L g3806 ( 
.A(n_3685),
.B(n_3581),
.C(n_3550),
.Y(n_3806)
);

HB1xp67_ASAP7_75t_L g3807 ( 
.A(n_3658),
.Y(n_3807)
);

NOR3xp33_ASAP7_75t_L g3808 ( 
.A(n_3646),
.B(n_3523),
.C(n_3517),
.Y(n_3808)
);

XNOR2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3694),
.B(n_3732),
.Y(n_3809)
);

OA211x2_ASAP7_75t_L g3810 ( 
.A1(n_3685),
.A2(n_3517),
.B(n_3528),
.C(n_3523),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3716),
.B(n_3528),
.Y(n_3811)
);

AOI211xp5_ASAP7_75t_L g3812 ( 
.A1(n_3714),
.A2(n_3581),
.B(n_3578),
.C(n_3533),
.Y(n_3812)
);

OR2x2_ASAP7_75t_L g3813 ( 
.A(n_3712),
.B(n_3578),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3645),
.Y(n_3814)
);

OR2x2_ASAP7_75t_L g3815 ( 
.A(n_3698),
.B(n_3533),
.Y(n_3815)
);

NOR3xp33_ASAP7_75t_L g3816 ( 
.A(n_3648),
.B(n_111),
.C(n_113),
.Y(n_3816)
);

OAI22xp33_ASAP7_75t_L g3817 ( 
.A1(n_3642),
.A2(n_3253),
.B1(n_3254),
.B2(n_2880),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_SL g3818 ( 
.A(n_3745),
.B(n_3747),
.Y(n_3818)
);

NAND3xp33_ASAP7_75t_L g3819 ( 
.A(n_3731),
.B(n_111),
.C(n_115),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3659),
.Y(n_3820)
);

AO21x1_ASAP7_75t_SL g3821 ( 
.A1(n_3665),
.A2(n_116),
.B(n_117),
.Y(n_3821)
);

OR2x2_ASAP7_75t_SL g3822 ( 
.A(n_3680),
.B(n_3253),
.Y(n_3822)
);

NAND3xp33_ASAP7_75t_L g3823 ( 
.A(n_3731),
.B(n_116),
.C(n_119),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3716),
.B(n_120),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3720),
.B(n_120),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3666),
.Y(n_3826)
);

NAND3xp33_ASAP7_75t_L g3827 ( 
.A(n_3675),
.B(n_121),
.C(n_123),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3688),
.A2(n_3253),
.B1(n_1021),
.B2(n_1045),
.Y(n_3828)
);

OR2x2_ASAP7_75t_L g3829 ( 
.A(n_3671),
.B(n_121),
.Y(n_3829)
);

AOI22xp33_ASAP7_75t_L g3830 ( 
.A1(n_3688),
.A2(n_1021),
.B1(n_1045),
.B2(n_1032),
.Y(n_3830)
);

AOI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3681),
.A2(n_3700),
.B1(n_3677),
.B2(n_3696),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3651),
.B(n_123),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3669),
.B(n_124),
.Y(n_3833)
);

INVx2_ASAP7_75t_L g3834 ( 
.A(n_3658),
.Y(n_3834)
);

NAND4xp25_ASAP7_75t_L g3835 ( 
.A(n_3717),
.B(n_126),
.C(n_124),
.D(n_125),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3655),
.B(n_126),
.Y(n_3836)
);

OA211x2_ASAP7_75t_L g3837 ( 
.A1(n_3675),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_3837)
);

OAI211xp5_ASAP7_75t_L g3838 ( 
.A1(n_3739),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3689),
.B(n_130),
.Y(n_3839)
);

NAND3xp33_ASAP7_75t_L g3840 ( 
.A(n_3668),
.B(n_130),
.C(n_131),
.Y(n_3840)
);

NAND3xp33_ASAP7_75t_L g3841 ( 
.A(n_3670),
.B(n_131),
.C(n_132),
.Y(n_3841)
);

OR2x2_ASAP7_75t_L g3842 ( 
.A(n_3785),
.B(n_3674),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_SL g3843 ( 
.A(n_3782),
.B(n_3752),
.Y(n_3843)
);

HB1xp67_ASAP7_75t_L g3844 ( 
.A(n_3786),
.Y(n_3844)
);

AOI221xp5_ASAP7_75t_L g3845 ( 
.A1(n_3790),
.A2(n_3700),
.B1(n_3709),
.B2(n_3748),
.C(n_3736),
.Y(n_3845)
);

NOR2xp33_ASAP7_75t_L g3846 ( 
.A(n_3751),
.B(n_3758),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_SL g3847 ( 
.A(n_3754),
.B(n_3681),
.Y(n_3847)
);

OAI221xp5_ASAP7_75t_L g3848 ( 
.A1(n_3796),
.A2(n_3695),
.B1(n_3642),
.B2(n_3704),
.C(n_3724),
.Y(n_3848)
);

INVx1_ASAP7_75t_SL g3849 ( 
.A(n_3757),
.Y(n_3849)
);

BUFx2_ASAP7_75t_L g3850 ( 
.A(n_3770),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3769),
.B(n_3705),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3804),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3770),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3772),
.B(n_3722),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3807),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3768),
.Y(n_3856)
);

HB1xp67_ASAP7_75t_L g3857 ( 
.A(n_3786),
.Y(n_3857)
);

OAI31xp33_ASAP7_75t_L g3858 ( 
.A1(n_3762),
.A2(n_3838),
.A3(n_3799),
.B(n_3823),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3772),
.B(n_3693),
.Y(n_3859)
);

AOI221xp5_ASAP7_75t_L g3860 ( 
.A1(n_3762),
.A2(n_3715),
.B1(n_3724),
.B2(n_3738),
.C(n_3735),
.Y(n_3860)
);

INVx1_ASAP7_75t_SL g3861 ( 
.A(n_3755),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3776),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3803),
.B(n_3734),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3786),
.Y(n_3864)
);

AOI221xp5_ASAP7_75t_L g3865 ( 
.A1(n_3765),
.A2(n_3715),
.B1(n_3741),
.B2(n_3711),
.C(n_3707),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3774),
.B(n_3683),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3781),
.Y(n_3867)
);

NOR3xp33_ASAP7_75t_SL g3868 ( 
.A(n_3750),
.B(n_3719),
.C(n_3691),
.Y(n_3868)
);

AOI221xp5_ASAP7_75t_L g3869 ( 
.A1(n_3761),
.A2(n_3729),
.B1(n_3732),
.B2(n_3730),
.C(n_3725),
.Y(n_3869)
);

INVxp67_ASAP7_75t_L g3870 ( 
.A(n_3821),
.Y(n_3870)
);

OAI221xp5_ASAP7_75t_SL g3871 ( 
.A1(n_3780),
.A2(n_3761),
.B1(n_3778),
.B2(n_3779),
.C(n_3831),
.Y(n_3871)
);

NAND4xp25_ASAP7_75t_SL g3872 ( 
.A(n_3789),
.B(n_3686),
.C(n_3728),
.D(n_3725),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3784),
.B(n_3734),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3798),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3814),
.Y(n_3875)
);

AOI22xp33_ASAP7_75t_L g3876 ( 
.A1(n_3810),
.A2(n_3642),
.B1(n_3740),
.B2(n_3687),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3767),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3820),
.Y(n_3878)
);

INVx3_ASAP7_75t_L g3879 ( 
.A(n_3767),
.Y(n_3879)
);

OAI221xp5_ASAP7_75t_L g3880 ( 
.A1(n_3753),
.A2(n_3687),
.B1(n_3730),
.B2(n_3702),
.C(n_3653),
.Y(n_3880)
);

AOI211xp5_ASAP7_75t_SL g3881 ( 
.A1(n_3812),
.A2(n_3740),
.B(n_3687),
.C(n_134),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3788),
.Y(n_3882)
);

BUFx2_ASAP7_75t_L g3883 ( 
.A(n_3809),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3794),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3775),
.B(n_132),
.Y(n_3885)
);

AND2x4_ASAP7_75t_L g3886 ( 
.A(n_3834),
.B(n_133),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3826),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3822),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3793),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3773),
.Y(n_3890)
);

NAND2xp33_ASAP7_75t_SL g3891 ( 
.A(n_3766),
.B(n_133),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3756),
.B(n_134),
.Y(n_3892)
);

INVx3_ASAP7_75t_L g3893 ( 
.A(n_3763),
.Y(n_3893)
);

NAND4xp25_ASAP7_75t_L g3894 ( 
.A(n_3764),
.B(n_137),
.C(n_135),
.D(n_136),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3777),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3802),
.B(n_135),
.Y(n_3896)
);

AND2x2_ASAP7_75t_L g3897 ( 
.A(n_3771),
.B(n_3791),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3783),
.B(n_138),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3815),
.Y(n_3899)
);

BUFx3_ASAP7_75t_L g3900 ( 
.A(n_3833),
.Y(n_3900)
);

OR2x2_ASAP7_75t_L g3901 ( 
.A(n_3829),
.B(n_138),
.Y(n_3901)
);

INVx2_ASAP7_75t_SL g3902 ( 
.A(n_3801),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3797),
.B(n_139),
.Y(n_3903)
);

AND2x4_ASAP7_75t_SL g3904 ( 
.A(n_3839),
.B(n_139),
.Y(n_3904)
);

NAND3xp33_ASAP7_75t_L g3905 ( 
.A(n_3819),
.B(n_140),
.C(n_141),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3818),
.B(n_141),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3759),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3808),
.B(n_142),
.Y(n_3908)
);

BUFx2_ASAP7_75t_L g3909 ( 
.A(n_3827),
.Y(n_3909)
);

INVx3_ASAP7_75t_L g3910 ( 
.A(n_3813),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3832),
.Y(n_3911)
);

OR2x2_ASAP7_75t_L g3912 ( 
.A(n_3795),
.B(n_143),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3824),
.Y(n_3913)
);

HB1xp67_ASAP7_75t_L g3914 ( 
.A(n_3760),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3819),
.A2(n_995),
.B1(n_1032),
.B2(n_1021),
.Y(n_3915)
);

BUFx2_ASAP7_75t_L g3916 ( 
.A(n_3827),
.Y(n_3916)
);

HB1xp67_ASAP7_75t_L g3917 ( 
.A(n_3811),
.Y(n_3917)
);

AOI22xp33_ASAP7_75t_L g3918 ( 
.A1(n_3823),
.A2(n_995),
.B1(n_1045),
.B2(n_1032),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3805),
.Y(n_3919)
);

AOI221xp5_ASAP7_75t_L g3920 ( 
.A1(n_3789),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.C(n_148),
.Y(n_3920)
);

OAI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3841),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3836),
.B(n_150),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3800),
.Y(n_3923)
);

AND2x4_ASAP7_75t_L g3924 ( 
.A(n_3841),
.B(n_151),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3787),
.Y(n_3925)
);

OAI31xp33_ASAP7_75t_L g3926 ( 
.A1(n_3792),
.A2(n_153),
.A3(n_151),
.B(n_152),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3812),
.B(n_155),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3825),
.B(n_155),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3792),
.B(n_156),
.Y(n_3929)
);

AOI221xp5_ASAP7_75t_L g3930 ( 
.A1(n_3835),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.C(n_159),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3840),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3806),
.Y(n_3932)
);

OR2x2_ASAP7_75t_L g3933 ( 
.A(n_3806),
.B(n_3830),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3864),
.Y(n_3934)
);

AOI22xp33_ASAP7_75t_L g3935 ( 
.A1(n_3843),
.A2(n_3816),
.B1(n_3837),
.B2(n_3817),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3859),
.B(n_3828),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3924),
.B(n_3883),
.Y(n_3937)
);

HB1xp67_ASAP7_75t_L g3938 ( 
.A(n_3850),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3850),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3844),
.Y(n_3940)
);

OAI322xp33_ASAP7_75t_L g3941 ( 
.A1(n_3932),
.A2(n_157),
.A3(n_159),
.B1(n_160),
.B2(n_163),
.C1(n_164),
.C2(n_165),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3924),
.B(n_160),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3864),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3857),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3902),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3870),
.Y(n_3946)
);

OAI322xp33_ASAP7_75t_L g3947 ( 
.A1(n_3893),
.A2(n_164),
.A3(n_166),
.B1(n_167),
.B2(n_168),
.C1(n_169),
.C2(n_170),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3924),
.B(n_3883),
.Y(n_3948)
);

AOI32xp33_ASAP7_75t_L g3949 ( 
.A1(n_3893),
.A2(n_166),
.A3(n_168),
.B1(n_170),
.B2(n_172),
.Y(n_3949)
);

NOR2x1p5_ASAP7_75t_SL g3950 ( 
.A(n_3853),
.B(n_172),
.Y(n_3950)
);

AND2x4_ASAP7_75t_L g3951 ( 
.A(n_3902),
.B(n_174),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3852),
.Y(n_3952)
);

OAI21xp33_ASAP7_75t_L g3953 ( 
.A1(n_3868),
.A2(n_174),
.B(n_175),
.Y(n_3953)
);

AOI32xp33_ASAP7_75t_L g3954 ( 
.A1(n_3893),
.A2(n_176),
.A3(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_3954)
);

AND2x2_ASAP7_75t_L g3955 ( 
.A(n_3859),
.B(n_177),
.Y(n_3955)
);

INVx1_ASAP7_75t_SL g3956 ( 
.A(n_3849),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3903),
.B(n_178),
.Y(n_3957)
);

OR2x2_ASAP7_75t_L g3958 ( 
.A(n_3912),
.B(n_179),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3900),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3855),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3892),
.Y(n_3961)
);

NAND4xp25_ASAP7_75t_L g3962 ( 
.A(n_3846),
.B(n_181),
.C(n_182),
.D(n_183),
.Y(n_3962)
);

OA222x2_ASAP7_75t_L g3963 ( 
.A1(n_3853),
.A2(n_181),
.B1(n_182),
.B2(n_184),
.C1(n_185),
.C2(n_186),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3854),
.B(n_184),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3892),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3900),
.Y(n_3966)
);

BUFx3_ASAP7_75t_L g3967 ( 
.A(n_3904),
.Y(n_3967)
);

AND2x4_ASAP7_75t_L g3968 ( 
.A(n_3884),
.B(n_185),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3910),
.Y(n_3969)
);

NAND2x1p5_ASAP7_75t_L g3970 ( 
.A(n_3843),
.B(n_187),
.Y(n_3970)
);

OAI21xp33_ASAP7_75t_L g3971 ( 
.A1(n_3871),
.A2(n_188),
.B(n_189),
.Y(n_3971)
);

OAI322xp33_ASAP7_75t_L g3972 ( 
.A1(n_3909),
.A2(n_188),
.A3(n_189),
.B1(n_190),
.B2(n_191),
.C1(n_192),
.C2(n_193),
.Y(n_3972)
);

INVx1_ASAP7_75t_SL g3973 ( 
.A(n_3851),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3854),
.B(n_190),
.Y(n_3974)
);

NAND4xp25_ASAP7_75t_L g3975 ( 
.A(n_3858),
.B(n_193),
.C(n_194),
.D(n_195),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3903),
.B(n_197),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3863),
.B(n_199),
.Y(n_3977)
);

OR2x2_ASAP7_75t_L g3978 ( 
.A(n_3912),
.B(n_199),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3863),
.B(n_3896),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3909),
.B(n_200),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3896),
.B(n_201),
.Y(n_3981)
);

OR2x2_ASAP7_75t_L g3982 ( 
.A(n_3890),
.B(n_201),
.Y(n_3982)
);

AOI22xp5_ASAP7_75t_L g3983 ( 
.A1(n_3916),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_3983)
);

NAND4xp75_ASAP7_75t_L g3984 ( 
.A(n_3926),
.B(n_203),
.C(n_205),
.D(n_206),
.Y(n_3984)
);

AOI211xp5_ASAP7_75t_SL g3985 ( 
.A1(n_3848),
.A2(n_207),
.B(n_210),
.C(n_211),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3862),
.Y(n_3986)
);

AOI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3916),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_3987)
);

INVxp67_ASAP7_75t_SL g3988 ( 
.A(n_3879),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3898),
.B(n_213),
.Y(n_3989)
);

NAND2x1p5_ASAP7_75t_L g3990 ( 
.A(n_3898),
.B(n_213),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3890),
.B(n_3842),
.Y(n_3991)
);

OA222x2_ASAP7_75t_L g3992 ( 
.A1(n_3879),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.C1(n_217),
.C2(n_219),
.Y(n_3992)
);

O2A1O1Ixp33_ASAP7_75t_L g3993 ( 
.A1(n_3882),
.A2(n_214),
.B(n_215),
.C(n_216),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3862),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3910),
.Y(n_3995)
);

AOI32xp33_ASAP7_75t_L g3996 ( 
.A1(n_3927),
.A2(n_217),
.A3(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3910),
.Y(n_3997)
);

INVx1_ASAP7_75t_SL g3998 ( 
.A(n_3851),
.Y(n_3998)
);

OR2x2_ASAP7_75t_L g3999 ( 
.A(n_3842),
.B(n_220),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3901),
.Y(n_4000)
);

OAI22xp5_ASAP7_75t_L g4001 ( 
.A1(n_3905),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3886),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3901),
.Y(n_4003)
);

OR2x2_ASAP7_75t_L g4004 ( 
.A(n_3861),
.B(n_224),
.Y(n_4004)
);

AND2x2_ASAP7_75t_L g4005 ( 
.A(n_3895),
.B(n_3906),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3907),
.Y(n_4006)
);

NOR2xp33_ASAP7_75t_L g4007 ( 
.A(n_3931),
.B(n_225),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3907),
.Y(n_4008)
);

INVx2_ASAP7_75t_L g4009 ( 
.A(n_3886),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3895),
.B(n_226),
.Y(n_4010)
);

INVx2_ASAP7_75t_SL g4011 ( 
.A(n_3898),
.Y(n_4011)
);

OR2x2_ASAP7_75t_L g4012 ( 
.A(n_3885),
.B(n_226),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3899),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3929),
.B(n_228),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3899),
.Y(n_4015)
);

OAI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3881),
.A2(n_229),
.B(n_230),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3906),
.B(n_3847),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3917),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3884),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_SL g4020 ( 
.A(n_3845),
.B(n_229),
.Y(n_4020)
);

NAND2x1_ASAP7_75t_L g4021 ( 
.A(n_3886),
.B(n_231),
.Y(n_4021)
);

XNOR2x1_ASAP7_75t_L g4022 ( 
.A(n_3897),
.B(n_231),
.Y(n_4022)
);

AOI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_3894),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_4023)
);

OR2x2_ASAP7_75t_L g4024 ( 
.A(n_3937),
.B(n_3885),
.Y(n_4024)
);

NAND3xp33_ASAP7_75t_L g4025 ( 
.A(n_3985),
.B(n_3882),
.C(n_3927),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3946),
.B(n_3919),
.Y(n_4026)
);

INVx2_ASAP7_75t_SL g4027 ( 
.A(n_3967),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3990),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_4021),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3951),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3979),
.B(n_4017),
.Y(n_4031)
);

OR2x2_ASAP7_75t_L g4032 ( 
.A(n_3948),
.B(n_3919),
.Y(n_4032)
);

AND2x4_ASAP7_75t_L g4033 ( 
.A(n_3969),
.B(n_3856),
.Y(n_4033)
);

NOR3xp33_ASAP7_75t_L g4034 ( 
.A(n_3975),
.B(n_3891),
.C(n_3929),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3951),
.Y(n_4035)
);

AOI33xp33_ASAP7_75t_L g4036 ( 
.A1(n_3935),
.A2(n_3897),
.A3(n_3956),
.B1(n_3998),
.B2(n_3973),
.B3(n_3923),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_4005),
.B(n_3914),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_SL g4038 ( 
.A(n_4011),
.B(n_3891),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3995),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3953),
.B(n_3908),
.Y(n_4040)
);

OR2x6_ASAP7_75t_L g4041 ( 
.A(n_3970),
.B(n_3980),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3988),
.Y(n_4042)
);

OR2x2_ASAP7_75t_L g4043 ( 
.A(n_3991),
.B(n_3873),
.Y(n_4043)
);

NOR2xp33_ASAP7_75t_SL g4044 ( 
.A(n_3947),
.B(n_3975),
.Y(n_4044)
);

NAND2x1_ASAP7_75t_L g4045 ( 
.A(n_4002),
.B(n_3879),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_L g4046 ( 
.A(n_3953),
.B(n_3997),
.Y(n_4046)
);

NOR2xp33_ASAP7_75t_L g4047 ( 
.A(n_3971),
.B(n_3959),
.Y(n_4047)
);

NAND2xp33_ASAP7_75t_SL g4048 ( 
.A(n_4022),
.B(n_3921),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3950),
.B(n_3908),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3938),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3966),
.B(n_3925),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3971),
.B(n_3867),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3977),
.B(n_3911),
.Y(n_4053)
);

INVxp67_ASAP7_75t_SL g4054 ( 
.A(n_3939),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3961),
.B(n_3913),
.Y(n_4055)
);

AND2x2_ASAP7_75t_L g4056 ( 
.A(n_3965),
.B(n_3913),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3955),
.B(n_3928),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3981),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3945),
.Y(n_4059)
);

NAND3xp33_ASAP7_75t_L g4060 ( 
.A(n_4020),
.B(n_3920),
.C(n_3860),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3964),
.B(n_3928),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3940),
.Y(n_4062)
);

NAND2xp33_ASAP7_75t_R g4063 ( 
.A(n_4016),
.B(n_3933),
.Y(n_4063)
);

AND2x4_ASAP7_75t_SL g4064 ( 
.A(n_4009),
.B(n_3874),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_L g4065 ( 
.A(n_3957),
.B(n_3889),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3944),
.Y(n_4066)
);

NOR2x1_ASAP7_75t_L g4067 ( 
.A(n_3947),
.B(n_3877),
.Y(n_4067)
);

AND2x4_ASAP7_75t_L g4068 ( 
.A(n_4000),
.B(n_3866),
.Y(n_4068)
);

NOR3xp33_ASAP7_75t_SL g4069 ( 
.A(n_4018),
.B(n_3880),
.C(n_3872),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3968),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3968),
.Y(n_4071)
);

BUFx2_ASAP7_75t_L g4072 ( 
.A(n_4003),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3989),
.Y(n_4073)
);

HB1xp67_ASAP7_75t_L g4074 ( 
.A(n_4006),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3974),
.Y(n_4075)
);

OR2x2_ASAP7_75t_L g4076 ( 
.A(n_3986),
.B(n_3933),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_3994),
.B(n_3904),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3934),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3943),
.B(n_3875),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3999),
.Y(n_4080)
);

AO21x1_ASAP7_75t_L g4081 ( 
.A1(n_3993),
.A2(n_3877),
.B(n_3878),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_4010),
.Y(n_4082)
);

NOR4xp25_ASAP7_75t_SL g4083 ( 
.A(n_4013),
.B(n_3869),
.C(n_3865),
.D(n_3887),
.Y(n_4083)
);

OR2x2_ASAP7_75t_L g4084 ( 
.A(n_4015),
.B(n_3922),
.Y(n_4084)
);

OR2x2_ASAP7_75t_L g4085 ( 
.A(n_4008),
.B(n_3888),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3982),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3958),
.Y(n_4087)
);

NAND4xp25_ASAP7_75t_L g4088 ( 
.A(n_4007),
.B(n_3930),
.C(n_3918),
.D(n_3915),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3936),
.B(n_3888),
.Y(n_4089)
);

NAND2xp33_ASAP7_75t_L g4090 ( 
.A(n_3984),
.B(n_3876),
.Y(n_4090)
);

OR2x2_ASAP7_75t_L g4091 ( 
.A(n_4004),
.B(n_3952),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3949),
.B(n_232),
.Y(n_4092)
);

BUFx2_ASAP7_75t_L g4093 ( 
.A(n_3978),
.Y(n_4093)
);

AO21x1_ASAP7_75t_L g4094 ( 
.A1(n_3976),
.A2(n_234),
.B(n_235),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3960),
.B(n_235),
.Y(n_4095)
);

BUFx2_ASAP7_75t_L g4096 ( 
.A(n_4012),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_4019),
.Y(n_4097)
);

BUFx2_ASAP7_75t_L g4098 ( 
.A(n_3942),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3954),
.B(n_237),
.Y(n_4099)
);

NOR3xp33_ASAP7_75t_L g4100 ( 
.A(n_3962),
.B(n_238),
.C(n_240),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3996),
.B(n_240),
.Y(n_4101)
);

OR2x2_ASAP7_75t_L g4102 ( 
.A(n_4014),
.B(n_241),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3963),
.B(n_242),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_4023),
.B(n_243),
.Y(n_4104)
);

OAI221xp5_ASAP7_75t_L g4105 ( 
.A1(n_4023),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.C(n_246),
.Y(n_4105)
);

NOR3xp33_ASAP7_75t_L g4106 ( 
.A(n_3962),
.B(n_244),
.C(n_246),
.Y(n_4106)
);

AOI221xp5_ASAP7_75t_L g4107 ( 
.A1(n_3972),
.A2(n_3941),
.B1(n_4001),
.B2(n_3987),
.C(n_3983),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_4031),
.B(n_3983),
.Y(n_4108)
);

OR2x2_ASAP7_75t_L g4109 ( 
.A(n_4030),
.B(n_3987),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_4026),
.B(n_3963),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4027),
.B(n_3992),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_4035),
.B(n_3992),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_4057),
.B(n_3941),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4034),
.B(n_3972),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_4045),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_4034),
.B(n_4029),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_4061),
.B(n_248),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_4072),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_4100),
.B(n_250),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_4037),
.B(n_251),
.Y(n_4120)
);

INVx1_ASAP7_75t_SL g4121 ( 
.A(n_4064),
.Y(n_4121)
);

OR2x2_ASAP7_75t_L g4122 ( 
.A(n_4046),
.B(n_252),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_4060),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_4123)
);

NOR2x1_ASAP7_75t_L g4124 ( 
.A(n_4103),
.B(n_4025),
.Y(n_4124)
);

OR2x2_ASAP7_75t_L g4125 ( 
.A(n_4046),
.B(n_253),
.Y(n_4125)
);

NOR2x1_ASAP7_75t_L g4126 ( 
.A(n_4032),
.B(n_255),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_4077),
.Y(n_4127)
);

AOI22xp33_ASAP7_75t_SL g4128 ( 
.A1(n_4044),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_4128)
);

INVxp67_ASAP7_75t_L g4129 ( 
.A(n_4074),
.Y(n_4129)
);

OR2x2_ASAP7_75t_L g4130 ( 
.A(n_4040),
.B(n_256),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4074),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_4100),
.B(n_258),
.Y(n_4132)
);

OAI21xp5_ASAP7_75t_L g4133 ( 
.A1(n_4067),
.A2(n_259),
.B(n_260),
.Y(n_4133)
);

OAI21xp33_ASAP7_75t_L g4134 ( 
.A1(n_4044),
.A2(n_260),
.B(n_261),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4106),
.B(n_261),
.Y(n_4135)
);

OAI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_4069),
.A2(n_262),
.B(n_263),
.Y(n_4136)
);

AND2x2_ASAP7_75t_SL g4137 ( 
.A(n_4106),
.B(n_4036),
.Y(n_4137)
);

INVx1_ASAP7_75t_SL g4138 ( 
.A(n_4038),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4089),
.B(n_262),
.Y(n_4139)
);

O2A1O1Ixp33_ASAP7_75t_L g4140 ( 
.A1(n_4081),
.A2(n_263),
.B(n_264),
.C(n_265),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_4028),
.B(n_265),
.Y(n_4141)
);

OAI21xp5_ASAP7_75t_L g4142 ( 
.A1(n_4069),
.A2(n_266),
.B(n_267),
.Y(n_4142)
);

NOR3xp33_ASAP7_75t_SL g4143 ( 
.A(n_4063),
.B(n_266),
.C(n_267),
.Y(n_4143)
);

AOI211x1_ASAP7_75t_L g4144 ( 
.A1(n_4094),
.A2(n_269),
.B(n_270),
.C(n_271),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4054),
.Y(n_4145)
);

HB1xp67_ASAP7_75t_L g4146 ( 
.A(n_4041),
.Y(n_4146)
);

NOR2xp67_ASAP7_75t_SL g4147 ( 
.A(n_4024),
.B(n_269),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_4049),
.B(n_270),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_4070),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4054),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_4071),
.B(n_271),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4085),
.Y(n_4152)
);

OR2x2_ASAP7_75t_L g4153 ( 
.A(n_4040),
.B(n_274),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4047),
.B(n_274),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_4051),
.B(n_276),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4047),
.B(n_277),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_4075),
.B(n_277),
.Y(n_4157)
);

NAND4xp75_ASAP7_75t_L g4158 ( 
.A(n_4042),
.B(n_278),
.C(n_279),
.D(n_280),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_4041),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_4041),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_4053),
.B(n_278),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4107),
.B(n_279),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4096),
.Y(n_4163)
);

OR2x2_ASAP7_75t_L g4164 ( 
.A(n_4049),
.B(n_280),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4093),
.Y(n_4165)
);

NOR3xp33_ASAP7_75t_L g4166 ( 
.A(n_4048),
.B(n_4104),
.C(n_4101),
.Y(n_4166)
);

NOR2xp33_ASAP7_75t_L g4167 ( 
.A(n_4058),
.B(n_281),
.Y(n_4167)
);

INVxp67_ASAP7_75t_SL g4168 ( 
.A(n_4104),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_SL g4169 ( 
.A(n_4107),
.B(n_281),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_SL g4170 ( 
.A(n_4068),
.B(n_282),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_4068),
.B(n_283),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_4033),
.Y(n_4172)
);

OAI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_4083),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_4173)
);

OAI31xp33_ASAP7_75t_L g4174 ( 
.A1(n_4105),
.A2(n_286),
.A3(n_287),
.B(n_288),
.Y(n_4174)
);

OAI22xp33_ASAP7_75t_L g4175 ( 
.A1(n_4173),
.A2(n_4052),
.B1(n_4076),
.B2(n_4092),
.Y(n_4175)
);

OAI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_4140),
.A2(n_4090),
.B(n_4052),
.Y(n_4176)
);

OAI21xp33_ASAP7_75t_SL g4177 ( 
.A1(n_4169),
.A2(n_4050),
.B(n_4056),
.Y(n_4177)
);

AOI222xp33_ASAP7_75t_L g4178 ( 
.A1(n_4169),
.A2(n_4066),
.B1(n_4062),
.B2(n_4065),
.C1(n_4098),
.C2(n_4059),
.Y(n_4178)
);

AOI322xp5_ASAP7_75t_L g4179 ( 
.A1(n_4137),
.A2(n_4099),
.A3(n_4092),
.B1(n_4101),
.B2(n_4078),
.C1(n_4082),
.C2(n_4079),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4145),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_4162),
.A2(n_4043),
.B1(n_4099),
.B2(n_4105),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4121),
.B(n_4033),
.Y(n_4182)
);

NOR2xp33_ASAP7_75t_L g4183 ( 
.A(n_4138),
.B(n_4080),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4113),
.B(n_4124),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4110),
.B(n_4055),
.Y(n_4185)
);

OR2x2_ASAP7_75t_L g4186 ( 
.A(n_4118),
.B(n_4091),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_4128),
.B(n_4039),
.Y(n_4187)
);

OAI22xp5_ASAP7_75t_L g4188 ( 
.A1(n_4128),
.A2(n_4087),
.B1(n_4084),
.B2(n_4086),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4150),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_4172),
.B(n_4095),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4172),
.Y(n_4191)
);

AND2x2_ASAP7_75t_SL g4192 ( 
.A(n_4166),
.B(n_4073),
.Y(n_4192)
);

CKINVDCx8_ASAP7_75t_R g4193 ( 
.A(n_4148),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4146),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_SL g4195 ( 
.A(n_4118),
.B(n_4102),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_SL g4196 ( 
.A(n_4144),
.B(n_4097),
.Y(n_4196)
);

OAI332xp33_ASAP7_75t_L g4197 ( 
.A1(n_4114),
.A2(n_4088),
.A3(n_290),
.B1(n_291),
.B2(n_292),
.B3(n_293),
.C1(n_294),
.C2(n_295),
.Y(n_4197)
);

AOI22xp5_ASAP7_75t_L g4198 ( 
.A1(n_4137),
.A2(n_4088),
.B1(n_290),
.B2(n_295),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4146),
.Y(n_4199)
);

OAI21xp5_ASAP7_75t_SL g4200 ( 
.A1(n_4136),
.A2(n_4142),
.B(n_4133),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4129),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4129),
.Y(n_4202)
);

OAI21xp33_ASAP7_75t_SL g4203 ( 
.A1(n_4131),
.A2(n_287),
.B(n_296),
.Y(n_4203)
);

OAI22xp5_ASAP7_75t_L g4204 ( 
.A1(n_4123),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4126),
.Y(n_4205)
);

OA21x2_ASAP7_75t_L g4206 ( 
.A1(n_4170),
.A2(n_297),
.B(n_299),
.Y(n_4206)
);

OR2x2_ASAP7_75t_L g4207 ( 
.A(n_4108),
.B(n_300),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_L g4208 ( 
.A(n_4134),
.B(n_300),
.Y(n_4208)
);

INVxp67_ASAP7_75t_L g4209 ( 
.A(n_4147),
.Y(n_4209)
);

INVxp33_ASAP7_75t_L g4210 ( 
.A(n_4116),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4139),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4120),
.Y(n_4212)
);

OAI21xp5_ASAP7_75t_L g4213 ( 
.A1(n_4143),
.A2(n_301),
.B(n_302),
.Y(n_4213)
);

AOI22xp33_ASAP7_75t_SL g4214 ( 
.A1(n_4163),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4127),
.B(n_303),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_SL g4216 ( 
.A(n_4143),
.B(n_4152),
.Y(n_4216)
);

INVxp67_ASAP7_75t_SL g4217 ( 
.A(n_4115),
.Y(n_4217)
);

XNOR2xp5_ASAP7_75t_L g4218 ( 
.A(n_4166),
.B(n_304),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4115),
.Y(n_4219)
);

OR2x2_ASAP7_75t_L g4220 ( 
.A(n_4109),
.B(n_305),
.Y(n_4220)
);

NAND4xp25_ASAP7_75t_SL g4221 ( 
.A(n_4111),
.B(n_305),
.C(n_306),
.D(n_308),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4149),
.B(n_309),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_4149),
.B(n_309),
.Y(n_4223)
);

AOI21xp33_ASAP7_75t_L g4224 ( 
.A1(n_4165),
.A2(n_310),
.B(n_311),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4148),
.B(n_312),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4117),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4161),
.B(n_4155),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4164),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4170),
.Y(n_4229)
);

AOI21xp33_ASAP7_75t_SL g4230 ( 
.A1(n_4112),
.A2(n_312),
.B(n_313),
.Y(n_4230)
);

NAND4xp25_ASAP7_75t_L g4231 ( 
.A(n_4159),
.B(n_313),
.C(n_314),
.D(n_315),
.Y(n_4231)
);

INVx1_ASAP7_75t_SL g4232 ( 
.A(n_4130),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4168),
.B(n_314),
.Y(n_4233)
);

AND3x1_ASAP7_75t_L g4234 ( 
.A(n_4174),
.B(n_315),
.C(n_316),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_4123),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_4119),
.A2(n_318),
.B(n_319),
.Y(n_4236)
);

NAND3xp33_ASAP7_75t_SL g4237 ( 
.A(n_4159),
.B(n_319),
.C(n_321),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_4160),
.B(n_322),
.Y(n_4238)
);

NOR2x1_ASAP7_75t_L g4239 ( 
.A(n_4158),
.B(n_323),
.Y(n_4239)
);

OR2x2_ASAP7_75t_L g4240 ( 
.A(n_4153),
.B(n_4122),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_4194),
.B(n_4168),
.Y(n_4241)
);

OAI21xp33_ASAP7_75t_L g4242 ( 
.A1(n_4184),
.A2(n_4183),
.B(n_4210),
.Y(n_4242)
);

AND2x2_ASAP7_75t_L g4243 ( 
.A(n_4192),
.B(n_4160),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_4205),
.B(n_4125),
.Y(n_4244)
);

NAND2x1_ASAP7_75t_L g4245 ( 
.A(n_4223),
.B(n_4141),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4199),
.B(n_4157),
.Y(n_4246)
);

O2A1O1Ixp33_ASAP7_75t_SL g4247 ( 
.A1(n_4196),
.A2(n_4135),
.B(n_4132),
.C(n_4171),
.Y(n_4247)
);

NOR3xp33_ASAP7_75t_L g4248 ( 
.A(n_4175),
.B(n_4156),
.C(n_4154),
.Y(n_4248)
);

OAI21xp5_ASAP7_75t_SL g4249 ( 
.A1(n_4198),
.A2(n_4167),
.B(n_4151),
.Y(n_4249)
);

XOR2x2_ASAP7_75t_L g4250 ( 
.A(n_4234),
.B(n_4167),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4191),
.B(n_324),
.Y(n_4251)
);

OR2x2_ASAP7_75t_L g4252 ( 
.A(n_4185),
.B(n_324),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_4206),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4217),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4206),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4186),
.Y(n_4256)
);

OAI322xp33_ASAP7_75t_L g4257 ( 
.A1(n_4187),
.A2(n_4216),
.A3(n_4202),
.B1(n_4201),
.B2(n_4230),
.C1(n_4181),
.C2(n_4182),
.Y(n_4257)
);

NAND2x1_ASAP7_75t_L g4258 ( 
.A(n_4223),
.B(n_4219),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4190),
.Y(n_4259)
);

NOR2xp33_ASAP7_75t_L g4260 ( 
.A(n_4197),
.B(n_325),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4220),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4209),
.B(n_326),
.Y(n_4262)
);

OAI321xp33_ASAP7_75t_L g4263 ( 
.A1(n_4176),
.A2(n_327),
.A3(n_328),
.B1(n_329),
.B2(n_330),
.C(n_331),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4238),
.Y(n_4264)
);

NAND2xp33_ASAP7_75t_SL g4265 ( 
.A(n_4229),
.B(n_332),
.Y(n_4265)
);

OAI22xp5_ASAP7_75t_L g4266 ( 
.A1(n_4193),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_4266)
);

AND2x2_ASAP7_75t_L g4267 ( 
.A(n_4212),
.B(n_4226),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4227),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_4240),
.Y(n_4269)
);

NOR2xp33_ASAP7_75t_L g4270 ( 
.A(n_4177),
.B(n_334),
.Y(n_4270)
);

INVx1_ASAP7_75t_SL g4271 ( 
.A(n_4239),
.Y(n_4271)
);

INVx1_ASAP7_75t_SL g4272 ( 
.A(n_4215),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4218),
.Y(n_4273)
);

OR2x2_ASAP7_75t_L g4274 ( 
.A(n_4221),
.B(n_335),
.Y(n_4274)
);

OAI211xp5_ASAP7_75t_L g4275 ( 
.A1(n_4177),
.A2(n_336),
.B(n_337),
.C(n_339),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4222),
.Y(n_4276)
);

A2O1A1Ixp33_ASAP7_75t_L g4277 ( 
.A1(n_4203),
.A2(n_340),
.B(n_341),
.C(n_342),
.Y(n_4277)
);

HB1xp67_ASAP7_75t_L g4278 ( 
.A(n_4203),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4211),
.B(n_341),
.Y(n_4279)
);

AOI222xp33_ASAP7_75t_L g4280 ( 
.A1(n_4188),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.C1(n_346),
.C2(n_347),
.Y(n_4280)
);

INVx1_ASAP7_75t_SL g4281 ( 
.A(n_4207),
.Y(n_4281)
);

INVxp67_ASAP7_75t_L g4282 ( 
.A(n_4208),
.Y(n_4282)
);

OAI21xp33_ASAP7_75t_L g4283 ( 
.A1(n_4179),
.A2(n_4200),
.B(n_4178),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4233),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_4214),
.B(n_345),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4180),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4189),
.Y(n_4287)
);

NOR2xp33_ASAP7_75t_L g4288 ( 
.A(n_4237),
.B(n_346),
.Y(n_4288)
);

OR2x2_ASAP7_75t_L g4289 ( 
.A(n_4232),
.B(n_347),
.Y(n_4289)
);

XOR2x2_ASAP7_75t_L g4290 ( 
.A(n_4195),
.B(n_348),
.Y(n_4290)
);

INVxp67_ASAP7_75t_L g4291 ( 
.A(n_4225),
.Y(n_4291)
);

OAI21xp5_ASAP7_75t_SL g4292 ( 
.A1(n_4213),
.A2(n_349),
.B(n_350),
.Y(n_4292)
);

HB1xp67_ASAP7_75t_L g4293 ( 
.A(n_4228),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4204),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4236),
.B(n_349),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_4278),
.B(n_4235),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_R g4297 ( 
.A(n_4265),
.B(n_4256),
.Y(n_4297)
);

NOR2xp33_ASAP7_75t_L g4298 ( 
.A(n_4257),
.B(n_4231),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4255),
.Y(n_4299)
);

NOR3xp33_ASAP7_75t_SL g4300 ( 
.A(n_4283),
.B(n_4224),
.C(n_352),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4271),
.B(n_4243),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4271),
.B(n_351),
.Y(n_4302)
);

AOI31xp33_ASAP7_75t_L g4303 ( 
.A1(n_4293),
.A2(n_351),
.A3(n_353),
.B(n_354),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4270),
.B(n_353),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4267),
.B(n_4264),
.Y(n_4305)
);

NOR3xp33_ASAP7_75t_SL g4306 ( 
.A(n_4242),
.B(n_355),
.C(n_356),
.Y(n_4306)
);

NOR2xp33_ASAP7_75t_L g4307 ( 
.A(n_4245),
.B(n_355),
.Y(n_4307)
);

XOR2xp5_ASAP7_75t_L g4308 ( 
.A(n_4250),
.B(n_359),
.Y(n_4308)
);

INVx1_ASAP7_75t_SL g4309 ( 
.A(n_4274),
.Y(n_4309)
);

NOR3xp33_ASAP7_75t_SL g4310 ( 
.A(n_4249),
.B(n_359),
.C(n_362),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4253),
.Y(n_4311)
);

OR2x2_ASAP7_75t_L g4312 ( 
.A(n_4258),
.B(n_362),
.Y(n_4312)
);

OR2x2_ASAP7_75t_L g4313 ( 
.A(n_4252),
.B(n_363),
.Y(n_4313)
);

BUFx4f_ASAP7_75t_SL g4314 ( 
.A(n_4272),
.Y(n_4314)
);

CKINVDCx16_ASAP7_75t_R g4315 ( 
.A(n_4272),
.Y(n_4315)
);

INVxp67_ASAP7_75t_L g4316 ( 
.A(n_4288),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4254),
.B(n_363),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4279),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4260),
.B(n_364),
.Y(n_4319)
);

AOI21xp33_ASAP7_75t_L g4320 ( 
.A1(n_4241),
.A2(n_364),
.B(n_366),
.Y(n_4320)
);

OR2x2_ASAP7_75t_L g4321 ( 
.A(n_4246),
.B(n_366),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4262),
.Y(n_4322)
);

AND3x2_ASAP7_75t_L g4323 ( 
.A(n_4269),
.B(n_367),
.C(n_368),
.Y(n_4323)
);

NOR2xp33_ASAP7_75t_R g4324 ( 
.A(n_4261),
.B(n_368),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4277),
.B(n_4280),
.Y(n_4325)
);

BUFx10_ASAP7_75t_L g4326 ( 
.A(n_4286),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4292),
.B(n_369),
.Y(n_4327)
);

NAND3xp33_ASAP7_75t_L g4328 ( 
.A(n_4275),
.B(n_370),
.C(n_371),
.Y(n_4328)
);

OAI21xp5_ASAP7_75t_SL g4329 ( 
.A1(n_4292),
.A2(n_4249),
.B(n_4281),
.Y(n_4329)
);

XNOR2xp5_ASAP7_75t_L g4330 ( 
.A(n_4290),
.B(n_370),
.Y(n_4330)
);

NOR3xp33_ASAP7_75t_L g4331 ( 
.A(n_4244),
.B(n_371),
.C(n_372),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4289),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4287),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_4281),
.B(n_372),
.Y(n_4334)
);

XOR2x2_ASAP7_75t_L g4335 ( 
.A(n_4248),
.B(n_373),
.Y(n_4335)
);

NOR2xp33_ASAP7_75t_L g4336 ( 
.A(n_4285),
.B(n_374),
.Y(n_4336)
);

NOR2xp67_ASAP7_75t_L g4337 ( 
.A(n_4328),
.B(n_4263),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4301),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4312),
.Y(n_4339)
);

INVxp67_ASAP7_75t_L g4340 ( 
.A(n_4307),
.Y(n_4340)
);

NOR2x1_ASAP7_75t_L g4341 ( 
.A(n_4329),
.B(n_4251),
.Y(n_4341)
);

OAI22xp5_ASAP7_75t_L g4342 ( 
.A1(n_4315),
.A2(n_4294),
.B1(n_4259),
.B2(n_4268),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4323),
.B(n_4273),
.Y(n_4343)
);

NOR3xp33_ASAP7_75t_L g4344 ( 
.A(n_4329),
.B(n_4282),
.C(n_4291),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_4334),
.B(n_4284),
.Y(n_4345)
);

AOI21xp5_ASAP7_75t_L g4346 ( 
.A1(n_4296),
.A2(n_4247),
.B(n_4263),
.Y(n_4346)
);

NOR3xp33_ASAP7_75t_L g4347 ( 
.A(n_4319),
.B(n_4276),
.C(n_4295),
.Y(n_4347)
);

XNOR2xp5_ASAP7_75t_L g4348 ( 
.A(n_4308),
.B(n_4266),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4314),
.Y(n_4349)
);

OAI21xp33_ASAP7_75t_L g4350 ( 
.A1(n_4298),
.A2(n_374),
.B(n_995),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4302),
.Y(n_4351)
);

OAI21xp33_ASAP7_75t_SL g4352 ( 
.A1(n_4299),
.A2(n_2880),
.B(n_1032),
.Y(n_4352)
);

AOI211xp5_ASAP7_75t_L g4353 ( 
.A1(n_4328),
.A2(n_1094),
.B(n_1032),
.C(n_1045),
.Y(n_4353)
);

AOI211x1_ASAP7_75t_L g4354 ( 
.A1(n_4311),
.A2(n_2880),
.B(n_1045),
.C(n_1051),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_4304),
.A2(n_1094),
.B(n_1051),
.Y(n_4355)
);

XNOR2x1_ASAP7_75t_SL g4356 ( 
.A(n_4330),
.B(n_1094),
.Y(n_4356)
);

AOI21xp5_ASAP7_75t_L g4357 ( 
.A1(n_4327),
.A2(n_1094),
.B(n_1051),
.Y(n_4357)
);

AOI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_4325),
.A2(n_1094),
.B(n_1051),
.Y(n_4358)
);

OAI211xp5_ASAP7_75t_L g4359 ( 
.A1(n_4297),
.A2(n_1094),
.B(n_1051),
.C(n_1083),
.Y(n_4359)
);

NAND3xp33_ASAP7_75t_L g4360 ( 
.A(n_4306),
.B(n_1076),
.C(n_1051),
.Y(n_4360)
);

OAI21xp33_ASAP7_75t_SL g4361 ( 
.A1(n_4305),
.A2(n_1076),
.B(n_1083),
.Y(n_4361)
);

OAI22xp33_ASAP7_75t_L g4362 ( 
.A1(n_4349),
.A2(n_4309),
.B1(n_4321),
.B2(n_4317),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4337),
.B(n_4310),
.Y(n_4363)
);

OR2x2_ASAP7_75t_L g4364 ( 
.A(n_4339),
.B(n_4313),
.Y(n_4364)
);

OA22x2_ASAP7_75t_L g4365 ( 
.A1(n_4348),
.A2(n_4318),
.B1(n_4322),
.B2(n_4332),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4338),
.B(n_4303),
.Y(n_4366)
);

INVxp67_ASAP7_75t_L g4367 ( 
.A(n_4341),
.Y(n_4367)
);

OAI21xp33_ASAP7_75t_SL g4368 ( 
.A1(n_4356),
.A2(n_4343),
.B(n_4345),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4342),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_4346),
.B(n_4331),
.Y(n_4370)
);

XNOR2xp5_ASAP7_75t_L g4371 ( 
.A(n_4344),
.B(n_4335),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4340),
.Y(n_4372)
);

OAI221xp5_ASAP7_75t_L g4373 ( 
.A1(n_4350),
.A2(n_4300),
.B1(n_4316),
.B2(n_4333),
.C(n_4347),
.Y(n_4373)
);

INVx2_ASAP7_75t_SL g4374 ( 
.A(n_4351),
.Y(n_4374)
);

NOR2xp33_ASAP7_75t_L g4375 ( 
.A(n_4359),
.B(n_4320),
.Y(n_4375)
);

OAI21xp33_ASAP7_75t_L g4376 ( 
.A1(n_4353),
.A2(n_4336),
.B(n_4324),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4353),
.Y(n_4377)
);

AOI221xp5_ASAP7_75t_L g4378 ( 
.A1(n_4367),
.A2(n_4358),
.B1(n_4354),
.B2(n_4361),
.C(n_4360),
.Y(n_4378)
);

AOI22xp5_ASAP7_75t_L g4379 ( 
.A1(n_4369),
.A2(n_4326),
.B1(n_4352),
.B2(n_4355),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4363),
.Y(n_4380)
);

AOI22xp5_ASAP7_75t_L g4381 ( 
.A1(n_4365),
.A2(n_4326),
.B1(n_4357),
.B2(n_1072),
.Y(n_4381)
);

AOI22xp5_ASAP7_75t_L g4382 ( 
.A1(n_4372),
.A2(n_1076),
.B1(n_1083),
.B2(n_1072),
.Y(n_4382)
);

AOI22xp5_ASAP7_75t_L g4383 ( 
.A1(n_4371),
.A2(n_1076),
.B1(n_1083),
.B2(n_1072),
.Y(n_4383)
);

NOR3xp33_ASAP7_75t_L g4384 ( 
.A(n_4373),
.B(n_1076),
.C(n_1083),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_4362),
.B(n_1083),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4364),
.Y(n_4386)
);

AO22x2_ASAP7_75t_L g4387 ( 
.A1(n_4374),
.A2(n_1072),
.B1(n_1075),
.B2(n_1076),
.Y(n_4387)
);

NOR4xp25_ASAP7_75t_L g4388 ( 
.A(n_4368),
.B(n_1075),
.C(n_1072),
.D(n_973),
.Y(n_4388)
);

OAI211xp5_ASAP7_75t_L g4389 ( 
.A1(n_4386),
.A2(n_4370),
.B(n_4376),
.C(n_4366),
.Y(n_4389)
);

XNOR2xp5_ASAP7_75t_L g4390 ( 
.A(n_4380),
.B(n_4377),
.Y(n_4390)
);

OAI22xp5_ASAP7_75t_L g4391 ( 
.A1(n_4379),
.A2(n_4375),
.B1(n_1075),
.B2(n_1072),
.Y(n_4391)
);

AOI22xp5_ASAP7_75t_L g4392 ( 
.A1(n_4384),
.A2(n_1075),
.B1(n_1304),
.B2(n_1296),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4378),
.B(n_1075),
.Y(n_4393)
);

AO22x2_ASAP7_75t_L g4394 ( 
.A1(n_4385),
.A2(n_1075),
.B1(n_1304),
.B2(n_1296),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4387),
.Y(n_4395)
);

AND2x4_ASAP7_75t_L g4396 ( 
.A(n_4395),
.B(n_4381),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4390),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4389),
.Y(n_4398)
);

XOR2xp5_ASAP7_75t_L g4399 ( 
.A(n_4391),
.B(n_4383),
.Y(n_4399)
);

OAI22xp33_ASAP7_75t_L g4400 ( 
.A1(n_4393),
.A2(n_4382),
.B1(n_4388),
.B2(n_1298),
.Y(n_4400)
);

NOR2x1_ASAP7_75t_L g4401 ( 
.A(n_4394),
.B(n_1296),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4398),
.B(n_4392),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4397),
.B(n_973),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4403),
.Y(n_4404)
);

INVx3_ASAP7_75t_L g4405 ( 
.A(n_4402),
.Y(n_4405)
);

OAI211xp5_ASAP7_75t_SL g4406 ( 
.A1(n_4405),
.A2(n_4400),
.B(n_4401),
.C(n_4396),
.Y(n_4406)
);

XNOR2x1_ASAP7_75t_L g4407 ( 
.A(n_4406),
.B(n_4405),
.Y(n_4407)
);

XOR2xp5_ASAP7_75t_L g4408 ( 
.A(n_4407),
.B(n_4399),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4408),
.B(n_4404),
.Y(n_4409)
);

CKINVDCx20_ASAP7_75t_R g4410 ( 
.A(n_4409),
.Y(n_4410)
);

NAND4xp75_ASAP7_75t_L g4411 ( 
.A(n_4410),
.B(n_1298),
.C(n_1304),
.D(n_1266),
.Y(n_4411)
);

OAI322xp33_ASAP7_75t_L g4412 ( 
.A1(n_4411),
.A2(n_1298),
.A3(n_1304),
.B1(n_1266),
.B2(n_973),
.C1(n_1347),
.C2(n_1494),
.Y(n_4412)
);

AOI22xp33_ASAP7_75t_L g4413 ( 
.A1(n_4412),
.A2(n_1298),
.B1(n_1304),
.B2(n_973),
.Y(n_4413)
);

AOI322xp5_ASAP7_75t_L g4414 ( 
.A1(n_4413),
.A2(n_1298),
.A3(n_973),
.B1(n_1347),
.B2(n_1494),
.C1(n_1053),
.C2(n_1197),
.Y(n_4414)
);

OR2x2_ASAP7_75t_L g4415 ( 
.A(n_4414),
.B(n_1053),
.Y(n_4415)
);

AOI21xp5_ASAP7_75t_L g4416 ( 
.A1(n_4415),
.A2(n_1053),
.B(n_1197),
.Y(n_4416)
);

AOI211xp5_ASAP7_75t_L g4417 ( 
.A1(n_4416),
.A2(n_1053),
.B(n_4398),
.C(n_4397),
.Y(n_4417)
);


endmodule