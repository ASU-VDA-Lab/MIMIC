module fake_jpeg_827_n_513 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_513);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_513;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_22),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_65),
.Y(n_117)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_53),
.Y(n_105)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_54),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_19),
.B(n_15),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_99),
.Y(n_113)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_95),
.Y(n_119)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_90),
.Y(n_140)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_15),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_39),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_101),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_55),
.A2(n_30),
.B1(n_48),
.B2(n_47),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_107),
.A2(n_154),
.B1(n_41),
.B2(n_24),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_49),
.B(n_45),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_114),
.B(n_34),
.Y(n_188)
);

FAx1_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_35),
.CI(n_39),
.CON(n_115),
.SN(n_115)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_115),
.A2(n_149),
.B(n_114),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_63),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_25),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_145),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_51),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_70),
.Y(n_131)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_88),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_54),
.B(n_47),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_58),
.A2(n_48),
.B1(n_30),
.B2(n_35),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_150),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_59),
.A2(n_48),
.B1(n_30),
.B2(n_36),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_36),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_100),
.Y(n_181)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_167),
.A2(n_196),
.B1(n_105),
.B2(n_155),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_115),
.A2(n_67),
.B1(n_102),
.B2(n_74),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_168),
.A2(n_175),
.B1(n_190),
.B2(n_203),
.Y(n_245)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_171),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_175)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_113),
.B(n_44),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_177),
.B(n_187),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_86),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_180),
.Y(n_234)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_183),
.Y(n_259)
);

OR2x6_ASAP7_75t_SL g246 ( 
.A(n_184),
.B(n_162),
.Y(n_246)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_34),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_193),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_149),
.A2(n_141),
.B1(n_128),
.B2(n_123),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_189),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_151),
.A2(n_83),
.B1(n_101),
.B2(n_48),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_191),
.Y(n_265)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_79),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_120),
.A2(n_82),
.B1(n_91),
.B2(n_90),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_109),
.Y(n_199)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_205),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_116),
.A2(n_89),
.B1(n_87),
.B2(n_41),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_106),
.B(n_38),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_204),
.B(n_215),
.Y(n_258)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_98),
.B1(n_35),
.B2(n_45),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_137),
.B(n_49),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_142),
.B(n_44),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_98),
.B1(n_35),
.B2(n_38),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_116),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_104),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_212),
.Y(n_250)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_26),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_217),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_141),
.B(n_35),
.Y(n_217)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_136),
.Y(n_238)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_133),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_122),
.B(n_15),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_109),
.C(n_155),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_175),
.A2(n_124),
.B1(n_26),
.B2(n_111),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_222),
.A2(n_231),
.B1(n_244),
.B2(n_252),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_225),
.A2(n_132),
.B1(n_189),
.B2(n_185),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_188),
.A2(n_111),
.B1(n_140),
.B2(n_122),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_232),
.B(n_2),
.Y(n_300)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_163),
.B(n_129),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_266),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_190),
.A2(n_211),
.B1(n_203),
.B2(n_206),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_194),
.B(n_183),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_196),
.A2(n_136),
.B1(n_120),
.B2(n_138),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_225),
.B1(n_245),
.B2(n_238),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_143),
.B1(n_138),
.B2(n_133),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_217),
.B(n_132),
.CI(n_158),
.CON(n_263),
.SN(n_263)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_199),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_166),
.B(n_143),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_221),
.B(n_179),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_269),
.B(n_283),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_272),
.A2(n_280),
.B1(n_287),
.B2(n_304),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_172),
.B1(n_219),
.B2(n_212),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_306),
.B1(n_307),
.B2(n_254),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_275),
.A2(n_298),
.B1(n_302),
.B2(n_224),
.Y(n_320)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_279),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_223),
.B1(n_228),
.B2(n_250),
.Y(n_280)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

AND2x6_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_164),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_294),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_237),
.B(n_201),
.Y(n_283)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_218),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_290),
.Y(n_315)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_243),
.B(n_198),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_288),
.B(n_291),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_295),
.B(n_270),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_173),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_165),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_228),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_293),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_202),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_191),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_133),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_301),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_1),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_303),
.Y(n_338)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_224),
.Y(n_297)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_246),
.A2(n_183),
.B1(n_192),
.B2(n_4),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_242),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_232),
.B(n_2),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_229),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_3),
.Y(n_303)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_5),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_308),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_248),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_265),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_227),
.B(n_7),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_230),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_251),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_292),
.A2(n_263),
.B1(n_240),
.B2(n_236),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_310),
.A2(n_336),
.B1(n_342),
.B2(n_306),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_249),
.C(n_262),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_316),
.C(n_322),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_312),
.A2(n_319),
.B(n_293),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_230),
.C(n_239),
.Y(n_316)
);

AO22x1_ASAP7_75t_L g318 ( 
.A1(n_298),
.A2(n_263),
.B1(n_265),
.B2(n_224),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_318),
.A2(n_302),
.B(n_273),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_289),
.A2(n_264),
.B(n_260),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_320),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_272),
.A2(n_236),
.B1(n_264),
.B2(n_260),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_321),
.A2(n_327),
.B1(n_337),
.B2(n_279),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_235),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_335),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_235),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_330),
.C(n_295),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_274),
.A2(n_265),
.B1(n_239),
.B2(n_242),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

MAJx2_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_251),
.C(n_254),
.Y(n_330)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_270),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_271),
.A2(n_261),
.B1(n_259),
.B2(n_10),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_274),
.A2(n_259),
.B1(n_9),
.B2(n_10),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_271),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_332),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_351),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_333),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_339),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_286),
.C(n_277),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_357),
.C(n_362),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_268),
.B(n_282),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_355),
.A2(n_358),
.B(n_365),
.Y(n_386)
);

BUFx2_ASAP7_75t_SL g356 ( 
.A(n_325),
.Y(n_356)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_293),
.C(n_278),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_366),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_311),
.C(n_326),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_309),
.C(n_285),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_371),
.C(n_376),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_283),
.B(n_297),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_315),
.Y(n_367)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_367),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_287),
.Y(n_368)
);

AO21x1_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_341),
.B(n_340),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_276),
.B1(n_304),
.B2(n_299),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_369),
.A2(n_373),
.B1(n_320),
.B2(n_361),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_281),
.C(n_299),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_338),
.B(n_11),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_372),
.B(n_374),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_310),
.A2(n_279),
.B1(n_12),
.B2(n_13),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_279),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_375),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_340),
.C(n_330),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_344),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_377),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_378),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_379),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_340),
.C(n_346),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_348),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_387),
.B(n_389),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_354),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_334),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_393),
.C(n_398),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_359),
.A2(n_321),
.B1(n_314),
.B2(n_327),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_392),
.A2(n_360),
.B1(n_363),
.B2(n_351),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_334),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_317),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_350),
.B(n_317),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_401),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_379),
.A2(n_318),
.B1(n_314),
.B2(n_337),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_403),
.A2(n_405),
.B1(n_378),
.B2(n_360),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_318),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_407),
.C(n_357),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_379),
.A2(n_344),
.B1(n_343),
.B2(n_14),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_343),
.C(n_12),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_411),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_410),
.A2(n_415),
.B1(n_420),
.B2(n_421),
.Y(n_445)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_397),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_402),
.B(n_366),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_428),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_395),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_352),
.C(n_376),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_395),
.C(n_390),
.Y(n_449)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_397),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_388),
.B(n_370),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_417),
.B(n_425),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_380),
.A2(n_360),
.B1(n_347),
.B2(n_355),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_396),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_422),
.A2(n_424),
.B1(n_426),
.B2(n_403),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_386),
.A2(n_385),
.B(n_381),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_423),
.A2(n_433),
.B(n_400),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_386),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_399),
.B(n_375),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_408),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_404),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_394),
.B(n_364),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_431),
.A2(n_432),
.B1(n_400),
.B2(n_377),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_381),
.A2(n_363),
.B1(n_358),
.B2(n_365),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_385),
.A2(n_373),
.B(n_368),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_424),
.A2(n_394),
.B(n_402),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_434),
.B(n_448),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_435),
.Y(n_463)
);

MAJx2_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_384),
.C(n_387),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_438),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_382),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_442),
.Y(n_455)
);

XNOR2x2_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_406),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_439),
.A2(n_433),
.B(n_418),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_389),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_453),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_451),
.C(n_452),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_390),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_406),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_399),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_407),
.C(n_383),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_430),
.C(n_449),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_461),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_435),
.A2(n_423),
.B(n_416),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_458),
.A2(n_425),
.B(n_392),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_459),
.A2(n_452),
.B(n_445),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_412),
.C(n_422),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_464),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_444),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_467),
.Y(n_480)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_466),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_409),
.C(n_410),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_442),
.C(n_437),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_472),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_471),
.A2(n_481),
.B(n_483),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_456),
.B(n_453),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_463),
.A2(n_415),
.B1(n_451),
.B2(n_426),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_468),
.B1(n_11),
.B2(n_14),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_446),
.Y(n_477)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_477),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_436),
.Y(n_478)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_478),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_482),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_457),
.A2(n_421),
.B(n_440),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_463),
.A2(n_431),
.B1(n_405),
.B2(n_369),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_458),
.A2(n_459),
.B(n_461),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_457),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_486),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_460),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_455),
.C(n_460),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_490),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_455),
.C(n_468),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_494),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_482),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_11),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_475),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_500),
.Y(n_502)
);

AOI21xp33_ASAP7_75t_L g498 ( 
.A1(n_485),
.A2(n_478),
.B(n_471),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_501),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_473),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_490),
.C(n_499),
.Y(n_504)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_504),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_492),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_505),
.B(n_491),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_506),
.A2(n_504),
.B1(n_503),
.B2(n_502),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_507),
.Y(n_509)
);

MAJx2_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_500),
.C(n_488),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_510),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_511),
.B(n_488),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_493),
.Y(n_513)
);


endmodule