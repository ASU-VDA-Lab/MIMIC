module fake_jpeg_16335_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx10_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_19),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_25),
.B1(n_18),
.B2(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_15),
.B(n_0),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_60),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_27),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_27),
.B(n_23),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_19),
.B1(n_24),
.B2(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_58),
.B1(n_16),
.B2(n_20),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_53),
.B1(n_30),
.B2(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_39),
.B1(n_42),
.B2(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_25),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_42),
.B(n_30),
.C(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_18),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_22),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_72),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_17),
.B1(n_21),
.B2(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_42),
.B1(n_38),
.B2(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_80),
.B1(n_64),
.B2(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_31),
.B1(n_21),
.B2(n_17),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_77),
.B(n_60),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_57),
.B1(n_20),
.B2(n_22),
.Y(n_108)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_37),
.B1(n_34),
.B2(n_29),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_74),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_49),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_97),
.B(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_104),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_44),
.B1(n_43),
.B2(n_21),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_103),
.B1(n_111),
.B2(n_91),
.Y(n_115)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_107),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_55),
.B(n_62),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_55),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_65),
.C(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_61),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_77),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_34),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_57),
.B1(n_22),
.B2(n_20),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_113),
.B(n_121),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_129),
.B1(n_72),
.B2(n_85),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_80),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_103),
.C(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_86),
.B1(n_84),
.B2(n_69),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_89),
.B1(n_108),
.B2(n_101),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_88),
.B1(n_37),
.B2(n_71),
.Y(n_150)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_67),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_134),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_46),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_137),
.C(n_112),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_97),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_150),
.B1(n_154),
.B2(n_131),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_90),
.C(n_101),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_132),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_107),
.B(n_90),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_152),
.B(n_144),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_128),
.B1(n_133),
.B2(n_123),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_96),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_123),
.Y(n_172)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_155),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_46),
.B1(n_109),
.B2(n_36),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_163),
.C(n_164),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_170),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_162),
.B1(n_175),
.B2(n_127),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_128),
.B1(n_115),
.B2(n_112),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_125),
.C(n_124),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_125),
.C(n_117),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_10),
.B(n_14),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_148),
.C(n_141),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_174),
.C(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

XNOR2x2_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_156),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_120),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_119),
.B1(n_127),
.B2(n_46),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_127),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_150),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_50),
.C(n_29),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_136),
.B1(n_154),
.B2(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_181),
.B1(n_186),
.B2(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_163),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_151),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_165),
.B1(n_176),
.B2(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_172),
.C(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_203),
.Y(n_214)
);

AOI22x1_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_158),
.B1(n_174),
.B2(n_164),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_198),
.A2(n_184),
.B1(n_186),
.B2(n_189),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_50),
.C(n_36),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_50),
.C(n_23),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_50),
.C(n_23),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_23),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_178),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_28),
.B(n_1),
.C(n_2),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_207),
.B1(n_190),
.B2(n_4),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_180),
.B(n_177),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_207),
.B(n_9),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_200),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_184),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_207),
.C(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_199),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_202),
.B1(n_203),
.B2(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_206),
.B(n_179),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_212),
.C(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_225),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_223),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_29),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_232),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_213),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_214),
.A3(n_226),
.B1(n_218),
.B2(n_215),
.C1(n_6),
.C2(n_7),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_237),
.Y(n_242)
);

NAND2x1_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_218),
.Y(n_237)
);

AOI31xp33_ASAP7_75t_SL g238 ( 
.A1(n_229),
.A2(n_9),
.A3(n_13),
.B(n_12),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_239),
.B(n_231),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_29),
.A3(n_28),
.B1(n_36),
.B2(n_5),
.C1(n_6),
.C2(n_8),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_243),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_234),
.B(n_5),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_2),
.B(n_3),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_5),
.B(n_12),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_3),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_23),
.C(n_4),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_4),
.Y(n_250)
);


endmodule