module real_jpeg_25805_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_72),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_69),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_69),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_6),
.A2(n_26),
.B1(n_103),
.B2(n_108),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_6),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_6),
.A2(n_26),
.B1(n_51),
.B2(n_52),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_8),
.B(n_51),
.C(n_63),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_116),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_8),
.A2(n_56),
.B1(n_85),
.B2(n_156),
.Y(n_155)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_58),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_13),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_20),
.B(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.C(n_74),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_21),
.A2(n_22),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_42),
.C(n_59),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_32),
.B2(n_38),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_25),
.A2(n_31),
.B1(n_77),
.B2(n_116),
.Y(n_178)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

HAxp5_ASAP7_75t_SL g77 ( 
.A(n_27),
.B(n_78),
.CON(n_77),
.SN(n_77)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_34),
.C(n_36),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_27),
.A2(n_46),
.B(n_92),
.C(n_95),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_47),
.C(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_31),
.A2(n_39),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_33),
.A2(n_35),
.B(n_77),
.C(n_79),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_35),
.B(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_59),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_102),
.B1(n_106),
.B2(n_111),
.Y(n_101)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_107),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_46),
.A2(n_47),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_53),
.B(n_55),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_49),
.Y(n_97)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_54),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_52),
.B1(n_63),
.B2(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_52),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_53),
.A2(n_83),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_54),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_85),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_56),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_56),
.A2(n_149),
.B1(n_156),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_60),
.A2(n_74),
.B1(n_75),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_60),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_67),
.B(n_70),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_61),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_61),
.A2(n_66),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_61),
.A2(n_66),
.B1(n_134),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_66),
.B(n_78),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_68),
.A2(n_73),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_76),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_93),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_92),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_78),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_82),
.B(n_86),
.Y(n_144)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_100),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_113),
.Y(n_100)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_181),
.B(n_187),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_170),
.B(n_180),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_145),
.B(n_169),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_131),
.B1(n_132),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_153),
.B(n_168),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_151),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_162),
.B(n_167),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_164),
.Y(n_167)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_179),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_175),
.C(n_178),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_182),
.B(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);


endmodule