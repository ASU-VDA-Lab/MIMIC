module fake_netlist_1_6772_n_28 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_10), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
AO31x2_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_15), .A3(n_12), .B(n_11), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_17), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_16), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
OAI21xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_16), .B(n_1), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
NAND5xp2_ASAP7_75t_L g25 ( .A(n_23), .B(n_0), .C(n_3), .D(n_4), .E(n_7), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
XNOR2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_24), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
endmodule