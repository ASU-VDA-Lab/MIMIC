module fake_jpeg_9616_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_12),
.B1(n_17),
.B2(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

A2O1A1O1Ixp25_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_25),
.B(n_19),
.C(n_21),
.D(n_10),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_45),
.C(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_15),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_17),
.B1(n_36),
.B2(n_11),
.Y(n_52)
);

AO22x2_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_36),
.B1(n_37),
.B2(n_31),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

XNOR2x2_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_41),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_43),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_58),
.B(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_42),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_40),
.B(n_45),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_20),
.C(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_62),
.B1(n_39),
.B2(n_20),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_55),
.C(n_34),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_68),
.C(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_57),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_14),
.Y(n_74)
);

AO221x1_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_59),
.C(n_7),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_14),
.B1(n_8),
.B2(n_9),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_65),
.C(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_9),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_76),
.B(n_6),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_8),
.Y(n_79)
);


endmodule