module real_jpeg_33774_n_4 (n_3, n_1, n_0, n_2, n_4);

input n_3;
input n_1;
input n_0;
input n_2;

output n_4;

wire n_5;
wire n_8;
wire n_12;
wire n_10;
wire n_15;
wire n_11;
wire n_14;
wire n_6;
wire n_7;
wire n_13;
wire n_9;

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_13),
.Y(n_14)
);

BUFx2_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_L g4 ( 
.A1(n_5),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_4)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g5 ( 
.A1(n_6),
.A2(n_7),
.B(n_8),
.Y(n_5)
);

NAND2xp33_ASAP7_75t_SL g8 ( 
.A(n_6),
.B(n_7),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

AO21x1_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_13),
.B(n_14),
.Y(n_10)
);

INVx2_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);


endmodule