module fake_jpeg_10068_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_67),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_35),
.B1(n_34),
.B2(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_22),
.B1(n_21),
.B2(n_43),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_35),
.B1(n_34),
.B2(n_25),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_84),
.B1(n_31),
.B2(n_30),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_42),
.B1(n_34),
.B2(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_88),
.B1(n_94),
.B2(n_69),
.Y(n_102)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_85),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_22),
.B(n_21),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_26),
.B(n_27),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_34),
.B1(n_21),
.B2(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_28),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_28),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_93),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_29),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_38),
.B1(n_40),
.B2(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_16),
.C(n_11),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_115),
.C(n_7),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_104),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_102),
.B1(n_87),
.B2(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_45),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_113),
.B1(n_87),
.B2(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_54),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_93),
.C(n_71),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_77),
.C(n_78),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_38),
.B(n_13),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_124),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_54),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_82),
.Y(n_142)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_126),
.B(n_15),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_75),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_127),
.A2(n_32),
.B(n_33),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_128),
.A2(n_129),
.B1(n_138),
.B2(n_143),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_75),
.B1(n_58),
.B2(n_76),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_97),
.C(n_55),
.Y(n_169)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_121),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_80),
.B1(n_73),
.B2(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_153),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_92),
.B1(n_95),
.B2(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_54),
.B1(n_50),
.B2(n_47),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_82),
.B1(n_72),
.B2(n_47),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_50),
.B1(n_78),
.B2(n_61),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_64),
.B1(n_45),
.B2(n_30),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_45),
.B1(n_31),
.B2(n_26),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_113),
.B(n_106),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_159),
.B(n_163),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_122),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_169),
.C(n_170),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_106),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_165),
.B(n_171),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_104),
.B1(n_119),
.B2(n_121),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_98),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

XOR2x2_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_97),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_167),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_105),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_18),
.Y(n_170)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_18),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_176),
.B1(n_178),
.B2(n_181),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_17),
.B(n_30),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_183),
.B(n_27),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_142),
.A2(n_149),
.B(n_131),
.C(n_150),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_125),
.C(n_118),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_152),
.C(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_203),
.C(n_210),
.Y(n_215)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_118),
.B1(n_125),
.B2(n_135),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_192),
.B1(n_202),
.B2(n_209),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_135),
.B1(n_27),
.B2(n_31),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_201),
.B(n_161),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_32),
.B(n_28),
.C(n_12),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_197),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_204),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_32),
.B(n_17),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_155),
.A2(n_168),
.B1(n_172),
.B2(n_166),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_165),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_133),
.B1(n_152),
.B2(n_19),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_211),
.B1(n_24),
.B2(n_23),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_155),
.A2(n_19),
.B1(n_133),
.B2(n_24),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_32),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_159),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_186),
.B(n_154),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_217),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_216),
.C(n_219),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_157),
.C(n_162),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_183),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_218),
.B(n_9),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_173),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_229),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_157),
.B(n_179),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_228),
.B(n_222),
.Y(n_247)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_175),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_227),
.C(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_180),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_181),
.C(n_161),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_193),
.B1(n_231),
.B2(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_193),
.B(n_207),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_252),
.B(n_256),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_213),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_255),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_207),
.B(n_189),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_190),
.B1(n_189),
.B2(n_196),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_217),
.A2(n_194),
.B(n_196),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_201),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_192),
.B1(n_200),
.B2(n_24),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_200),
.B1(n_19),
.B2(n_9),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_8),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_215),
.C(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_275),
.C(n_249),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_243),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_227),
.B1(n_214),
.B2(n_215),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_246),
.B1(n_258),
.B2(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_8),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_32),
.C(n_9),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_274),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_277),
.Y(n_289)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_252),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_17),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_17),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_7),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_17),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_248),
.B1(n_251),
.B2(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_247),
.B(n_244),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_282),
.A2(n_288),
.B(n_14),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_292),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_244),
.B1(n_251),
.B2(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_264),
.B(n_279),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_269),
.B(n_256),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_295),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_257),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_293),
.C(n_294),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_255),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_242),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_276),
.C(n_275),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_306),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_243),
.B1(n_267),
.B2(n_272),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_0),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_14),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_268),
.B(n_7),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_305),
.B(n_0),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_295),
.C(n_293),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_17),
.C(n_2),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_286),
.C(n_292),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_287),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_14),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_314),
.C(n_316),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_286),
.B(n_10),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_2),
.B(n_3),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_313),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_17),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_299),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_298),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_12),
.C(n_11),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_317),
.A2(n_318),
.B(n_2),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_296),
.B(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_321),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_298),
.B(n_3),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_4),
.B(n_5),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_2),
.B(n_4),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_328),
.B(n_329),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_327),
.C(n_330),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_322),
.B(n_320),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_4),
.B(n_5),
.Y(n_334)
);

OAI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_321),
.C(n_317),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_6),
.Y(n_336)
);


endmodule