module fake_jpeg_24218_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_30),
.B1(n_36),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_34),
.B1(n_26),
.B2(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NOR4xp25_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_18),
.C(n_26),
.D(n_2),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_19),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_31),
.B1(n_25),
.B2(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_66),
.B1(n_30),
.B2(n_23),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_43),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_42),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_74),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_78),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_30),
.B1(n_25),
.B2(n_36),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_57),
.B1(n_66),
.B2(n_52),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_93),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_26),
.B1(n_18),
.B2(n_43),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_90),
.B1(n_81),
.B2(n_88),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_23),
.B1(n_39),
.B2(n_44),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_92),
.B1(n_94),
.B2(n_21),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_26),
.B1(n_43),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_57),
.B1(n_53),
.B2(n_62),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_61),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_100),
.Y(n_103)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_0),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_108),
.B1(n_110),
.B2(n_123),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_57),
.B1(n_52),
.B2(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_124),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_52),
.B1(n_70),
.B2(n_49),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_100),
.B1(n_73),
.B2(n_82),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_70),
.B1(n_49),
.B2(n_62),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_95),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_62),
.B1(n_53),
.B2(n_49),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_56),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_73),
.A2(n_53),
.B1(n_55),
.B2(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_72),
.B(n_41),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_37),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_73),
.A2(n_55),
.B1(n_69),
.B2(n_48),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_90),
.B1(n_88),
.B2(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_133),
.B(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_146),
.B1(n_151),
.B2(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_141),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_88),
.B1(n_100),
.B2(n_77),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_148),
.B1(n_152),
.B2(n_158),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_77),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_161),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_100),
.B1(n_101),
.B2(n_99),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_86),
.C(n_55),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_123),
.C(n_124),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_96),
.B1(n_71),
.B2(n_89),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_86),
.B1(n_89),
.B2(n_45),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_89),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_157),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_41),
.B(n_45),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_136),
.B(n_137),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_48),
.B1(n_37),
.B2(n_32),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_109),
.B(n_29),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_103),
.A2(n_32),
.B1(n_20),
.B2(n_85),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_106),
.A2(n_32),
.B1(n_20),
.B2(n_85),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_160),
.B1(n_117),
.B2(n_118),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_20),
.B1(n_74),
.B2(n_29),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_114),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_177),
.C(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_169),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_168),
.A2(n_170),
.B(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_119),
.C(n_111),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_173),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_127),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_181),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_117),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_176),
.B(n_186),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_114),
.C(n_113),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_129),
.B1(n_113),
.B2(n_115),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_180),
.B1(n_160),
.B2(n_156),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_115),
.B1(n_102),
.B2(n_105),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_126),
.C(n_116),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_116),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_74),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_126),
.C(n_116),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_158),
.C(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_126),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_191),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_198),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_132),
.B(n_157),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_196),
.A2(n_214),
.B(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_178),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_162),
.A2(n_140),
.B1(n_146),
.B2(n_135),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_206),
.B1(n_211),
.B2(n_217),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_207),
.C(n_212),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_162),
.A2(n_140),
.B1(n_146),
.B2(n_148),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_132),
.C(n_140),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_156),
.B1(n_149),
.B2(n_160),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_149),
.C(n_139),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_29),
.B(n_1),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_216),
.B(n_220),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_104),
.B1(n_2),
.B2(n_3),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_183),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_164),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_166),
.A2(n_185),
.B(n_165),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_174),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_104),
.C(n_29),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_188),
.C(n_182),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_104),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_169),
.B1(n_15),
.B2(n_14),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_181),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_232),
.B1(n_244),
.B2(n_209),
.Y(n_254)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_235),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_173),
.B1(n_172),
.B2(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_164),
.Y(n_233)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_238),
.C(n_207),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_166),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_182),
.C(n_171),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_214),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_176),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_171),
.B1(n_167),
.B2(n_193),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_211),
.B1(n_206),
.B2(n_201),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_235),
.B1(n_239),
.B2(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_15),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_14),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_221),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_14),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_248),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_210),
.B(n_195),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_200),
.B(n_214),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_251),
.A2(n_262),
.B1(n_242),
.B2(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_265),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_242),
.A2(n_240),
.B1(n_250),
.B2(n_234),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_230),
.B1(n_194),
.B2(n_247),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_195),
.B(n_210),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_266),
.B(n_224),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_264),
.C(n_236),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_208),
.B1(n_200),
.B2(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_212),
.C(n_219),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_196),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_0),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g272 ( 
.A(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_238),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_279),
.C(n_282),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_255),
.B(n_3),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_267),
.B1(n_261),
.B2(n_268),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_225),
.C(n_246),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_262),
.B1(n_251),
.B2(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_220),
.C(n_218),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_227),
.C(n_243),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_287),
.C(n_288),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_258),
.C(n_252),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_0),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_268),
.Y(n_293)
);

OAI321xp33_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_266),
.A3(n_263),
.B1(n_260),
.B2(n_267),
.C(n_257),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_297),
.B(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_8),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_304),
.B1(n_297),
.B2(n_305),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_0),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_299),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_282),
.A2(n_4),
.B(n_5),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_4),
.C(n_5),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_302),
.A2(n_279),
.B(n_8),
.Y(n_311)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_6),
.B(n_7),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_289),
.B1(n_274),
.B2(n_9),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_277),
.A2(n_6),
.B(n_7),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_302),
.B(n_287),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_296),
.C(n_10),
.Y(n_322)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_314),
.C(n_9),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_273),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_281),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_315),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_303),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_9),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_298),
.C(n_295),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_316),
.B(n_318),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_322),
.B(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_326),
.B(n_10),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_335),
.C(n_327),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_333),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_310),
.B(n_317),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_332),
.A2(n_334),
.B(n_323),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_307),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_314),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_338),
.C(n_11),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_330),
.A2(n_328),
.B(n_324),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_10),
.B(n_11),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_341),
.B(n_336),
.C(n_12),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_12),
.C(n_13),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_13),
.Y(n_344)
);


endmodule