module fake_netlist_1_811_n_682 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_682);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_682;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_606;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_18), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_12), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_33), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_65), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_10), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_61), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_47), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_59), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_1), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_2), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_27), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_5), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_34), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_23), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_60), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_6), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_73), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_6), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_64), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_43), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_37), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_42), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_16), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_15), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_0), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_31), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_57), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_52), .Y(n_106) );
OR2x2_ASAP7_75t_L g107 ( .A(n_1), .B(n_22), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_45), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_49), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_50), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_25), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_4), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_38), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_30), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_44), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_46), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_48), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_63), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_20), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_74), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_88), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_90), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_116), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_92), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
NAND2xp33_ASAP7_75t_SL g132 ( .A(n_78), .B(n_0), .Y(n_132) );
CKINVDCx8_ASAP7_75t_R g133 ( .A(n_76), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_85), .B(n_2), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_97), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_110), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_106), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_94), .B(n_3), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_111), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_112), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_113), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_107), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_114), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_115), .Y(n_158) );
BUFx8_ASAP7_75t_L g159 ( .A(n_117), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_76), .B(n_3), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
INVxp67_ASAP7_75t_SL g164 ( .A(n_150), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_150), .B(n_121), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_150), .B(n_109), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_156), .B(n_83), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_123), .B(n_83), .Y(n_170) );
OAI221xp5_ASAP7_75t_L g171 ( .A1(n_154), .A2(n_98), .B1(n_104), .B2(n_93), .C(n_81), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_136), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
BUFx12f_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_127), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_123), .B(n_100), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_156), .B(n_91), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_161), .Y(n_183) );
BUFx8_ASAP7_75t_L g184 ( .A(n_161), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_124), .B(n_100), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_130), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_126), .B(n_91), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_127), .Y(n_189) );
AOI22x1_ASAP7_75t_L g190 ( .A1(n_130), .A2(n_89), .B1(n_108), .B2(n_101), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_134), .A2(n_122), .B(n_108), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_149), .B(n_122), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_141), .B(n_110), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_157), .B(n_80), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_158), .B(n_80), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_134), .B(n_36), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_137), .B(n_4), .Y(n_200) );
INVxp67_ASAP7_75t_SL g201 ( .A(n_140), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_137), .B(n_39), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_143), .B(n_35), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_125), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_143), .B(n_5), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_160), .B(n_40), .Y(n_206) );
AO221x1_ASAP7_75t_L g207 ( .A1(n_162), .A2(n_7), .B1(n_8), .B2(n_9), .C(n_10), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_125), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_160), .B(n_7), .Y(n_209) );
INVx8_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_139), .B(n_53), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_145), .B(n_8), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_139), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_142), .B(n_54), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_162), .B(n_9), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_133), .B(n_55), .Y(n_217) );
NOR2xp33_ASAP7_75t_R g218 ( .A(n_133), .B(n_51), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_131), .B(n_11), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_146), .B(n_11), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_131), .B(n_17), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_142), .B(n_19), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_181), .B(n_159), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_210), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_183), .A2(n_132), .B1(n_159), .B2(n_151), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_166), .B(n_163), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_169), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_183), .B(n_163), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_164), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_187), .B(n_155), .Y(n_232) );
BUFx8_ASAP7_75t_SL g233 ( .A(n_175), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_210), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_182), .A2(n_155), .B(n_152), .C(n_135), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_166), .B(n_152), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_199), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_165), .A2(n_132), .B1(n_135), .B2(n_142), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_167), .B(n_129), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_174), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_201), .B(n_148), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_172), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_199), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_166), .B(n_128), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_194), .B(n_148), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_188), .B(n_128), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_176), .A2(n_148), .B(n_147), .Y(n_247) );
NAND2xp33_ASAP7_75t_SL g248 ( .A(n_218), .B(n_148), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_186), .B(n_148), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_179), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_195), .Y(n_251) );
BUFx8_ASAP7_75t_L g252 ( .A(n_175), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_210), .B(n_147), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_196), .B(n_128), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_197), .B(n_147), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_212), .B(n_147), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_204), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_210), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_208), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_199), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_165), .B(n_147), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_171), .A2(n_21), .B(n_24), .C(n_26), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_185), .B(n_28), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_191), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_193), .B(n_29), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_191), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_195), .A2(n_32), .B1(n_56), .B2(n_58), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_165), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_165), .A2(n_62), .B1(n_66), .B2(n_68), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_165), .A2(n_69), .B1(n_70), .B2(n_72), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_216), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_220), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_200), .Y(n_274) );
INVx4_ASAP7_75t_L g275 ( .A(n_165), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_184), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_209), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_192), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_170), .B(n_75), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_170), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_192), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_178), .B(n_190), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_178), .B(n_206), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_184), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_198), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_213), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_214), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_213), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_257), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_274), .B(n_184), .Y(n_291) );
BUFx5_ASAP7_75t_L g292 ( .A(n_242), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_278), .B(n_222), .Y(n_293) );
INVx3_ASAP7_75t_SL g294 ( .A(n_252), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_231), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_230), .Y(n_296) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_247), .A2(n_203), .B(n_202), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_230), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_229), .B(n_221), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_252), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_240), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_234), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_251), .B(n_207), .Y(n_303) );
NOR2x1p5_ASAP7_75t_SL g304 ( .A(n_286), .B(n_168), .Y(n_304) );
OA21x2_ASAP7_75t_L g305 ( .A1(n_247), .A2(n_203), .B(n_202), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_285), .B(n_218), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_226), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_277), .B(n_219), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_272), .B(n_217), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_244), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_234), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_253), .A2(n_223), .B1(n_224), .B2(n_215), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_262), .A2(n_224), .B(n_215), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_226), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_226), .B(n_211), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g316 ( .A1(n_225), .A2(n_211), .B(n_173), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_232), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g318 ( .A1(n_225), .A2(n_168), .B1(n_173), .B2(n_177), .Y(n_318) );
CKINVDCx16_ASAP7_75t_R g319 ( .A(n_233), .Y(n_319) );
BUFx12f_ASAP7_75t_L g320 ( .A(n_244), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_273), .B(n_189), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_275), .B(n_177), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_238), .A2(n_180), .B1(n_189), .B2(n_275), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_234), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_226), .Y(n_325) );
CKINVDCx11_ASAP7_75t_R g326 ( .A(n_268), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_257), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_255), .B(n_180), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_239), .B(n_281), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_232), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_284), .A2(n_283), .B(n_241), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_284), .A2(n_283), .B(n_241), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_258), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_254), .A2(n_245), .B(n_228), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_250), .B(n_260), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_246), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_256), .B(n_236), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_259), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_317), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_330), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_335), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_335), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_293), .B(n_276), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_333), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_321), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_292), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_293), .B(n_276), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_328), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_291), .B(n_227), .Y(n_352) );
OA21x2_ASAP7_75t_L g353 ( .A1(n_316), .A2(n_313), .B(n_332), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_331), .A2(n_268), .B(n_280), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_291), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_331), .A2(n_280), .B(n_262), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_336), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_296), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_332), .A2(n_271), .B(n_270), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_299), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_292), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_292), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_292), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_290), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_327), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_342), .B(n_303), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_346), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_342), .B(n_329), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_343), .B(n_329), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_348), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_343), .B(n_326), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_356), .B(n_310), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_339), .B(n_309), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_364), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_341), .B(n_309), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_344), .B(n_276), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_350), .B(n_307), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_352), .A2(n_264), .B1(n_314), .B2(n_307), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_345), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_363), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_350), .B(n_314), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_340), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_351), .B(n_337), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_381), .Y(n_396) );
OR2x6_ASAP7_75t_L g397 ( .A(n_371), .B(n_364), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_381), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
INVx5_ASAP7_75t_L g400 ( .A(n_382), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_384), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_372), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_387), .B(n_367), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_384), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_352), .B1(n_361), .B2(n_264), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_390), .Y(n_408) );
AOI222xp33_ASAP7_75t_L g409 ( .A1(n_376), .A2(n_294), .B1(n_359), .B2(n_368), .C1(n_358), .C2(n_300), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_387), .B(n_367), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_389), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_392), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_378), .B(n_366), .Y(n_414) );
OA21x2_ASAP7_75t_L g415 ( .A1(n_378), .A2(n_360), .B(n_357), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_389), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_382), .Y(n_417) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_374), .A2(n_319), .A3(n_306), .B(n_325), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_374), .A2(n_365), .B1(n_349), .B2(n_362), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
INVx4_ASAP7_75t_SL g421 ( .A(n_390), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_395), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_369), .B(n_355), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_380), .B(n_355), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_369), .A2(n_355), .B1(n_349), .B2(n_362), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_392), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
BUFx2_ASAP7_75t_SL g429 ( .A(n_390), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_370), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_413), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_427), .B(n_393), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_418), .A2(n_388), .B(n_379), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_423), .B(n_391), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_430), .B(n_393), .Y(n_439) );
INVxp33_ASAP7_75t_L g440 ( .A(n_404), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_423), .B(n_391), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_416), .B(n_386), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_398), .B(n_383), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_398), .B(n_383), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_402), .B(n_379), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_405), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_412), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_399), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_400), .B(n_382), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_416), .B(n_386), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_409), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_405), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_399), .B(n_385), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_420), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_401), .B(n_385), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_424), .B(n_373), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_428), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_407), .B(n_320), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_401), .B(n_353), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_428), .B(n_377), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_420), .Y(n_465) );
OAI321xp33_ASAP7_75t_L g466 ( .A1(n_424), .A2(n_263), .A3(n_312), .B1(n_249), .B2(n_363), .C(n_235), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_422), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_400), .B(n_365), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_422), .Y(n_469) );
NAND2xp33_ASAP7_75t_L g470 ( .A(n_400), .B(n_354), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_403), .B(n_353), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_403), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_404), .B(n_337), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_406), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_406), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_410), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_410), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_415), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_415), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_408), .B(n_308), .Y(n_480) );
AND2x4_ASAP7_75t_SL g481 ( .A(n_397), .B(n_354), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_411), .B(n_353), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_437), .B(n_397), .Y(n_483) );
AND2x2_ASAP7_75t_SL g484 ( .A(n_470), .B(n_481), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_457), .B(n_425), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_435), .B(n_400), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_432), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_457), .B(n_415), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_437), .B(n_397), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_444), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_408), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_441), .B(n_411), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_440), .B(n_442), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_446), .Y(n_496) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_432), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_448), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_449), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_480), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_448), .B(n_415), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_481), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_460), .B(n_429), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_442), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_460), .B(n_429), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_440), .B(n_421), .Y(n_506) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_453), .B(n_400), .C(n_419), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_468), .B(n_421), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_465), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_452), .B(n_421), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_449), .Y(n_511) );
AO21x1_ASAP7_75t_L g512 ( .A1(n_451), .A2(n_414), .B(n_431), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_467), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_452), .B(n_421), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_439), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_469), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_450), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_436), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_456), .B(n_414), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_470), .B(n_417), .Y(n_520) );
NAND4xp25_ASAP7_75t_SL g521 ( .A(n_443), .B(n_431), .C(n_318), .D(n_417), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_438), .B(n_414), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_454), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_455), .B(n_417), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_458), .B(n_304), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_461), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_450), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_472), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_456), .B(n_324), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_445), .B(n_353), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_447), .B(n_360), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_462), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_474), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_474), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_476), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_459), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_472), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_459), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_464), .A2(n_266), .B1(n_322), .B2(n_315), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_475), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_504), .B(n_482), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_484), .A2(n_434), .B(n_473), .C(n_466), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_537), .B(n_479), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_500), .B(n_475), .Y(n_545) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_497), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_515), .B(n_482), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_539), .B(n_477), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_492), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_494), .B(n_477), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_519), .B(n_471), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_491), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_509), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_493), .B(n_479), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_483), .B(n_463), .Y(n_556) );
OR2x6_ASAP7_75t_L g557 ( .A(n_508), .B(n_478), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_491), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_513), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_490), .B(n_463), .Y(n_560) );
BUFx2_ASAP7_75t_SL g561 ( .A(n_502), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_516), .B(n_471), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_532), .B(n_266), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_518), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_523), .B(n_478), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_495), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_510), .B(n_357), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_521), .A2(n_312), .B1(n_315), .B2(n_297), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_514), .B(n_338), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_506), .B(n_338), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_503), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_505), .B(n_297), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_496), .B(n_249), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_524), .B(n_338), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_486), .B(n_324), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_522), .B(n_311), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_498), .B(n_305), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_526), .Y(n_578) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_527), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_533), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_507), .A2(n_322), .B(n_324), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_522), .B(n_305), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_534), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_535), .B(n_334), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_536), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_524), .B(n_311), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_541), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_531), .B(n_311), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_527), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_488), .B(n_302), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_531), .B(n_302), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_499), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_511), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_561), .B(n_485), .Y(n_594) );
NOR2xp33_ASAP7_75t_SL g595 ( .A(n_546), .B(n_507), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_563), .B(n_540), .C(n_485), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_549), .B(n_530), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_545), .B(n_529), .Y(n_598) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_543), .A2(n_512), .B(n_540), .C(n_489), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_542), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_547), .B(n_489), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_552), .A2(n_501), .B(n_525), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_552), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_581), .B(n_558), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_553), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_554), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_555), .B(n_501), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_551), .B(n_538), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_574), .B(n_520), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_559), .B(n_529), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_564), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_573), .B(n_525), .C(n_538), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_574), .B(n_528), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_578), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_584), .B(n_517), .C(n_248), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_566), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_575), .B(n_323), .C(n_254), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_592), .Y(n_618) );
NOR2x1p5_ASAP7_75t_L g619 ( .A(n_579), .B(n_269), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_544), .B(n_323), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_571), .B(n_322), .Y(n_621) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_557), .B(n_269), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_589), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_544), .B(n_288), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_550), .B(n_269), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_557), .B(n_259), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g628 ( .A1(n_568), .A2(n_259), .B(n_289), .C(n_267), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_583), .Y(n_629) );
NAND2xp33_ASAP7_75t_L g630 ( .A(n_612), .B(n_548), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_601), .B(n_562), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_600), .A2(n_557), .B1(n_556), .B2(n_560), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_596), .A2(n_567), .B1(n_585), .B2(n_587), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_604), .A2(n_569), .B(n_576), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_605), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_599), .A2(n_565), .B1(n_593), .B2(n_586), .C(n_582), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_594), .B(n_573), .C(n_588), .Y(n_637) );
INVxp67_ASAP7_75t_SL g638 ( .A(n_612), .Y(n_638) );
AOI31xp33_ASAP7_75t_L g639 ( .A1(n_627), .A2(n_570), .A3(n_572), .B(n_591), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_607), .B(n_590), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_608), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_603), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_606), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_622), .B(n_570), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_602), .A2(n_577), .B(n_279), .Y(n_645) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_623), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_596), .A2(n_282), .B1(n_265), .B2(n_287), .Y(n_647) );
OAI322xp33_ASAP7_75t_L g648 ( .A1(n_597), .A2(n_237), .A3(n_243), .B1(n_261), .B2(n_282), .C1(n_623), .C2(n_614), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_618), .B(n_611), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_616), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_626), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_636), .B(n_628), .C(n_624), .Y(n_652) );
AO22x2_ASAP7_75t_L g653 ( .A1(n_638), .A2(n_629), .B1(n_609), .B2(n_613), .Y(n_653) );
NAND4xp25_ASAP7_75t_SL g654 ( .A(n_633), .B(n_595), .C(n_615), .D(n_620), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_651), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_641), .Y(n_656) );
INVx2_ASAP7_75t_SL g657 ( .A(n_649), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_637), .A2(n_598), .B1(n_610), .B2(n_621), .Y(n_658) );
NOR3x2_ASAP7_75t_L g659 ( .A(n_630), .B(n_619), .C(n_617), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_635), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_634), .B(n_625), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_644), .B(n_642), .Y(n_662) );
NAND4xp75_ASAP7_75t_L g663 ( .A(n_631), .B(n_640), .C(n_650), .D(n_643), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_646), .Y(n_664) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_652), .B(n_647), .C(n_637), .D(n_642), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_664), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_664), .Y(n_667) );
AND3x2_ASAP7_75t_L g668 ( .A(n_662), .B(n_648), .C(n_639), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_662), .Y(n_669) );
NOR4xp25_ASAP7_75t_L g670 ( .A(n_654), .B(n_632), .C(n_645), .D(n_655), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_653), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_669), .A2(n_661), .B1(n_663), .B2(n_653), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_670), .A2(n_657), .B1(n_661), .B2(n_660), .C(n_656), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_671), .B(n_658), .C(n_659), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_671), .A2(n_656), .B1(n_667), .B2(n_666), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_675), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_672), .B(n_668), .Y(n_677) );
XNOR2xp5_ASAP7_75t_L g678 ( .A(n_674), .B(n_665), .Y(n_678) );
OA21x2_ASAP7_75t_L g679 ( .A1(n_677), .A2(n_673), .B(n_676), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_678), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_680), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_679), .B(n_678), .Y(n_682) );
endmodule