module fake_jpeg_7269_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx8_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_9),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_13),
.B1(n_8),
.B2(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_16),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_20),
.B(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_11),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_26),
.B(n_17),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_42),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_14),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_19),
.B1(n_12),
.B2(n_11),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_17),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_43),
.C(n_42),
.Y(n_50)
);

OAI321xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_10),
.A3(n_13),
.B1(n_8),
.B2(n_9),
.C(n_6),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.C(n_22),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

OAI321xp33_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_2),
.C(n_1),
.Y(n_54)
);

BUFx24_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_56),
.B(n_50),
.C(n_3),
.D(n_2),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_1),
.Y(n_60)
);


endmodule