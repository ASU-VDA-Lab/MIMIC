module fake_aes_7698_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_10;
wire n_7;
INVx2_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx3_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_0), .B(n_1), .Y(n_5) );
AND2x2_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
OAI21xp5_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
NOR2x1_ASAP7_75t_L g11 ( .A(n_9), .B(n_7), .Y(n_11) );
XOR2x2_ASAP7_75t_L g12 ( .A(n_11), .B(n_2), .Y(n_12) );
OAI211xp5_ASAP7_75t_L g13 ( .A1(n_10), .A2(n_5), .B(n_3), .C(n_2), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
OAI321xp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_13), .A3(n_5), .B1(n_12), .B2(n_1), .C(n_2), .Y(n_15) );
endmodule