module fake_jpeg_17686_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_15),
.CON(n_26),
.SN(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_19),
.B(n_18),
.C(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_10),
.Y(n_36)
);

AOI22x1_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_37),
.B1(n_25),
.B2(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_20),
.B1(n_11),
.B2(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_11),
.B1(n_20),
.B2(n_25),
.Y(n_47)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_30),
.B(n_22),
.C(n_17),
.D(n_29),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_27),
.C(n_23),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_23),
.C(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_14),
.B1(n_23),
.B2(n_2),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_14),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_22),
.B(n_17),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_29),
.C(n_27),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_10),
.C(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVxp33_ASAP7_75t_SL g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_68),
.B1(n_0),
.B2(n_2),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_10),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_55),
.B1(n_41),
.B2(n_40),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_48),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_64),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_78),
.B(n_61),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_81),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_67),
.B1(n_62),
.B2(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_46),
.Y(n_79)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_85),
.B(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_85),
.B1(n_68),
.B2(n_75),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_70),
.B(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_56),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_74),
.C(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_74),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_95),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_90),
.B(n_93),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_102),
.B(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_103),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_96),
.B(n_99),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_78),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.C(n_3),
.Y(n_107)
);

AOI21x1_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_3),
.B(n_4),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.C(n_3),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_57),
.B(n_4),
.C(n_5),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_7),
.Y(n_110)
);


endmodule