module fake_jpeg_9600_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_34),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_30),
.B1(n_28),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_20),
.B1(n_19),
.B2(n_22),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_28),
.B1(n_20),
.B2(n_17),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_73),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_85),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_75),
.B(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_97),
.B1(n_23),
.B2(n_27),
.Y(n_117)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_21),
.B1(n_29),
.B2(n_17),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_18),
.B(n_22),
.C(n_23),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_34),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_34),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_21),
.B1(n_20),
.B2(n_33),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_26),
.B1(n_25),
.B2(n_33),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_69),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_104),
.B1(n_111),
.B2(n_80),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_59),
.B1(n_57),
.B2(n_66),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_120),
.B1(n_83),
.B2(n_24),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_65),
.C(n_64),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_57),
.B1(n_66),
.B2(n_60),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_61),
.C(n_55),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_94),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_95),
.B(n_72),
.C(n_89),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_60),
.B1(n_51),
.B2(n_58),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_125),
.B1(n_126),
.B2(n_81),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_85),
.B(n_42),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_74),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_31),
.B1(n_25),
.B2(n_26),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_31),
.B1(n_27),
.B2(n_24),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_72),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_84),
.C(n_1),
.Y(n_188)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_136),
.Y(n_181)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_139),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_84),
.B1(n_82),
.B2(n_9),
.Y(n_183)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_72),
.B1(n_89),
.B2(n_91),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_16),
.B(n_15),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_146),
.B1(n_101),
.B2(n_110),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_71),
.B1(n_92),
.B2(n_90),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_150),
.B1(n_67),
.B2(n_32),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_83),
.B1(n_94),
.B2(n_88),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_147),
.B(n_16),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_154),
.B1(n_9),
.B2(n_16),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_89),
.B1(n_88),
.B2(n_85),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_155),
.Y(n_185)
);

AO21x2_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_104),
.B(n_102),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_106),
.B1(n_109),
.B2(n_113),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_121),
.B(n_105),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_117),
.B1(n_102),
.B2(n_119),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_177),
.B(n_140),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_159),
.A2(n_0),
.B(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_160),
.B(n_166),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_167),
.B1(n_170),
.B2(n_175),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_168),
.B1(n_176),
.B2(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_99),
.B1(n_109),
.B2(n_106),
.Y(n_167)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_106),
.B1(n_108),
.B2(n_113),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_106),
.B1(n_79),
.B2(n_126),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_14),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_174),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_32),
.B(n_67),
.C(n_55),
.D(n_61),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_79),
.B1(n_27),
.B2(n_24),
.Y(n_175)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_67),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_187),
.C(n_188),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_84),
.B1(n_82),
.B2(n_2),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_137),
.B1(n_134),
.B2(n_127),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_138),
.A2(n_143),
.B1(n_130),
.B2(n_137),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_141),
.B1(n_127),
.B2(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_130),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_186),
.B(n_150),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_133),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_197),
.B(n_199),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_139),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_208),
.B(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_205),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_176),
.B1(n_158),
.B2(n_172),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_207),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_129),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_217),
.B1(n_177),
.B2(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_148),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_167),
.B1(n_187),
.B2(n_177),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_0),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_3),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_231),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_178),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_216),
.A2(n_163),
.B1(n_168),
.B2(n_173),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_163),
.B1(n_158),
.B2(n_170),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_224),
.B(n_197),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_194),
.B1(n_203),
.B2(n_204),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_166),
.B1(n_159),
.B2(n_162),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_162),
.B1(n_188),
.B2(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_9),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_15),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_241),
.C(n_245),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_10),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_190),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_211),
.B(n_212),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_202),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_4),
.C(n_5),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_213),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_192),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_257),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_200),
.B(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

OAI22x1_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_267),
.B1(n_196),
.B2(n_217),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_214),
.B1(n_195),
.B2(n_197),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_228),
.B1(n_227),
.B2(n_243),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_199),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_263),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_208),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_266),
.C(n_233),
.Y(n_268)
);

XOR2x2_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_229),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_197),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_191),
.C(n_206),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_196),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_232),
.C(n_234),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_274),
.C(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_284),
.B(n_255),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_266),
.C(n_261),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_241),
.C(n_239),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_227),
.B1(n_220),
.B2(n_191),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_267),
.B1(n_253),
.B2(n_237),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_231),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

BUFx12_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_219),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_220),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_235),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_245),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_282),
.A2(n_252),
.B(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_284),
.B(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_295),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_262),
.C(n_256),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_293),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_294),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_250),
.C(n_226),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_235),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_226),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_250),
.C(n_267),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_273),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_270),
.B1(n_280),
.B2(n_272),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_306),
.B1(n_290),
.B2(n_299),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_274),
.B1(n_276),
.B2(n_275),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_293),
.Y(n_314)
);

NOR2x1_ASAP7_75t_R g308 ( 
.A(n_288),
.B(n_279),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_308),
.A2(n_285),
.B(n_12),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_242),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_311),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_10),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_298),
.Y(n_313)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_320),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_285),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_305),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_302),
.B(n_308),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_304),
.B(n_12),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_326),
.B(n_327),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_317),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_309),
.B(n_306),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_300),
.B(n_13),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_329),
.A2(n_330),
.B(n_322),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_15),
.C(n_6),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_328),
.B(n_321),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_8),
.B1(n_328),
.B2(n_329),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_8),
.Y(n_335)
);


endmodule