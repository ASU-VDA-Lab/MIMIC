module real_aes_1468_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_0), .B(n_142), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_1), .A2(n_151), .B(n_156), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_2), .B(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_3), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_4), .B(n_158), .Y(n_196) );
INVx1_ASAP7_75t_L g149 ( .A(n_5), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_6), .B(n_158), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_7), .B(n_168), .Y(n_551) );
INVx1_ASAP7_75t_L g531 ( .A(n_8), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_9), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g810 ( .A(n_10), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_11), .Y(n_497) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_12), .B(n_160), .Y(n_185) );
INVx2_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_14), .A2(n_27), .B1(n_142), .B2(n_151), .C(n_232), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_15), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_16), .B(n_142), .Y(n_181) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_17), .A2(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g559 ( .A(n_18), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_19), .B(n_162), .Y(n_235) );
INVxp33_ASAP7_75t_L g812 ( .A(n_20), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_21), .B(n_158), .Y(n_172) );
AO21x1_ASAP7_75t_L g191 ( .A1(n_22), .A2(n_142), .B(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g118 ( .A(n_23), .Y(n_118) );
INVx1_ASAP7_75t_L g557 ( .A(n_24), .Y(n_557) );
INVx1_ASAP7_75t_SL g479 ( .A(n_25), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_26), .B(n_143), .Y(n_547) );
NAND2x1_ASAP7_75t_L g204 ( .A(n_28), .B(n_158), .Y(n_204) );
AOI33xp33_ASAP7_75t_L g517 ( .A1(n_29), .A2(n_55), .A3(n_462), .B1(n_467), .B2(n_518), .B3(n_519), .Y(n_517) );
NAND2x1_ASAP7_75t_L g223 ( .A(n_30), .B(n_160), .Y(n_223) );
INVx1_ASAP7_75t_L g490 ( .A(n_31), .Y(n_490) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_32), .A2(n_88), .B(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g164 ( .A(n_32), .B(n_88), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_33), .B(n_470), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_34), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_35), .B(n_158), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_36), .B(n_160), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_37), .A2(n_151), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g148 ( .A(n_38), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g152 ( .A(n_38), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g461 ( .A(n_38), .Y(n_461) );
OR2x6_ASAP7_75t_L g116 ( .A(n_39), .B(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_40), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_41), .B(n_142), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_42), .B(n_470), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_43), .A2(n_137), .B1(n_168), .B2(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_44), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_45), .B(n_143), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_46), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_47), .B(n_160), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_48), .B(n_179), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_49), .B(n_143), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_50), .A2(n_151), .B(n_222), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_51), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_52), .A2(n_85), .B1(n_796), .B2(n_797), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_52), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_53), .A2(n_80), .B1(n_779), .B2(n_780), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_53), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_54), .B(n_160), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_56), .B(n_143), .Y(n_508) );
INVx1_ASAP7_75t_L g145 ( .A(n_57), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_57), .Y(n_155) );
AND2x2_ASAP7_75t_L g509 ( .A(n_58), .B(n_162), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_59), .A2(n_75), .B1(n_459), .B2(n_470), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_60), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_61), .B(n_158), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_62), .B(n_137), .Y(n_499) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_63), .A2(n_459), .B(n_464), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_64), .A2(n_151), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g554 ( .A(n_65), .Y(n_554) );
AO21x1_ASAP7_75t_L g193 ( .A1(n_66), .A2(n_151), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_67), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g507 ( .A(n_68), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_69), .B(n_142), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_70), .A2(n_459), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g216 ( .A(n_71), .B(n_163), .Y(n_216) );
INVx1_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
INVx1_ASAP7_75t_L g153 ( .A(n_72), .Y(n_153) );
AND2x2_ASAP7_75t_L g227 ( .A(n_73), .B(n_136), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_74), .B(n_470), .Y(n_520) );
AND2x2_ASAP7_75t_L g481 ( .A(n_76), .B(n_136), .Y(n_481) );
INVx1_ASAP7_75t_L g555 ( .A(n_77), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_78), .A2(n_459), .B(n_478), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_79), .A2(n_459), .B(n_512), .C(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_80), .Y(n_779) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
AND2x2_ASAP7_75t_L g135 ( .A(n_82), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_83), .B(n_142), .Y(n_174) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_84), .B(n_136), .Y(n_456) );
INVx1_ASAP7_75t_L g796 ( .A(n_85), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_86), .A2(n_459), .B1(n_515), .B2(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_L g192 ( .A(n_87), .B(n_168), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_89), .B(n_160), .Y(n_173) );
AND2x2_ASAP7_75t_L g208 ( .A(n_90), .B(n_136), .Y(n_208) );
INVx1_ASAP7_75t_L g465 ( .A(n_91), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_92), .B(n_158), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_93), .A2(n_151), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_94), .B(n_160), .Y(n_233) );
AND2x2_ASAP7_75t_L g521 ( .A(n_95), .B(n_136), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_96), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_97), .A2(n_488), .B(n_489), .C(n_492), .Y(n_487) );
BUFx2_ASAP7_75t_L g106 ( .A(n_98), .Y(n_106) );
BUFx2_ASAP7_75t_SL g791 ( .A(n_98), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_99), .A2(n_151), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_100), .B(n_143), .Y(n_468) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_803), .B(n_811), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_121), .B(n_789), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_108), .A2(n_793), .B(n_800), .Y(n_792) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_120), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_R g802 ( .A(n_113), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x6_ASAP7_75t_SL g125 ( .A(n_114), .B(n_116), .Y(n_125) );
OR2x6_ASAP7_75t_SL g445 ( .A(n_114), .B(n_115), .Y(n_445) );
OR2x2_ASAP7_75t_L g787 ( .A(n_114), .B(n_116), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
OAI222xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_778), .B1(n_781), .B2(n_782), .C1(n_787), .C2(n_788), .Y(n_121) );
AOI22x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B1(n_444), .B2(n_446), .Y(n_122) );
INVx3_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
CKINVDCx11_ASAP7_75t_R g786 ( .A(n_125), .Y(n_786) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g785 ( .A(n_127), .Y(n_785) );
INVx1_ASAP7_75t_L g794 ( .A(n_127), .Y(n_794) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_353), .Y(n_127) );
NOR4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_271), .C(n_297), .D(n_337), .Y(n_128) );
OAI211xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_186), .B(n_217), .C(n_257), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_165), .Y(n_131) );
AND2x2_ASAP7_75t_L g424 ( .A(n_132), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_133), .B(n_165), .Y(n_291) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g218 ( .A(n_134), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_134), .B(n_244), .Y(n_243) );
INVx5_ASAP7_75t_L g277 ( .A(n_134), .Y(n_277) );
NOR2x1_ASAP7_75t_SL g319 ( .A(n_134), .B(n_166), .Y(n_319) );
AND2x2_ASAP7_75t_L g375 ( .A(n_134), .B(n_178), .Y(n_375) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
INVx3_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_136), .A2(n_207), .B1(n_487), .B2(n_493), .Y(n_486) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_137), .B(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_139), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g168 ( .A(n_139), .B(n_164), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_150), .B(n_162), .Y(n_140) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
INVx1_ASAP7_75t_L g491 ( .A(n_143), .Y(n_491) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
AND2x6_ASAP7_75t_L g160 ( .A(n_144), .B(n_153), .Y(n_160) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g158 ( .A(n_146), .B(n_155), .Y(n_158) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx5_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_148), .Y(n_492) );
AND2x2_ASAP7_75t_L g154 ( .A(n_149), .B(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_149), .Y(n_472) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
BUFx3_ASAP7_75t_L g473 ( .A(n_152), .Y(n_473) );
INVx2_ASAP7_75t_L g463 ( .A(n_153), .Y(n_463) );
AND2x4_ASAP7_75t_L g459 ( .A(n_154), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g467 ( .A(n_155), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_161), .Y(n_156) );
INVxp67_ASAP7_75t_L g560 ( .A(n_158), .Y(n_560) );
INVxp67_ASAP7_75t_L g558 ( .A(n_160), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_161), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_161), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_161), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_161), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_161), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_161), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_161), .A2(n_233), .B(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_161), .A2(n_465), .B(n_466), .C(n_468), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_161), .A2(n_466), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_161), .A2(n_466), .B(n_507), .C(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g515 ( .A(n_161), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_161), .A2(n_466), .B(n_531), .C(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_161), .A2(n_547), .B(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_161), .B(n_168), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_162), .Y(n_226) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_162), .A2(n_231), .B(n_235), .Y(n_230) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_162), .A2(n_231), .B(n_235), .Y(n_270) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_177), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_166), .B(n_178), .Y(n_247) );
AND2x2_ASAP7_75t_L g308 ( .A(n_166), .B(n_277), .Y(n_308) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_175), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_167), .B(n_176), .Y(n_175) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_167), .A2(n_169), .B(n_175), .Y(n_261) );
INVx1_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_168), .A2(n_181), .B(n_182), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_168), .B(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_168), .A2(n_458), .B(n_469), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
AND2x2_ASAP7_75t_L g320 ( .A(n_177), .B(n_244), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_177), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g364 ( .A(n_177), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g397 ( .A(n_177), .B(n_218), .Y(n_397) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g241 ( .A(n_178), .Y(n_241) );
AND2x2_ASAP7_75t_L g274 ( .A(n_178), .B(n_275), .Y(n_274) );
BUFx3_ASAP7_75t_L g309 ( .A(n_178), .Y(n_309) );
OR2x2_ASAP7_75t_L g385 ( .A(n_178), .B(n_244), .Y(n_385) );
INVx2_ASAP7_75t_SL g512 ( .A(n_179), .Y(n_512) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_179), .A2(n_529), .B(n_533), .Y(n_528) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
AOI211x1_ASAP7_75t_SL g314 ( .A1(n_188), .A2(n_306), .B(n_315), .C(n_317), .Y(n_314) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_188), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_188), .B(n_357), .Y(n_404) );
BUFx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g229 ( .A(n_190), .Y(n_229) );
OAI21x1_ASAP7_75t_SL g190 ( .A1(n_191), .A2(n_193), .B(n_197), .Y(n_190) );
INVx1_ASAP7_75t_L g198 ( .A(n_192), .Y(n_198) );
AOI322xp5_ASAP7_75t_L g217 ( .A1(n_199), .A2(n_218), .A3(n_228), .B1(n_236), .B2(n_239), .C1(n_245), .C2(n_248), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_199), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
INVx2_ASAP7_75t_L g252 ( .A(n_200), .Y(n_252) );
INVxp67_ASAP7_75t_L g294 ( .A(n_200), .Y(n_294) );
BUFx3_ASAP7_75t_L g358 ( .A(n_200), .Y(n_358) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_207), .B(n_208), .Y(n_200) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_201), .A2(n_207), .B(n_208), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_206), .Y(n_201) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_207), .A2(n_210), .B(n_216), .Y(n_209) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_207), .A2(n_210), .B(n_216), .Y(n_256) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_207), .A2(n_503), .B(n_509), .Y(n_502) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_207), .A2(n_503), .B(n_509), .Y(n_525) );
INVx2_ASAP7_75t_L g267 ( .A(n_209), .Y(n_267) );
AND2x2_ASAP7_75t_L g316 ( .A(n_209), .B(n_230), .Y(n_316) );
AND2x2_ASAP7_75t_L g360 ( .A(n_209), .B(n_269), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_211), .B(n_215), .Y(n_210) );
AND2x2_ASAP7_75t_L g245 ( .A(n_218), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_218), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_218), .B(n_274), .Y(n_439) );
INVx4_ASAP7_75t_L g244 ( .A(n_219), .Y(n_244) );
AND2x2_ASAP7_75t_L g276 ( .A(n_219), .B(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_219), .Y(n_329) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_226), .B(n_227), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_226), .A2(n_475), .B(n_481), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_228), .B(n_313), .Y(n_338) );
INVx1_ASAP7_75t_SL g377 ( .A(n_228), .Y(n_377) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AND2x4_ASAP7_75t_L g268 ( .A(n_229), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_229), .B(n_267), .Y(n_336) );
AND2x2_ASAP7_75t_L g388 ( .A(n_229), .B(n_238), .Y(n_388) );
OR2x2_ASAP7_75t_L g412 ( .A(n_229), .B(n_230), .Y(n_412) );
AND2x2_ASAP7_75t_L g236 ( .A(n_230), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g286 ( .A(n_230), .B(n_267), .Y(n_286) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_230), .B(n_254), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_236), .B(n_349), .Y(n_366) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
BUFx2_ASAP7_75t_L g301 ( .A(n_238), .Y(n_301) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_238), .B(n_255), .Y(n_341) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
OR2x2_ASAP7_75t_L g289 ( .A(n_240), .B(n_243), .Y(n_289) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g258 ( .A(n_241), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g406 ( .A(n_241), .B(n_319), .Y(n_406) );
AND2x2_ASAP7_75t_L g422 ( .A(n_241), .B(n_276), .Y(n_422) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AOI311xp33_ASAP7_75t_L g392 ( .A1(n_243), .A2(n_331), .A3(n_393), .B(n_395), .C(n_402), .Y(n_392) );
AND2x4_ASAP7_75t_L g259 ( .A(n_244), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g263 ( .A(n_244), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_244), .B(n_277), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_244), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g376 ( .A(n_244), .B(n_363), .Y(n_376) );
AND2x2_ASAP7_75t_L g262 ( .A(n_246), .B(n_263), .Y(n_262) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
INVxp67_ASAP7_75t_SL g280 ( .A(n_247), .Y(n_280) );
OR2x2_ASAP7_75t_L g369 ( .A(n_247), .B(n_333), .Y(n_369) );
INVx1_ASAP7_75t_L g425 ( .A(n_247), .Y(n_425) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g334 ( .A(n_251), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g348 ( .A(n_251), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g423 ( .A(n_251), .B(n_296), .Y(n_423) );
BUFx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g266 ( .A(n_252), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g285 ( .A(n_252), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g347 ( .A(n_253), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_253), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_402) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g296 ( .A(n_254), .B(n_267), .Y(n_296) );
AND2x4_ASAP7_75t_L g349 ( .A(n_254), .B(n_256), .Y(n_349) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI21xp33_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_262), .B(n_264), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_258), .A2(n_344), .B1(n_348), .B2(n_350), .Y(n_343) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_259), .B(n_277), .Y(n_303) );
INVx2_ASAP7_75t_L g365 ( .A(n_259), .Y(n_365) );
AND2x2_ASAP7_75t_L g379 ( .A(n_259), .B(n_375), .Y(n_379) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g275 ( .A(n_261), .Y(n_275) );
INVx1_ASAP7_75t_L g328 ( .A(n_261), .Y(n_328) );
INVx1_ASAP7_75t_L g279 ( .A(n_263), .Y(n_279) );
AND3x2_ASAP7_75t_L g307 ( .A(n_263), .B(n_308), .C(n_309), .Y(n_307) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g371 ( .A(n_266), .Y(n_371) );
AND2x2_ASAP7_75t_L g299 ( .A(n_268), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g370 ( .A(n_268), .B(n_371), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_268), .A2(n_382), .B1(n_386), .B2(n_389), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_268), .B(n_416), .Y(n_420) );
BUFx2_ASAP7_75t_L g311 ( .A(n_269), .Y(n_311) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g282 ( .A(n_270), .Y(n_282) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_270), .Y(n_401) );
OAI221xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_281), .B1(n_283), .B2(n_284), .C(n_287), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_278), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g363 ( .A(n_275), .Y(n_363) );
INVx2_ASAP7_75t_SL g352 ( .A(n_276), .Y(n_352) );
AND2x2_ASAP7_75t_L g434 ( .A(n_276), .B(n_301), .Y(n_434) );
INVx4_ASAP7_75t_L g325 ( .A(n_277), .Y(n_325) );
INVx1_ASAP7_75t_L g283 ( .A(n_278), .Y(n_283) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x4_ASAP7_75t_L g394 ( .A(n_282), .B(n_349), .Y(n_394) );
INVx1_ASAP7_75t_SL g433 ( .A(n_282), .Y(n_433) );
AND2x2_ASAP7_75t_L g438 ( .A(n_282), .B(n_341), .Y(n_438) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g380 ( .A(n_286), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_290), .B(n_292), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g313 ( .A(n_294), .Y(n_313) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g310 ( .A(n_296), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g400 ( .A(n_296), .B(n_401), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_302), .B(n_304), .C(n_321), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g393 ( .A(n_300), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_301), .B(n_316), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_301), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g426 ( .A(n_301), .B(n_349), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g337 ( .A1(n_302), .A2(n_326), .B1(n_338), .B2(n_339), .C(n_343), .Y(n_337) );
INVx3_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g408 ( .A(n_303), .B(n_309), .Y(n_408) );
OAI32xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_310), .A3(n_312), .B1(n_314), .B2(n_318), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_308), .Y(n_398) );
INVx2_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_309), .A2(n_361), .B(n_441), .C(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g346 ( .A(n_311), .Y(n_346) );
OR2x2_ASAP7_75t_L g442 ( .A(n_311), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_315), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g403 ( .A(n_318), .Y(n_403) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g384 ( .A(n_319), .Y(n_384) );
OAI21xp33_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_330), .B(n_334), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
OR2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_325), .B(n_328), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_327), .A2(n_359), .B1(n_428), .B2(n_431), .C(n_435), .Y(n_427) );
INVx2_ASAP7_75t_L g430 ( .A(n_327), .Y(n_430) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OR2x2_ASAP7_75t_L g351 ( .A(n_331), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g418 ( .A(n_331), .B(n_376), .Y(n_418) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g416 ( .A(n_341), .Y(n_416) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_349), .B(n_379), .Y(n_436) );
INVx2_ASAP7_75t_L g443 ( .A(n_349), .Y(n_443) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_351), .A2(n_414), .B1(n_417), .B2(n_419), .C(n_421), .Y(n_413) );
AND5x1_ASAP7_75t_L g353 ( .A(n_354), .B(n_392), .C(n_407), .D(n_427), .E(n_437), .Y(n_353) );
NOR2xp33_ASAP7_75t_SL g354 ( .A(n_355), .B(n_372), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_361), .B1(n_364), .B2(n_366), .C(n_367), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_377), .B1(n_378), .B2(n_380), .C(n_381), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_377), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
OR2x2_ASAP7_75t_L g390 ( .A(n_385), .B(n_391), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B(n_399), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B(n_413), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_424), .B2(n_426), .Y(n_421) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_423), .A2(n_438), .B(n_439), .C(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g441 ( .A(n_434), .Y(n_441) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g784 ( .A(n_444), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
OAI22x1_ASAP7_75t_L g783 ( .A1(n_446), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_783) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
AND3x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_668), .C(n_731), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_632), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_573), .C(n_602), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_452), .B(n_562), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_482), .B1(n_522), .B2(n_534), .Y(n_452) );
NAND2x1_ASAP7_75t_L g717 ( .A(n_453), .B(n_563), .Y(n_717) );
INVx2_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_474), .Y(n_454) );
INVx2_ASAP7_75t_L g536 ( .A(n_455), .Y(n_536) );
INVx4_ASAP7_75t_L g578 ( .A(n_455), .Y(n_578) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_455), .Y(n_598) );
AND2x4_ASAP7_75t_L g609 ( .A(n_455), .B(n_577), .Y(n_609) );
AND2x2_ASAP7_75t_L g615 ( .A(n_455), .B(n_539), .Y(n_615) );
NOR2x1_ASAP7_75t_SL g745 ( .A(n_455), .B(n_550), .Y(n_745) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVxp67_ASAP7_75t_L g498 ( .A(n_459), .Y(n_498) );
NOR2x1p5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g519 ( .A(n_462), .Y(n_519) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x6_ASAP7_75t_L g466 ( .A(n_463), .B(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g488 ( .A(n_466), .Y(n_488) );
INVx2_ASAP7_75t_L g549 ( .A(n_466), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_466), .A2(n_491), .B1(n_554), .B2(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g471 ( .A(n_467), .B(n_472), .Y(n_471) );
INVxp33_ASAP7_75t_L g518 ( .A(n_467), .Y(n_518) );
INVx1_ASAP7_75t_L g500 ( .A(n_470), .Y(n_500) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g542 ( .A(n_471), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
INVx2_ASAP7_75t_L g581 ( .A(n_474), .Y(n_581) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_474), .Y(n_595) );
INVx1_ASAP7_75t_L g606 ( .A(n_474), .Y(n_606) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_474), .Y(n_618) );
AND2x2_ASAP7_75t_L g650 ( .A(n_474), .B(n_550), .Y(n_650) );
AND2x2_ASAP7_75t_L g682 ( .A(n_474), .B(n_566), .Y(n_682) );
INVx1_ASAP7_75t_L g689 ( .A(n_474), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_501), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g631 ( .A(n_484), .B(n_570), .Y(n_631) );
INVx2_ASAP7_75t_L g705 ( .A(n_484), .Y(n_705) );
AND2x2_ASAP7_75t_L g728 ( .A(n_484), .B(n_501), .Y(n_728) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_485), .B(n_525), .Y(n_569) );
INVx2_ASAP7_75t_L g590 ( .A(n_485), .Y(n_590) );
AND2x4_ASAP7_75t_L g612 ( .A(n_485), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g647 ( .A(n_485), .Y(n_647) );
AND2x2_ASAP7_75t_L g724 ( .A(n_485), .B(n_528), .Y(n_724) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g695 ( .A(n_501), .Y(n_695) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
NOR2xp67_ASAP7_75t_L g620 ( .A(n_502), .B(n_590), .Y(n_620) );
AND2x2_ASAP7_75t_L g625 ( .A(n_502), .B(n_590), .Y(n_625) );
INVx2_ASAP7_75t_L g638 ( .A(n_502), .Y(n_638) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_502), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AND2x4_ASAP7_75t_L g611 ( .A(n_510), .B(n_524), .Y(n_611) );
AND2x2_ASAP7_75t_L g626 ( .A(n_510), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g679 ( .A(n_510), .Y(n_679) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_511), .B(n_528), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_511), .B(n_525), .Y(n_683) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_521), .Y(n_511) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_512), .A2(n_513), .B(n_521), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_514), .B(n_520), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVxp33_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
INVx3_ASAP7_75t_L g587 ( .A(n_524), .Y(n_587) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
AND2x2_ASAP7_75t_L g754 ( .A(n_525), .B(n_755), .Y(n_754) );
INVx3_ASAP7_75t_L g642 ( .A(n_526), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_526), .B(n_679), .Y(n_774) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g589 ( .A(n_527), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g570 ( .A(n_528), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g613 ( .A(n_528), .Y(n_613) );
INVxp67_ASAP7_75t_L g627 ( .A(n_528), .Y(n_627) );
INVx1_ASAP7_75t_L g687 ( .A(n_528), .Y(n_687) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_528), .Y(n_755) );
INVx1_ASAP7_75t_L g739 ( .A(n_534), .Y(n_739) );
NOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_535), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g693 ( .A(n_536), .B(n_565), .Y(n_693) );
OR2x2_ASAP7_75t_L g729 ( .A(n_537), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g711 ( .A(n_538), .B(n_689), .Y(n_711) );
AND2x2_ASAP7_75t_L g763 ( .A(n_538), .B(n_598), .Y(n_763) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_550), .Y(n_538) );
AND2x4_ASAP7_75t_L g565 ( .A(n_539), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g577 ( .A(n_539), .Y(n_577) );
INVx2_ASAP7_75t_L g594 ( .A(n_539), .Y(n_594) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_539), .Y(n_772) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_545), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .C(n_544), .Y(n_541) );
INVx3_ASAP7_75t_L g566 ( .A(n_550), .Y(n_566) );
INVx2_ASAP7_75t_L g660 ( .A(n_550), .Y(n_660) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_556), .B(n_561), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B1(n_559), .B2(n_560), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_564), .B(n_640), .Y(n_657) );
NOR2x1_ASAP7_75t_L g699 ( .A(n_564), .B(n_578), .Y(n_699) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_565), .B(n_640), .Y(n_777) );
AND2x2_ASAP7_75t_L g593 ( .A(n_566), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g607 ( .A(n_566), .Y(n_607) );
AOI22xp5_ASAP7_75t_SL g655 ( .A1(n_567), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_568), .B(n_626), .Y(n_652) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g713 ( .A(n_569), .B(n_601), .Y(n_713) );
AND2x2_ASAP7_75t_L g583 ( .A(n_570), .B(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g619 ( .A(n_570), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g715 ( .A(n_570), .B(n_705), .Y(n_715) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g637 ( .A(n_572), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g663 ( .A(n_572), .Y(n_663) );
AND2x2_ASAP7_75t_L g753 ( .A(n_572), .B(n_590), .Y(n_753) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_582), .B1(n_586), .B2(n_591), .C(n_596), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g654 ( .A(n_576), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_576), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_576), .B(n_650), .Y(n_769) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NOR2xp67_ASAP7_75t_SL g622 ( .A(n_578), .B(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_578), .Y(n_635) );
OR2x2_ASAP7_75t_L g719 ( .A(n_578), .B(n_720), .Y(n_719) );
AND2x4_ASAP7_75t_SL g771 ( .A(n_578), .B(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g640 ( .A(n_580), .Y(n_640) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_581), .Y(n_730) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI221x1_ASAP7_75t_L g670 ( .A1(n_583), .A2(n_671), .B1(n_673), .B2(n_676), .C(n_680), .Y(n_670) );
AND2x2_ASAP7_75t_L g656 ( .A(n_584), .B(n_612), .Y(n_656) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
AND2x2_ASAP7_75t_L g599 ( .A(n_587), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_587), .B(n_589), .Y(n_726) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_593), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_593), .B(n_606), .Y(n_623) );
INVx2_ASAP7_75t_L g630 ( .A(n_593), .Y(n_630) );
INVx1_ASAP7_75t_L g675 ( .A(n_594), .Y(n_675) );
BUFx2_ASAP7_75t_L g764 ( .A(n_595), .Y(n_764) );
NAND2xp33_ASAP7_75t_SL g596 ( .A(n_597), .B(n_599), .Y(n_596) );
OR2x6_ASAP7_75t_L g629 ( .A(n_598), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g710 ( .A(n_598), .B(n_650), .Y(n_710) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_621), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_610), .B1(n_614), .B2(n_619), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
AND2x2_ASAP7_75t_SL g667 ( .A(n_605), .B(n_609), .Y(n_667) );
AND2x4_ASAP7_75t_L g673 ( .A(n_605), .B(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_SL g605 ( .A(n_606), .B(n_607), .Y(n_605) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_606), .Y(n_698) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_609), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_609), .B(n_640), .Y(n_672) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_609), .Y(n_756) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g703 ( .A(n_611), .B(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g664 ( .A(n_612), .Y(n_664) );
NAND2x1_ASAP7_75t_SL g708 ( .A(n_612), .B(n_663), .Y(n_708) );
AND2x2_ASAP7_75t_L g742 ( .A(n_612), .B(n_637), .Y(n_742) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_628), .B2(n_631), .Y(n_621) );
BUFx2_ASAP7_75t_L g737 ( .A(n_623), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_624), .A2(n_693), .B1(n_767), .B2(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g678 ( .A(n_625), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g645 ( .A(n_626), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_630), .B(n_762), .C(n_764), .Y(n_761) );
INVx1_ASAP7_75t_L g665 ( .A(n_631), .Y(n_665) );
AOI211x1_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_641), .B(n_643), .C(n_661), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_636), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AND2x2_ASAP7_75t_L g723 ( .A(n_637), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_637), .B(n_704), .Y(n_735) );
AND2x2_ASAP7_75t_L g767 ( .A(n_637), .B(n_705), .Y(n_767) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g748 ( .A(n_640), .Y(n_748) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g677 ( .A(n_642), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_655), .Y(n_643) );
AOI22xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_648), .B1(n_651), .B2(n_653), .Y(n_644) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g685 ( .A(n_647), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g700 ( .A(n_647), .Y(n_700) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_SL g770 ( .A(n_650), .B(n_771), .Y(n_770) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g706 ( .A(n_659), .B(n_689), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_666), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_663), .B(n_685), .Y(n_760) );
OR2x2_ASAP7_75t_L g738 ( .A(n_664), .B(n_683), .Y(n_738) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND3x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_690), .C(n_714), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_673), .A2(n_703), .B1(n_706), .B2(n_707), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_674), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_SL g747 ( .A(n_674), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_674), .B(n_748), .Y(n_751) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI222xp33_ASAP7_75t_L g734 ( .A1(n_678), .A2(n_735), .B1(n_736), .B2(n_737), .C1(n_738), .C2(n_739), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_684), .B2(n_688), .Y(n_680) );
INVx1_ASAP7_75t_SL g720 ( .A(n_682), .Y(n_720) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g757 ( .A(n_686), .B(n_753), .Y(n_757) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_701), .Y(n_690) );
AOI21xp5_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_694), .B(n_700), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_709), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_708), .B(n_722), .Y(n_721) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_710), .A2(n_711), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g736 ( .A(n_711), .Y(n_736) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_718), .B2(n_721), .C(n_725), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NAND3x1_ASAP7_75t_L g732 ( .A(n_733), .B(n_758), .C(n_765), .Y(n_732) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_740), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_749), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_742), .B(n_743), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_744), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B1(n_756), .B2(n_757), .Y(n_749) );
AND2x4_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_775), .Y(n_765) );
AOI22xp5_ASAP7_75t_SL g766 ( .A1(n_767), .A2(n_768), .B1(n_770), .B2(n_773), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVxp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g781 ( .A(n_778), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g798 ( .A(n_785), .Y(n_798) );
INVx3_ASAP7_75t_L g807 ( .A(n_787), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
OAI22xp5_ASAP7_75t_SL g793 ( .A1(n_794), .A2(n_795), .B1(n_798), .B2(n_799), .Y(n_793) );
INVx1_ASAP7_75t_L g799 ( .A(n_795), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx4_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g813 ( .A(n_806), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
endmodule