module fake_jpeg_25196_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_33),
.B1(n_22),
.B2(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_27),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_18),
.B(n_24),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_48),
.B1(n_25),
.B2(n_21),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_0),
.B(n_1),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_33),
.B1(n_21),
.B2(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_31),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_19),
.CON(n_60),
.SN(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_34),
.B(n_19),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_40),
.B1(n_39),
.B2(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_81),
.B1(n_58),
.B2(n_47),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_44),
.B1(n_56),
.B2(n_49),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_34),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_86),
.B1(n_90),
.B2(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_84),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_33),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_46),
.B(n_50),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_16),
.B(n_22),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_95),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_110),
.B1(n_90),
.B2(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_103),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_91),
.B1(n_105),
.B2(n_108),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_55),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_61),
.C(n_62),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_108),
.C(n_86),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_43),
.C(n_56),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_48),
.B1(n_59),
.B2(n_49),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_19),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_53),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_53),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_119),
.B(n_141),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_137),
.B1(n_97),
.B2(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_125),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_128),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_59),
.B1(n_83),
.B2(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_85),
.B1(n_82),
.B2(n_16),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_92),
.A2(n_64),
.B1(n_65),
.B2(n_74),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_140),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_110),
.B1(n_112),
.B2(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_142),
.B1(n_94),
.B2(n_59),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_66),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_65),
.B1(n_20),
.B2(n_66),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_73),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_114),
.B(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_30),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_59),
.B1(n_36),
.B2(n_28),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_42),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_16),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_179),
.B(n_32),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_158),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_132),
.B1(n_135),
.B2(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_174),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_104),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_163),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_104),
.B(n_109),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_159),
.B(n_164),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_109),
.B1(n_102),
.B2(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_161),
.B(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_96),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_127),
.B(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_102),
.B1(n_28),
.B2(n_70),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_30),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_171),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_30),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_140),
.B1(n_131),
.B2(n_145),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_120),
.B1(n_20),
.B2(n_31),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_122),
.A2(n_24),
.B(n_20),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_120),
.B1(n_122),
.B2(n_125),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_188),
.B1(n_193),
.B2(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_191),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_167),
.B1(n_148),
.B2(n_160),
.Y(n_215)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_159),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_23),
.A3(n_18),
.B1(n_32),
.B2(n_42),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_199),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_156),
.C(n_163),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_200),
.C(n_170),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_166),
.Y(n_234)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_42),
.C(n_14),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_172),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_207),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_206),
.B1(n_179),
.B2(n_160),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_152),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_209),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_213),
.B(n_203),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_221),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_223),
.B1(n_189),
.B2(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_225),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_183),
.A2(n_210),
.B1(n_191),
.B2(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_168),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_230),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_158),
.C(n_159),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_185),
.C(n_209),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_162),
.B(n_150),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_231),
.C(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_199),
.B(n_197),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_171),
.B(n_150),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_223),
.B(n_211),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_219),
.B(n_235),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_187),
.B(n_192),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_234),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_205),
.B1(n_183),
.B2(n_193),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_227),
.B1(n_214),
.B2(n_203),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_174),
.C(n_184),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_215),
.C(n_222),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_253),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_206),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_224),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_203),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_3),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_266),
.C(n_271),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_256),
.B(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_3),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_219),
.C(n_212),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_273),
.B(n_247),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_244),
.B1(n_248),
.B2(n_247),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_11),
.C(n_9),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_281),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_264),
.B(n_271),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_286),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_243),
.C(n_240),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_242),
.C(n_250),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_284),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_248),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_260),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_254),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_6),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_262),
.C(n_269),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_294),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_297),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_269),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_3),
.C(n_4),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_5),
.C(n_6),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.C(n_287),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_6),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_281),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_303),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_278),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_282),
.B1(n_277),
.B2(n_274),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_300),
.B(n_305),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_292),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_314),
.B(n_298),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_289),
.B(n_7),
.Y(n_317)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_275),
.B(n_287),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_315),
.A2(n_316),
.B(n_317),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_289),
.B(n_7),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_312),
.C(n_311),
.Y(n_320)
);

NAND4xp25_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_310),
.C(n_7),
.D(n_8),
.Y(n_321)
);

NAND4xp25_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_7),
.C(n_8),
.D(n_297),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_8),
.Y(n_323)
);


endmodule