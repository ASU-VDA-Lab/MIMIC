module fake_netlist_1_4449_n_524 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_524);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_524;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_70), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_33), .Y(n_76) );
BUFx2_ASAP7_75t_SL g77 ( .A(n_73), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_12), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_41), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_38), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_37), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_42), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_61), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_49), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_40), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_39), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_60), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_34), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_2), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_15), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_28), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_23), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_62), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_53), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_52), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_24), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_21), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_44), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_71), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_46), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_50), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_65), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_59), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_80), .B(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_80), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_107), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_107), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_84), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_98), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_75), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_100), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_98), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_84), .Y(n_119) );
XOR2x2_ASAP7_75t_L g120 ( .A(n_78), .B(n_0), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_88), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_98), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_75), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_96), .B(n_1), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_99), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_94), .B(n_1), .Y(n_127) );
NOR2xp33_ASAP7_75t_SL g128 ( .A(n_81), .B(n_29), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_88), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_76), .Y(n_130) );
NOR2xp33_ASAP7_75t_SL g131 ( .A(n_102), .B(n_30), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_116), .B(n_95), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_123), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_116), .B(n_79), .Y(n_134) );
INVx4_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_130), .B(n_79), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_111), .B(n_99), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_130), .A2(n_90), .B1(n_91), .B2(n_103), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_112), .B(n_90), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_110), .B(n_93), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_123), .A2(n_91), .B1(n_103), .B2(n_77), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_112), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_125), .B(n_92), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_113), .B(n_92), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_125), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
INVx4_ASAP7_75t_SL g147 ( .A(n_115), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_114), .B(n_77), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_121), .B(n_83), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_119), .B(n_82), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_115), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_119), .B(n_82), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_118), .Y(n_156) );
NOR3x1_ASAP7_75t_L g157 ( .A(n_151), .B(n_120), .C(n_109), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_148), .A2(n_127), .B1(n_124), .B2(n_129), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
OR2x6_ASAP7_75t_L g161 ( .A(n_148), .B(n_105), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_149), .B(n_97), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_148), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_155), .B(n_131), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_149), .B(n_105), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_149), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_139), .B(n_144), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_155), .B(n_104), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_141), .A2(n_128), .B1(n_129), .B2(n_104), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_140), .B(n_117), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_141), .B(n_85), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_132), .B(n_85), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_132), .B(n_86), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_138), .A2(n_117), .B1(n_120), .B2(n_87), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_145), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_134), .B(n_86), .Y(n_181) );
NOR2xp67_ASAP7_75t_L g182 ( .A(n_135), .B(n_87), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_138), .B(n_106), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_142), .B(n_106), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_171), .A2(n_136), .B1(n_142), .B2(n_143), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_163), .A2(n_139), .B1(n_137), .B2(n_146), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_185), .A2(n_136), .B(n_143), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_169), .A2(n_146), .B(n_139), .C(n_137), .Y(n_192) );
AND3x1_ASAP7_75t_SL g193 ( .A(n_157), .B(n_2), .C(n_3), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_163), .A2(n_139), .B(n_137), .C(n_83), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_176), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_171), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_160), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_176), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_161), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_137), .B1(n_101), .B2(n_89), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_186), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_161), .A2(n_89), .B1(n_101), .B2(n_98), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_186), .B(n_98), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_165), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_158), .A2(n_108), .B1(n_152), .B2(n_122), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_167), .Y(n_211) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_186), .B(n_108), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_167), .B(n_3), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_185), .A2(n_154), .B(n_152), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_170), .B(n_4), .Y(n_216) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_169), .A2(n_154), .B(n_156), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_158), .A2(n_108), .B1(n_122), .B2(n_118), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_170), .A2(n_108), .B1(n_122), .B2(n_118), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_186), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_197), .B(n_165), .Y(n_221) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_194), .A2(n_164), .B(n_181), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_197), .Y(n_223) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_207), .A2(n_178), .B(n_177), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_203), .A2(n_179), .B1(n_172), .B2(n_166), .Y(n_225) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_192), .A2(n_182), .B(n_175), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_207), .A2(n_182), .B(n_184), .Y(n_228) );
OAI21x1_ASAP7_75t_SL g229 ( .A1(n_202), .A2(n_180), .B(n_173), .Y(n_229) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_218), .A2(n_180), .B(n_188), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_201), .Y(n_231) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_219), .A2(n_156), .B(n_150), .Y(n_232) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_204), .A2(n_168), .B(n_162), .Y(n_233) );
AO21x1_ASAP7_75t_L g234 ( .A1(n_210), .A2(n_170), .B(n_183), .Y(n_234) );
AOI21xp5_ASAP7_75t_SL g235 ( .A1(n_202), .A2(n_170), .B(n_159), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_201), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_216), .A2(n_179), .B1(n_183), .B2(n_187), .Y(n_237) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_217), .A2(n_168), .B(n_150), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_199), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_209), .B(n_159), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_217), .A2(n_168), .B(n_150), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_219), .A2(n_156), .B(n_187), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
OAI211xp5_ASAP7_75t_L g246 ( .A1(n_225), .A2(n_196), .B(n_174), .C(n_190), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_216), .B1(n_206), .B2(n_203), .Y(n_247) );
CKINVDCx6p67_ASAP7_75t_R g248 ( .A(n_231), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_223), .B(n_215), .Y(n_249) );
CKINVDCx14_ASAP7_75t_R g250 ( .A(n_231), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_221), .A2(n_215), .B(n_189), .Y(n_251) );
OAI21xp33_ASAP7_75t_L g252 ( .A1(n_237), .A2(n_212), .B(n_213), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_223), .B(n_206), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_221), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_243), .Y(n_256) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_237), .A2(n_198), .B1(n_211), .B2(n_216), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_224), .A2(n_212), .B(n_216), .C(n_191), .Y(n_258) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_208), .B(n_214), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_227), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_243), .B(n_213), .Y(n_261) );
AOI222xp33_ASAP7_75t_L g262 ( .A1(n_229), .A2(n_212), .B1(n_157), .B2(n_193), .C1(n_227), .C2(n_239), .Y(n_262) );
AOI222xp33_ASAP7_75t_L g263 ( .A1(n_229), .A2(n_205), .B1(n_200), .B2(n_195), .C1(n_220), .C2(n_201), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_234), .A2(n_205), .B1(n_195), .B2(n_220), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g265 ( .A1(n_239), .A2(n_200), .B1(n_168), .B2(n_217), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_239), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_256), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_255), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_255), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_262), .B(n_235), .C(n_108), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_256), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_260), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_266), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_248), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_250), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_254), .B(n_224), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_266), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_260), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_249), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_248), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_253), .B(n_224), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_247), .A2(n_234), .B1(n_229), .B2(n_226), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_249), .B(n_233), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_253), .B(n_245), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_261), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_267), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
OAI33xp33_ASAP7_75t_L g290 ( .A1(n_271), .A2(n_257), .A3(n_252), .B1(n_265), .B2(n_261), .B3(n_262), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_286), .B(n_246), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_270), .B(n_264), .C(n_263), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_271), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_273), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_268), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_273), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_282), .B(n_258), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_272), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_282), .B(n_231), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_263), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_280), .B(n_233), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_274), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_252), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_277), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_278), .B(n_245), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_268), .B(n_245), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_284), .A2(n_251), .B(n_240), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_269), .B(n_245), .Y(n_310) );
OAI21xp5_ASAP7_75t_SL g311 ( .A1(n_274), .A2(n_245), .B(n_240), .Y(n_311) );
AOI211xp5_ASAP7_75t_L g312 ( .A1(n_286), .A2(n_234), .B(n_228), .C(n_242), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_279), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_315), .B(n_272), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_297), .B(n_276), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_297), .B(n_276), .Y(n_321) );
AO21x1_ASAP7_75t_L g322 ( .A1(n_294), .A2(n_269), .B(n_285), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_296), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_315), .B(n_283), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_292), .A2(n_275), .B1(n_281), .B2(n_274), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_303), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_291), .B(n_285), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_316), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_299), .B(n_259), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_290), .B(n_288), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_299), .B(n_281), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_299), .B(n_281), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_316), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_308), .Y(n_337) );
NAND4xp25_ASAP7_75t_L g338 ( .A(n_312), .B(n_281), .C(n_274), .D(n_7), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_299), .B(n_4), .Y(n_339) );
AOI21xp33_ASAP7_75t_SL g340 ( .A1(n_302), .A2(n_5), .B(n_7), .Y(n_340) );
OR2x4_ASAP7_75t_L g341 ( .A(n_311), .B(n_118), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_302), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_301), .B(n_259), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_288), .B(n_231), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_308), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_313), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_306), .Y(n_348) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_312), .B(n_118), .C(n_122), .Y(n_349) );
AND3x2_ASAP7_75t_L g350 ( .A(n_300), .B(n_5), .C(n_8), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_317), .B(n_8), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_300), .A2(n_226), .B1(n_244), .B2(n_228), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_305), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_289), .B(n_236), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_305), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_301), .B(n_259), .Y(n_356) );
OR2x6_ASAP7_75t_L g357 ( .A(n_289), .B(n_242), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_293), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_293), .B(n_236), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_306), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_317), .B(n_9), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_333), .B(n_304), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_348), .B(n_304), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_320), .B(n_321), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_360), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_320), .B(n_314), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
NOR2x1p5_ASAP7_75t_L g369 ( .A(n_338), .B(n_295), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_321), .B(n_307), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_319), .B(n_307), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_333), .B(n_295), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_332), .B(n_314), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_337), .B(n_313), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_326), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_331), .B(n_314), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_328), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_336), .B(n_313), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_341), .A2(n_309), .B1(n_310), .B2(n_236), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_348), .B(n_310), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_346), .B(n_122), .Y(n_382) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_327), .B(n_244), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_329), .B(n_9), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_332), .B(n_244), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_343), .B(n_244), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_322), .B(n_241), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_347), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_325), .B(n_10), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_343), .B(n_244), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_325), .B(n_11), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_356), .B(n_232), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_339), .B(n_11), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_356), .B(n_232), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_347), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_323), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_330), .B(n_12), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_330), .B(n_13), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_358), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_351), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_348), .B(n_241), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_357), .B(n_232), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_357), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_361), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_357), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_344), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_341), .A2(n_241), .B1(n_232), .B2(n_226), .Y(n_409) );
NOR2x1_ASAP7_75t_L g410 ( .A(n_349), .B(n_232), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_342), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_352), .B(n_232), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_362), .B(n_344), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_372), .B(n_344), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_402), .A2(n_340), .B1(n_354), .B2(n_359), .C(n_342), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_398), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_368), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_364), .B(n_335), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_383), .A2(n_334), .B(n_354), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_365), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_403), .A2(n_350), .B1(n_354), .B2(n_359), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_369), .A2(n_350), .B1(n_359), .B2(n_226), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_363), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_403), .A2(n_228), .B(n_238), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_411), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_407), .A2(n_222), .B(n_230), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_364), .B(n_13), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_367), .B(n_14), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_406), .B(n_15), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_367), .B(n_16), .Y(n_431) );
AOI32xp33_ASAP7_75t_L g432 ( .A1(n_395), .A2(n_238), .A3(n_242), .B1(n_222), .B2(n_230), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_405), .A2(n_238), .B(n_222), .C(n_230), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_375), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_409), .A2(n_226), .B(n_217), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_377), .B(n_16), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_390), .A2(n_226), .B1(n_17), .B2(n_241), .C(n_153), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_392), .A2(n_241), .B1(n_153), .B2(n_17), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_378), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_363), .B(n_241), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_381), .Y(n_443) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_405), .B(n_241), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_385), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_399), .B(n_241), .C(n_153), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_394), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_363), .A2(n_153), .B1(n_185), .B2(n_147), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_405), .A2(n_153), .B(n_19), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_371), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_401), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_399), .A2(n_153), .B1(n_159), .B2(n_22), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_401), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_370), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_382), .Y(n_455) );
AOI221x1_ASAP7_75t_L g456 ( .A1(n_420), .A2(n_376), .B1(n_379), .B2(n_408), .C(n_404), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_445), .A2(n_404), .B1(n_386), .B2(n_391), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_422), .A2(n_408), .B1(n_373), .B2(n_387), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_450), .B(n_373), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_443), .A2(n_387), .B1(n_391), .B2(n_386), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_416), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_418), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_421), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_417), .B(n_400), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_426), .A2(n_380), .B1(n_400), .B2(n_412), .C(n_388), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_454), .B(n_370), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_444), .A2(n_388), .B(n_382), .Y(n_467) );
INVxp33_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_434), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_415), .A2(n_412), .B1(n_396), .B2(n_393), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_455), .B(n_371), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_439), .Y(n_472) );
O2A1O1Ixp5_ASAP7_75t_L g473 ( .A1(n_424), .A2(n_374), .B(n_397), .C(n_389), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_440), .Y(n_474) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_421), .A2(n_410), .B1(n_397), .B2(n_389), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_447), .Y(n_476) );
O2A1O1Ixp5_ASAP7_75t_L g477 ( .A1(n_424), .A2(n_413), .B(n_414), .C(n_430), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_417), .A2(n_393), .B(n_396), .C(n_25), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_451), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_429), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_423), .A2(n_153), .B1(n_147), .B2(n_159), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_419), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_471), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_458), .A2(n_468), .B1(n_456), .B2(n_463), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_480), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_457), .A2(n_441), .B(n_431), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_457), .B(n_436), .Y(n_488) );
OAI21xp5_ASAP7_75t_SL g489 ( .A1(n_478), .A2(n_470), .B(n_465), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_477), .A2(n_446), .B(n_449), .C(n_442), .Y(n_490) );
AOI211x1_ASAP7_75t_SL g491 ( .A1(n_467), .A2(n_452), .B(n_435), .C(n_425), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_470), .A2(n_437), .B1(n_438), .B2(n_432), .C(n_448), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_464), .Y(n_493) );
OAI211xp5_ASAP7_75t_SL g494 ( .A1(n_481), .A2(n_427), .B(n_425), .C(n_433), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_460), .A2(n_442), .B1(n_159), .B2(n_26), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_483), .A2(n_159), .B1(n_20), .B2(n_27), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_464), .A2(n_18), .B1(n_31), .B2(n_32), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_461), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_475), .A2(n_147), .B1(n_36), .B2(n_43), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_459), .A2(n_147), .B1(n_45), .B2(n_47), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_484), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_489), .A2(n_473), .B(n_462), .Y(n_502) );
OAI21xp33_ASAP7_75t_L g503 ( .A1(n_485), .A2(n_466), .B(n_476), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_485), .A2(n_474), .B1(n_472), .B2(n_469), .C(n_479), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_498), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_493), .A2(n_482), .B(n_48), .C(n_51), .Y(n_506) );
OAI211xp5_ASAP7_75t_SL g507 ( .A1(n_491), .A2(n_35), .B(n_54), .C(n_55), .Y(n_507) );
OAI311xp33_ASAP7_75t_L g508 ( .A1(n_487), .A2(n_56), .A3(n_57), .B1(n_58), .C1(n_63), .Y(n_508) );
AOI222xp33_ASAP7_75t_L g509 ( .A1(n_488), .A2(n_147), .B1(n_66), .B2(n_68), .C1(n_69), .C2(n_72), .Y(n_509) );
NOR2x1p5_ASAP7_75t_L g510 ( .A(n_501), .B(n_486), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_507), .B(n_497), .C(n_492), .Y(n_511) );
NOR2x1p5_ASAP7_75t_L g512 ( .A(n_505), .B(n_490), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_502), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_504), .B(n_499), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_510), .B(n_500), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_514), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_512), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_515), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_515), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g520 ( .A1(n_518), .A2(n_513), .B1(n_517), .B2(n_516), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_520), .A2(n_518), .B1(n_511), .B2(n_519), .C(n_503), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_521), .A2(n_506), .B(n_509), .Y(n_522) );
OAI22xp33_ASAP7_75t_L g523 ( .A1(n_522), .A2(n_496), .B1(n_495), .B2(n_508), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_523), .A2(n_494), .B1(n_64), .B2(n_74), .Y(n_524) );
endmodule