module fake_jpeg_3123_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_7),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_56),
.Y(n_62)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_38),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_43),
.B1(n_41),
.B2(n_50),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_70),
.B1(n_59),
.B2(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_47),
.B1(n_40),
.B2(n_50),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_0),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_47),
.B1(n_40),
.B2(n_45),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_79),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_59),
.B1(n_42),
.B2(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_100),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_77),
.B1(n_4),
.B2(n_5),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_42),
.B1(n_1),
.B2(n_3),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_98),
.B1(n_0),
.B2(n_6),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_20),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_6),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_74),
.B(n_77),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_9),
.B(n_10),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_110),
.C(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_7),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_8),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_8),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_11),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_93),
.C(n_98),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_103),
.B1(n_127),
.B2(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_134),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_118),
.B(n_102),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_136),
.A2(n_120),
.B1(n_123),
.B2(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_131),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_119),
.C(n_126),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_143),
.C(n_144),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_133),
.B1(n_123),
.B2(n_137),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_114),
.B1(n_130),
.B2(n_13),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.C(n_15),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_111),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_111),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.C1(n_25),
.C2(n_27),
.Y(n_149)
);

AOI322xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_29),
.A3(n_30),
.B1(n_32),
.B2(n_33),
.C1(n_34),
.C2(n_35),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_14),
.B(n_148),
.Y(n_151)
);


endmodule