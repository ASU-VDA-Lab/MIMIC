module fake_netlist_6_2901_n_1219 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1219);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1219;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_1079;
wire n_341;
wire n_362;
wire n_1212;
wire n_828;
wire n_462;
wire n_671;
wire n_726;
wire n_607;
wire n_1033;
wire n_419;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1217;
wire n_751;
wire n_449;
wire n_749;
wire n_1208;
wire n_798;
wire n_1164;
wire n_509;
wire n_1209;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_1214;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_823;
wire n_557;
wire n_1132;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_1192;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_517;
wire n_718;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_1206;
wire n_621;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_923;
wire n_504;
wire n_1078;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_1015;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_1205;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_1216;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_1004;
wire n_953;
wire n_1094;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_1213;
wire n_638;
wire n_1181;
wire n_910;
wire n_1211;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_1215;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_492;
wire n_972;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_1041;
wire n_686;
wire n_796;
wire n_1195;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_731;
wire n_570;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_811;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_630;
wire n_958;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_1218;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_1198;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1146;
wire n_1141;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_550;
wire n_487;
wire n_1125;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1207;
wire n_1111;
wire n_511;
wire n_715;
wire n_467;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_1167;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_1153;
wire n_439;
wire n_518;
wire n_1210;
wire n_679;
wire n_1069;
wire n_1185;
wire n_612;
wire n_453;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_825;
wire n_636;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_434;
wire n_515;
wire n_983;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_736;
wire n_613;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_410;
wire n_398;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;

BUFx10_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_312),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_314),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_48),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_44),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_132),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_34),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_183),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_140),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_105),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_256),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_15),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_85),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_24),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_231),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_145),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_206),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_14),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_172),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_98),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_217),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_297),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_93),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_194),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_232),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_19),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_12),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_15),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_56),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_6),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_60),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_213),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_181),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_311),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_135),
.Y(n_353)
);

BUFx2_ASAP7_75t_SL g354 ( 
.A(n_293),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_158),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_171),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_100),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_199),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_185),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_262),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_69),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_198),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_125),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_66),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_267),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_218),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_76),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_196),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_0),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_316),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_290),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_146),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_5),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_62),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_219),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_167),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_168),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_77),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_236),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_144),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_113),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_123),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_226),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_156),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_137),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_46),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_280),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_225),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_243),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_306),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_67),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_114),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_253),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_223),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_273),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_11),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_307),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_192),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_107),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_242),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_265),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_63),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_108),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_96),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_64),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_275),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_16),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_1),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_304),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_186),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_189),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_6),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_119),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_294),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_264),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_133),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_12),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_30),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_188),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_215),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_261),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_224),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_278),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_155),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_251),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_55),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_86),
.Y(n_429)
);

BUFx8_ASAP7_75t_SL g430 ( 
.A(n_45),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_94),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_241),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_187),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_208),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_249),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_143),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_161),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_31),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_120),
.Y(n_439)
);

BUFx2_ASAP7_75t_SL g440 ( 
.A(n_173),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_303),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_233),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_51),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_17),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_22),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_33),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_301),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_266),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_295),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_175),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_43),
.Y(n_451)
);

BUFx5_ASAP7_75t_L g452 ( 
.A(n_82),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_50),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_263),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_170),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_229),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_220),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_23),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_7),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_216),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_37),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_197),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_26),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_90),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_152),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_260),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_147),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_210),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_287),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_202),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_97),
.Y(n_471)
);

BUFx2_ASAP7_75t_SL g472 ( 
.A(n_87),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_24),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_35),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_88),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_130),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_221),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_227),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_110),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_104),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_10),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_61),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_214),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_248),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_259),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_284),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_238),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_272),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_9),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_124),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_240),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_33),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_117),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_176),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_179),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_308),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_184),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_277),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_203),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_292),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_305),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_165),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_129),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_200),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_72),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_148),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_39),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_164),
.Y(n_508)
);

BUFx8_ASAP7_75t_SL g509 ( 
.A(n_247),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_78),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_41),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_222),
.Y(n_512)
);

INVxp33_ASAP7_75t_R g513 ( 
.A(n_115),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_35),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_257),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_174),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_296),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_178),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_38),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_28),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_149),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_212),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_3),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_250),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_57),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_302),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_157),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_328),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_338),
.B(n_0),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_433),
.B(n_499),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_343),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_338),
.B(n_442),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_385),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_330),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_369),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_391),
.B(n_1),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_385),
.Y(n_540)
);

BUFx12f_ASAP7_75t_L g541 ( 
.A(n_323),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_385),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_410),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_444),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_442),
.B(n_352),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_433),
.B(n_2),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_393),
.B(n_2),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_334),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_445),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_471),
.B(n_3),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_385),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_499),
.B(n_4),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_392),
.B(n_36),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_317),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_423),
.B(n_4),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_392),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_392),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_323),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_392),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_481),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_317),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_452),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_485),
.B(n_5),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_371),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_452),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_321),
.B(n_7),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_355),
.B(n_8),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_448),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_371),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_372),
.B(n_8),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_434),
.B(n_9),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_478),
.B(n_10),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_448),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_520),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_448),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_320),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_344),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_443),
.B(n_11),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_395),
.B(n_13),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_405),
.B(n_13),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_500),
.B(n_14),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_40),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_345),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_16),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_455),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_519),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_455),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_322),
.B(n_17),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_347),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_465),
.B(n_18),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_519),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_452),
.B(n_18),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_467),
.B(n_19),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_519),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_519),
.Y(n_597)
);

AND2x4_ASAP7_75t_SL g598 ( 
.A(n_498),
.B(n_42),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_498),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_324),
.B(n_20),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_329),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_333),
.B(n_20),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g604 ( 
.A(n_501),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_373),
.B(n_397),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_335),
.Y(n_606)
);

NOR2x1_ASAP7_75t_L g607 ( 
.A(n_337),
.B(n_47),
.Y(n_607)
);

XNOR2x1_ASAP7_75t_L g608 ( 
.A(n_409),
.B(n_21),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_341),
.B(n_342),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_332),
.B(n_21),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_414),
.B(n_22),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_348),
.B(n_401),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_349),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_350),
.B(n_23),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_420),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_430),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_509),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_356),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_357),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_359),
.B(n_25),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_318),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_429),
.B(n_25),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_319),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_362),
.B(n_364),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_325),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_446),
.B(n_26),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_365),
.Y(n_627)
);

NOR2x1_ASAP7_75t_L g628 ( 
.A(n_367),
.B(n_49),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_368),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_376),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_354),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_435),
.B(n_27),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_462),
.B(n_27),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_378),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_380),
.B(n_28),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_327),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_459),
.B(n_463),
.Y(n_637)
);

BUFx12f_ASAP7_75t_L g638 ( 
.A(n_473),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_382),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_331),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_336),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_474),
.Y(n_642)
);

AO22x2_ASAP7_75t_L g643 ( 
.A1(n_534),
.A2(n_472),
.B1(n_440),
.B2(n_389),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_605),
.B(n_339),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_612),
.A2(n_351),
.B1(n_358),
.B2(n_326),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_579),
.A2(n_379),
.B1(n_384),
.B2(n_363),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_592),
.A2(n_422),
.B1(n_457),
.B2(n_412),
.Y(n_647)
);

OA22x2_ASAP7_75t_L g648 ( 
.A1(n_564),
.A2(n_578),
.B1(n_585),
.B2(n_548),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_551),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_637),
.B(n_340),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_595),
.A2(n_491),
.B1(n_510),
.B2(n_461),
.Y(n_651)
);

AO22x2_ASAP7_75t_L g652 ( 
.A1(n_546),
.A2(n_400),
.B1(n_402),
.B2(n_387),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_R g653 ( 
.A1(n_530),
.A2(n_458),
.B1(n_438),
.B2(n_513),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_551),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_556),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_539),
.A2(n_514),
.B1(n_523),
.B2(n_489),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_615),
.B(n_642),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_556),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_576),
.Y(n_659)
);

OA22x2_ASAP7_75t_L g660 ( 
.A1(n_529),
.A2(n_408),
.B1(n_417),
.B2(n_403),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_SL g661 ( 
.A1(n_611),
.A2(n_421),
.B1(n_427),
.B2(n_418),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_545),
.A2(n_516),
.B1(n_353),
.B2(n_360),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_610),
.A2(n_346),
.B1(n_361),
.B2(n_525),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_529),
.B(n_366),
.Y(n_664)
);

OAI22x1_ASAP7_75t_L g665 ( 
.A1(n_561),
.A2(n_527),
.B1(n_526),
.B2(n_524),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_631),
.B(n_439),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_576),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_633),
.A2(n_522),
.B1(n_521),
.B2(n_518),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_588),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_588),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_537),
.B(n_370),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_638),
.A2(n_454),
.B1(n_515),
.B2(n_512),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_L g673 ( 
.A1(n_622),
.A2(n_632),
.B1(n_599),
.B2(n_602),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_537),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_591),
.B(n_374),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_SL g676 ( 
.A(n_555),
.B(n_375),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_597),
.Y(n_677)
);

AO22x2_ASAP7_75t_L g678 ( 
.A1(n_546),
.A2(n_493),
.B1(n_507),
.B2(n_505),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_626),
.A2(n_451),
.B1(n_508),
.B2(n_506),
.Y(n_679)
);

AO22x2_ASAP7_75t_L g680 ( 
.A1(n_552),
.A2(n_480),
.B1(n_497),
.B2(n_495),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_602),
.A2(n_517),
.B1(n_456),
.B2(n_470),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_SL g682 ( 
.A1(n_550),
.A2(n_475),
.B1(n_486),
.B2(n_502),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_541),
.B(n_29),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_591),
.B(n_29),
.Y(n_685)
);

AO22x2_ASAP7_75t_L g686 ( 
.A1(n_552),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_559),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_568),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_547),
.A2(n_436),
.B1(n_503),
.B2(n_496),
.Y(n_689)
);

AO22x2_ASAP7_75t_L g690 ( 
.A1(n_608),
.A2(n_32),
.B1(n_34),
.B2(n_504),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_604),
.A2(n_431),
.B1(n_490),
.B2(n_488),
.Y(n_691)
);

AO22x2_ASAP7_75t_L g692 ( 
.A1(n_572),
.A2(n_494),
.B1(n_487),
.B2(n_484),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_563),
.A2(n_483),
.B1(n_482),
.B2(n_479),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_634),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_631),
.B(n_377),
.Y(n_695)
);

OA22x2_ASAP7_75t_L g696 ( 
.A1(n_575),
.A2(n_477),
.B1(n_476),
.B2(n_469),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_558),
.A2(n_468),
.B1(n_466),
.B2(n_464),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_SL g698 ( 
.A1(n_594),
.A2(n_460),
.B1(n_453),
.B2(n_450),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_SL g699 ( 
.A1(n_635),
.A2(n_449),
.B1(n_447),
.B2(n_441),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_574),
.Y(n_700)
);

AO22x2_ASAP7_75t_L g701 ( 
.A1(n_572),
.A2(n_437),
.B1(n_432),
.B2(n_428),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_616),
.B(n_381),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_623),
.B(n_383),
.Y(n_703)
);

AO22x2_ASAP7_75t_L g704 ( 
.A1(n_573),
.A2(n_426),
.B1(n_425),
.B2(n_424),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_554),
.B(n_386),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_573),
.A2(n_416),
.B1(n_415),
.B2(n_413),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_533),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_535),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_625),
.B(n_388),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_569),
.A2(n_411),
.B1(n_407),
.B2(n_406),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_624),
.A2(n_404),
.B1(n_399),
.B2(n_398),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_636),
.B(n_390),
.Y(n_712)
);

AOI22x1_ASAP7_75t_L g713 ( 
.A1(n_581),
.A2(n_396),
.B1(n_394),
.B2(n_54),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_587),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_59),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_589),
.B(n_65),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_577),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_562),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_565),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_606),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_SL g722 ( 
.A1(n_614),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_631),
.B(n_73),
.Y(n_723)
);

XNOR2xp5_ASAP7_75t_L g724 ( 
.A(n_598),
.B(n_315),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_531),
.B(n_74),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_620),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_639),
.Y(n_727)
);

AND2x2_ASAP7_75t_SL g728 ( 
.A(n_581),
.B(n_582),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_R g729 ( 
.A1(n_532),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_SL g730 ( 
.A(n_582),
.B(n_89),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_531),
.B(n_91),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_590),
.A2(n_92),
.B1(n_95),
.B2(n_99),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_725),
.B(n_609),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_649),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_717),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_645),
.Y(n_736)
);

XOR2x2_ASAP7_75t_L g737 ( 
.A(n_646),
.B(n_566),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_662),
.B(n_621),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_727),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_707),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_708),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_705),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_657),
.B(n_640),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_718),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_664),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_719),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_720),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_654),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_655),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_663),
.B(n_617),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_668),
.B(n_617),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_667),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_728),
.A2(n_609),
.B(n_600),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_677),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_684),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_659),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_689),
.B(n_617),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_647),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_658),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_731),
.A2(n_650),
.B(n_644),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_659),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_669),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_670),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_695),
.B(n_536),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_651),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_687),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_721),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_673),
.B(n_553),
.Y(n_768)
);

XNOR2x2_ASAP7_75t_L g769 ( 
.A(n_690),
.B(n_567),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_688),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_671),
.Y(n_771)
);

INVxp33_ASAP7_75t_L g772 ( 
.A(n_674),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_700),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_694),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_706),
.B(n_590),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_666),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_660),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_675),
.B(n_601),
.Y(n_778)
);

CKINVDCx16_ASAP7_75t_R g779 ( 
.A(n_691),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_685),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_703),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_679),
.B(n_600),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_709),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_712),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_713),
.Y(n_785)
);

INVxp33_ASAP7_75t_SL g786 ( 
.A(n_699),
.Y(n_786)
);

XNOR2xp5_ASAP7_75t_L g787 ( 
.A(n_724),
.B(n_603),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_696),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_665),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_652),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_656),
.B(n_603),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_652),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_715),
.Y(n_793)
);

INVx4_ASAP7_75t_SL g794 ( 
.A(n_683),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_678),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_686),
.B(n_586),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_678),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_680),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_680),
.Y(n_799)
);

XNOR2x2_ASAP7_75t_L g800 ( 
.A(n_690),
.B(n_571),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_676),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_710),
.B(n_583),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_698),
.B(n_536),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_732),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_723),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_730),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_643),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_643),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_L g810 ( 
.A(n_714),
.B(n_536),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_648),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_702),
.B(n_601),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_661),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_711),
.B(n_540),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_693),
.B(n_672),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_686),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_778),
.B(n_692),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_796),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_770),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_740),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_735),
.Y(n_821)
);

AND2x2_ASAP7_75t_SL g822 ( 
.A(n_791),
.B(n_586),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_793),
.B(n_692),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_793),
.B(n_753),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_806),
.B(n_701),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_770),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_782),
.B(n_701),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_739),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_770),
.Y(n_829)
);

BUFx12f_ASAP7_75t_SL g830 ( 
.A(n_796),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_771),
.B(n_745),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_776),
.B(n_704),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_772),
.B(n_704),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_767),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_774),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_767),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_780),
.B(n_702),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_742),
.B(n_697),
.Y(n_838)
);

AND2x2_ASAP7_75t_SL g839 ( 
.A(n_815),
.B(n_729),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_788),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_736),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_733),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_766),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_773),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_733),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_781),
.B(n_716),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_783),
.B(n_784),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_741),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_743),
.B(n_682),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_775),
.B(n_553),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_744),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_777),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_785),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_812),
.B(n_683),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_746),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_760),
.B(n_532),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_767),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_756),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_786),
.B(n_722),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_738),
.B(n_538),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_807),
.B(n_553),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_747),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_734),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_748),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_768),
.B(n_726),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_811),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_787),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_749),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_805),
.B(n_584),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_796),
.B(n_538),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_752),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_813),
.B(n_584),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_737),
.B(n_543),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_754),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_789),
.B(n_584),
.Y(n_875)
);

BUFx4f_ASAP7_75t_L g876 ( 
.A(n_801),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_790),
.B(n_607),
.Y(n_877)
);

CKINVDCx12_ASAP7_75t_R g878 ( 
.A(n_761),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_810),
.B(n_628),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_757),
.B(n_629),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_755),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_759),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_762),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_792),
.B(n_681),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_808),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_795),
.B(n_629),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_763),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_801),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_797),
.B(n_606),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_798),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_799),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_809),
.B(n_543),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_801),
.B(n_544),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_816),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_750),
.B(n_613),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_804),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_814),
.Y(n_897)
);

AND2x6_ASAP7_75t_L g898 ( 
.A(n_853),
.B(n_894),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_834),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_SL g900 ( 
.A(n_839),
.B(n_779),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_860),
.B(n_751),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_842),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_856),
.B(n_810),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_853),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_822),
.B(n_764),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_820),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_834),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_830),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_820),
.Y(n_909)
);

BUFx6f_ASAP7_75t_SL g910 ( 
.A(n_888),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_873),
.B(n_769),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_831),
.B(n_794),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_843),
.B(n_794),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_843),
.B(n_802),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_822),
.B(n_764),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_842),
.B(n_544),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_842),
.B(n_549),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_848),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_867),
.B(n_758),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_827),
.B(n_800),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_847),
.B(n_765),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_888),
.B(n_549),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_845),
.B(n_888),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_848),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_841),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_855),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_893),
.B(n_560),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_853),
.B(n_613),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_866),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_845),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_841),
.B(n_560),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_894),
.B(n_618),
.Y(n_932)
);

BUFx12f_ASAP7_75t_L g933 ( 
.A(n_818),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_889),
.B(n_570),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_855),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_891),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_830),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_876),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_894),
.B(n_618),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_854),
.B(n_570),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_896),
.B(n_653),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_876),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_866),
.Y(n_943)
);

AND2x6_ASAP7_75t_L g944 ( 
.A(n_824),
.B(n_528),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_870),
.B(n_528),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_896),
.B(n_619),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_839),
.B(n_619),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_891),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_838),
.B(n_627),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_845),
.Y(n_950)
);

BUFx5_ASAP7_75t_L g951 ( 
.A(n_857),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_871),
.Y(n_952)
);

AND2x6_ASAP7_75t_L g953 ( 
.A(n_850),
.B(n_627),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_880),
.B(n_630),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_896),
.B(n_630),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_883),
.B(n_540),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_829),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_923),
.Y(n_958)
);

CKINVDCx6p67_ASAP7_75t_R g959 ( 
.A(n_938),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_933),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_936),
.Y(n_961)
);

INVx5_ASAP7_75t_L g962 ( 
.A(n_898),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_957),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_931),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_923),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_901),
.A2(n_859),
.B1(n_849),
.B2(n_896),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_904),
.A2(n_868),
.B(n_883),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_936),
.Y(n_968)
);

INVx8_ASAP7_75t_L g969 ( 
.A(n_910),
.Y(n_969)
);

BUFx4f_ASAP7_75t_SL g970 ( 
.A(n_913),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_899),
.Y(n_971)
);

BUFx8_ASAP7_75t_SL g972 ( 
.A(n_925),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_948),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_921),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_948),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_929),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_899),
.Y(n_977)
);

BUFx24_ASAP7_75t_L g978 ( 
.A(n_914),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_913),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_916),
.B(n_821),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_908),
.Y(n_981)
);

INVx5_ASAP7_75t_SL g982 ( 
.A(n_940),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_940),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_942),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_907),
.Y(n_985)
);

INVx8_ASAP7_75t_L g986 ( 
.A(n_910),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_949),
.B(n_817),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_916),
.Y(n_988)
);

CKINVDCx6p67_ASAP7_75t_R g989 ( 
.A(n_941),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_904),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_927),
.B(n_833),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_943),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_917),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_951),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_907),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_903),
.B(n_902),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_902),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_914),
.Y(n_998)
);

CKINVDCx11_ASAP7_75t_R g999 ( 
.A(n_941),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_917),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_898),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_947),
.A2(n_897),
.B1(n_823),
.B2(n_825),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_930),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_961),
.Y(n_1004)
);

INVx6_ASAP7_75t_L g1005 ( 
.A(n_969),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_961),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_SL g1007 ( 
.A1(n_974),
.A2(n_900),
.B1(n_911),
.B2(n_920),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_968),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_991),
.A2(n_865),
.B1(n_900),
.B2(n_832),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_962),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_980),
.A2(n_865),
.B1(n_840),
.B2(n_919),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_980),
.A2(n_993),
.B1(n_1000),
.B2(n_988),
.Y(n_1012)
);

CKINVDCx11_ASAP7_75t_R g1013 ( 
.A(n_984),
.Y(n_1013)
);

INVx8_ASAP7_75t_L g1014 ( 
.A(n_969),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_966),
.B(n_945),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_969),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_973),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_964),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_962),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_SL g1020 ( 
.A1(n_994),
.A2(n_826),
.B(n_819),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_980),
.A2(n_840),
.B1(n_944),
.B2(n_846),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_999),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_975),
.Y(n_1023)
);

INVx6_ASAP7_75t_SL g1024 ( 
.A(n_978),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_987),
.B(n_912),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_1002),
.A2(n_944),
.B1(n_935),
.B2(n_924),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_976),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_990),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_SL g1029 ( 
.A1(n_998),
.A2(n_837),
.B(n_884),
.Y(n_1029)
);

INVx6_ASAP7_75t_L g1030 ( 
.A(n_986),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_990),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_997),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_996),
.A2(n_944),
.B1(n_909),
.B2(n_906),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_976),
.Y(n_1034)
);

CKINVDCx11_ASAP7_75t_R g1035 ( 
.A(n_984),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_SL g1036 ( 
.A1(n_978),
.A2(n_884),
.B1(n_892),
.B2(n_915),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_SL g1037 ( 
.A(n_959),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_997),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_992),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_992),
.Y(n_1040)
);

CKINVDCx11_ASAP7_75t_R g1041 ( 
.A(n_999),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_963),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_1007),
.A2(n_895),
.B(n_954),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_1036),
.A2(n_989),
.B1(n_944),
.B2(n_983),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_SL g1045 ( 
.A1(n_1015),
.A2(n_982),
.B1(n_986),
.B2(n_905),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1007),
.B(n_852),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_1037),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_SL g1048 ( 
.A1(n_1029),
.A2(n_879),
.B(n_937),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1025),
.B(n_852),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_SL g1050 ( 
.A1(n_1036),
.A2(n_879),
.B(n_828),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_1013),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_1022),
.A2(n_982),
.B1(n_986),
.B2(n_962),
.Y(n_1052)
);

OAI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_1009),
.A2(n_1011),
.B(n_1021),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1027),
.B(n_934),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_SL g1055 ( 
.A1(n_1009),
.A2(n_877),
.B(n_835),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1024),
.A2(n_996),
.B1(n_882),
.B2(n_946),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1018),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1024),
.A2(n_882),
.B1(n_955),
.B2(n_946),
.Y(n_1058)
);

OAI222xp33_ASAP7_75t_L g1059 ( 
.A1(n_1042),
.A2(n_955),
.B1(n_963),
.B2(n_885),
.C1(n_928),
.C2(n_952),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1008),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_1037),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1004),
.Y(n_1062)
);

BUFx12f_ASAP7_75t_L g1063 ( 
.A(n_1035),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_1016),
.Y(n_1064)
);

AOI222xp33_ASAP7_75t_L g1065 ( 
.A1(n_1034),
.A2(n_1041),
.B1(n_982),
.B2(n_1027),
.C1(n_1039),
.C2(n_1040),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1012),
.A2(n_882),
.B1(n_844),
.B2(n_869),
.Y(n_1066)
);

OAI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1016),
.A2(n_922),
.B1(n_981),
.B2(n_958),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_SL g1068 ( 
.A(n_1016),
.Y(n_1068)
);

OAI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1005),
.A2(n_981),
.B1(n_965),
.B2(n_958),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1026),
.A2(n_882),
.B1(n_883),
.B2(n_926),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1026),
.A2(n_918),
.B1(n_851),
.B2(n_862),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1017),
.A2(n_994),
.B1(n_1001),
.B2(n_962),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_SL g1073 ( 
.A(n_1010),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1023),
.A2(n_1001),
.B1(n_886),
.B2(n_890),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1033),
.A2(n_872),
.B1(n_887),
.B2(n_881),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_1014),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1033),
.A2(n_874),
.B1(n_930),
.B2(n_950),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1028),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1032),
.A2(n_950),
.B1(n_871),
.B2(n_877),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1038),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1057),
.B(n_1031),
.Y(n_1081)
);

AOI222xp33_ASAP7_75t_L g1082 ( 
.A1(n_1053),
.A2(n_864),
.B1(n_863),
.B2(n_875),
.C1(n_858),
.C2(n_960),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1060),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1046),
.A2(n_1006),
.B1(n_1030),
.B2(n_1005),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1078),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1044),
.A2(n_953),
.B1(n_868),
.B2(n_965),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1062),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_1043),
.A2(n_939),
.B(n_932),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1058),
.A2(n_1005),
.B1(n_1030),
.B2(n_1001),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1045),
.A2(n_953),
.B1(n_868),
.B2(n_857),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1065),
.A2(n_953),
.B1(n_1003),
.B2(n_858),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1048),
.A2(n_1030),
.B1(n_1001),
.B2(n_1014),
.Y(n_1092)
);

OAI222xp33_ASAP7_75t_L g1093 ( 
.A1(n_1056),
.A2(n_928),
.B1(n_1010),
.B2(n_1019),
.C1(n_1003),
.C2(n_861),
.Y(n_1093)
);

OAI222xp33_ASAP7_75t_L g1094 ( 
.A1(n_1054),
.A2(n_1052),
.B1(n_1074),
.B2(n_1069),
.C1(n_1067),
.C2(n_1071),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1066),
.A2(n_1014),
.B1(n_970),
.B2(n_960),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1050),
.A2(n_970),
.B1(n_979),
.B2(n_1019),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_SL g1097 ( 
.A1(n_1065),
.A2(n_1055),
.B(n_1059),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1049),
.A2(n_953),
.B1(n_979),
.B2(n_878),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1063),
.A2(n_972),
.B1(n_898),
.B2(n_951),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1074),
.A2(n_972),
.B1(n_898),
.B2(n_951),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1080),
.B(n_971),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1051),
.A2(n_878),
.B1(n_826),
.B2(n_819),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1072),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1075),
.B(n_977),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1073),
.B(n_1079),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1070),
.A2(n_829),
.B1(n_826),
.B2(n_819),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1072),
.A2(n_829),
.B1(n_951),
.B2(n_834),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1064),
.B(n_971),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1068),
.A2(n_1077),
.B1(n_1061),
.B2(n_1047),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1068),
.A2(n_829),
.B1(n_951),
.B2(n_834),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1047),
.A2(n_836),
.B1(n_971),
.B2(n_985),
.Y(n_1111)
);

OAI222xp33_ASAP7_75t_L g1112 ( 
.A1(n_1061),
.A2(n_995),
.B1(n_985),
.B2(n_977),
.C1(n_836),
.C2(n_956),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1064),
.B(n_971),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_SL g1114 ( 
.A1(n_1064),
.A2(n_995),
.B1(n_967),
.B2(n_836),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1076),
.A2(n_967),
.B1(n_596),
.B2(n_593),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1059),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1083),
.B(n_101),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1116),
.B(n_1020),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1085),
.B(n_540),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1092),
.A2(n_596),
.B1(n_593),
.B2(n_557),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1101),
.B(n_102),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1097),
.A2(n_103),
.B(n_106),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_1082),
.B(n_596),
.C(n_593),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1096),
.A2(n_557),
.B1(n_542),
.B2(n_112),
.Y(n_1124)
);

AOI211x1_ASAP7_75t_L g1125 ( 
.A1(n_1081),
.A2(n_109),
.B(n_111),
.C(n_116),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1087),
.B(n_118),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1088),
.A2(n_557),
.B1(n_542),
.B2(n_126),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1094),
.A2(n_542),
.B1(n_122),
.B2(n_127),
.C(n_128),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1084),
.B(n_1103),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_SL g1130 ( 
.A1(n_1099),
.A2(n_121),
.B(n_131),
.Y(n_1130)
);

NAND3xp33_ASAP7_75t_L g1131 ( 
.A(n_1084),
.B(n_1098),
.C(n_1091),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1104),
.B(n_134),
.Y(n_1132)
);

NAND4xp25_ASAP7_75t_L g1133 ( 
.A(n_1102),
.B(n_1099),
.C(n_1109),
.D(n_1100),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1095),
.A2(n_136),
.B(n_138),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1105),
.B(n_139),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1100),
.B(n_141),
.C(n_142),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1108),
.B(n_150),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1113),
.B(n_151),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1089),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1086),
.A2(n_153),
.B1(n_154),
.B2(n_159),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1107),
.B(n_160),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1119),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_L g1143 ( 
.A(n_1122),
.B(n_1093),
.C(n_1112),
.Y(n_1143)
);

AOI211xp5_ASAP7_75t_L g1144 ( 
.A1(n_1128),
.A2(n_1090),
.B(n_163),
.C(n_166),
.Y(n_1144)
);

NAND4xp75_ASAP7_75t_L g1145 ( 
.A(n_1125),
.B(n_1110),
.C(n_1114),
.D(n_1111),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_1119),
.B(n_1115),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1129),
.B(n_1115),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1139),
.B(n_1106),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1121),
.B(n_162),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1118),
.B(n_169),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1138),
.B(n_1118),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1117),
.B(n_177),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_L g1153 ( 
.A(n_1133),
.B(n_182),
.Y(n_1153)
);

NAND4xp75_ASAP7_75t_SL g1154 ( 
.A(n_1147),
.B(n_1130),
.C(n_1134),
.D(n_1123),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_1135),
.C(n_1131),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1142),
.Y(n_1156)
);

NAND4xp75_ASAP7_75t_SL g1157 ( 
.A(n_1153),
.B(n_1136),
.C(n_1124),
.D(n_1127),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1146),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1151),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_L g1160 ( 
.A(n_1150),
.B(n_1132),
.C(n_1137),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1148),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1143),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1145),
.Y(n_1163)
);

CKINVDCx14_ASAP7_75t_R g1164 ( 
.A(n_1163),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1158),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1156),
.Y(n_1166)
);

OA22x2_ASAP7_75t_SL g1167 ( 
.A1(n_1162),
.A2(n_1144),
.B1(n_1120),
.B2(n_1152),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1161),
.B(n_1149),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1159),
.B(n_1126),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1155),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1164),
.B(n_1160),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1166),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_1168),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1168),
.B(n_1141),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1165),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1169),
.Y(n_1176)
);

AOI22x1_ASAP7_75t_L g1177 ( 
.A1(n_1170),
.A2(n_1157),
.B1(n_1154),
.B2(n_1144),
.Y(n_1177)
);

AO22x1_ASAP7_75t_L g1178 ( 
.A1(n_1167),
.A2(n_1154),
.B1(n_1157),
.B2(n_1141),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1165),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1166),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1173),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1172),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1180),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1174),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1175),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1179),
.Y(n_1186)
);

AOI22x1_ASAP7_75t_L g1187 ( 
.A1(n_1182),
.A2(n_1178),
.B1(n_1177),
.B2(n_1176),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1182),
.Y(n_1188)
);

OAI322xp33_ASAP7_75t_L g1189 ( 
.A1(n_1183),
.A2(n_1177),
.A3(n_1171),
.B1(n_1140),
.B2(n_195),
.C1(n_201),
.C2(n_204),
.Y(n_1189)
);

NAND4xp75_ASAP7_75t_L g1190 ( 
.A(n_1181),
.B(n_190),
.C(n_191),
.D(n_193),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1186),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1184),
.A2(n_205),
.B1(n_207),
.B2(n_209),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1188),
.A2(n_1185),
.B1(n_228),
.B2(n_230),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1191),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_1192),
.A2(n_211),
.B(n_234),
.C(n_235),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1187),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1194),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1196),
.Y(n_1198)
);

AO22x2_ASAP7_75t_SL g1199 ( 
.A1(n_1193),
.A2(n_1190),
.B1(n_1189),
.B2(n_245),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1198),
.A2(n_1195),
.B1(n_244),
.B2(n_246),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1197),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1197),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1201),
.B(n_1199),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1202),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1203),
.A2(n_1200),
.B1(n_1204),
.B2(n_254),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1205),
.A2(n_310),
.B1(n_252),
.B2(n_255),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1205),
.B(n_237),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1206),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1207),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1208),
.A2(n_1209),
.B1(n_268),
.B2(n_269),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1208),
.A2(n_258),
.B1(n_270),
.B2(n_271),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1208),
.A2(n_274),
.B1(n_276),
.B2(n_279),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1210),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1213),
.A2(n_1212),
.B1(n_1211),
.B2(n_283),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1213),
.A2(n_281),
.B1(n_282),
.B2(n_285),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1215),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1214),
.Y(n_1217)
);

AOI221xp5_ASAP7_75t_L g1218 ( 
.A1(n_1216),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_1218)
);

AOI211xp5_ASAP7_75t_L g1219 ( 
.A1(n_1218),
.A2(n_1217),
.B(n_298),
.C(n_299),
.Y(n_1219)
);


endmodule