module fake_netlist_5_1359_n_473 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_473);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_473;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_451;
wire n_408;
wire n_376;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_467;
wire n_423;
wire n_284;
wire n_245;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_368;
wire n_247;
wire n_314;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_275;
wire n_252;
wire n_295;
wire n_330;
wire n_373;
wire n_307;
wire n_439;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_191;
wire n_171;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_470;
wire n_325;
wire n_449;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_457;
wire n_297;
wire n_225;
wire n_377;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_422;
wire n_415;
wire n_355;
wire n_336;
wire n_337;
wire n_430;
wire n_313;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_328;
wire n_214;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_165;
wire n_468;
wire n_213;
wire n_342;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_461;
wire n_333;
wire n_309;
wire n_462;
wire n_322;
wire n_258;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_463;
wire n_239;
wire n_466;
wire n_420;
wire n_310;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_441;
wire n_450;
wire n_312;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_410;
wire n_269;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_58),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_31),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_9),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_96),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_51),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_20),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_30),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_26),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_119),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_75),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_87),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_70),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_33),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_16),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_73),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_25),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_56),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_28),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_72),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_39),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_17),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_18),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_32),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_153),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_8),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_55),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_49),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_144),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_4),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_15),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_52),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_77),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_5),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_62),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_67),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_71),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_125),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_12),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_81),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_95),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_19),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_24),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_46),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_131),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_54),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_29),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_50),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_23),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_64),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_84),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_146),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_6),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_105),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_40),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_143),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_139),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_89),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_123),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_129),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_79),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_130),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_66),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_22),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_42),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_69),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_63),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_11),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_100),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_134),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_149),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_114),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_78),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_13),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_152),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_138),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_140),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_97),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_147),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_65),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_133),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_47),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_44),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_151),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_0),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_34),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_74),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_126),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_98),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_172),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_189),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_158),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_161),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_164),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_189),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_159),
.B(n_14),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_209),
.A2(n_21),
.B1(n_27),
.B2(n_35),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_189),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_162),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_167),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_170),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_166),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_266),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_174),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_176),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_186),
.B(n_59),
.Y(n_308)
);

XOR2x2_ASAP7_75t_SL g309 ( 
.A(n_177),
.B(n_60),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_184),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_179),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_193),
.A2(n_76),
.B1(n_80),
.B2(n_82),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_165),
.B(n_242),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_180),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_276),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_185),
.B(n_90),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_168),
.B(n_92),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_198),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_187),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_190),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_192),
.B(n_93),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_194),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_199),
.A2(n_94),
.B1(n_102),
.B2(n_103),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_196),
.B(n_104),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_201),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_202),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_243),
.B(n_109),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_203),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_204),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_205),
.A2(n_113),
.B(n_115),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_206),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_232),
.A2(n_256),
.B1(n_244),
.B2(n_265),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_207),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_211),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_216),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_240),
.B(n_118),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_218),
.Y(n_341)
);

OAI221xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_188),
.B1(n_173),
.B2(n_215),
.C(n_235),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_307),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_264),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_219),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_317),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_221),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

AO22x2_ASAP7_75t_L g354 ( 
.A1(n_309),
.A2(n_231),
.B1(n_281),
.B2(n_279),
.Y(n_354)
);

CKINVDCx11_ASAP7_75t_R g355 ( 
.A(n_310),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_320),
.Y(n_359)
);

OAI221xp5_ASAP7_75t_L g360 ( 
.A1(n_283),
.A2(n_260),
.B1(n_259),
.B2(n_257),
.C(n_253),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_258),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_288),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_285),
.B(n_175),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_241),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_169),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_319),
.B(n_213),
.Y(n_372)
);

OAI221xp5_ASAP7_75t_L g373 ( 
.A1(n_284),
.A2(n_208),
.B1(n_234),
.B2(n_226),
.C(n_237),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g375 ( 
.A1(n_308),
.A2(n_318),
.B1(n_340),
.B2(n_255),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g376 ( 
.A1(n_287),
.A2(n_251),
.B1(n_277),
.B2(n_275),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_296),
.B(n_225),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_249),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_298),
.Y(n_379)
);

OAI21x1_ASAP7_75t_L g380 ( 
.A1(n_352),
.A2(n_333),
.B(n_304),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_368),
.B(n_315),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_300),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_327),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_369),
.B(n_247),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_344),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_339),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_330),
.B1(n_337),
.B2(n_334),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_355),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_343),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_362),
.A2(n_314),
.B(n_329),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_316),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_321),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_305),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_301),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_359),
.Y(n_397)
);

AND3x1_ASAP7_75t_SL g398 ( 
.A(n_342),
.B(n_229),
.C(n_269),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_330),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_354),
.A2(n_217),
.B1(n_282),
.B2(n_212),
.Y(n_400)
);

NAND3xp33_ASAP7_75t_SL g401 ( 
.A(n_360),
.B(n_228),
.C(n_222),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_330),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_372),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_367),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_373),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_364),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_371),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_405),
.A2(n_345),
.B(n_377),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g412 ( 
.A1(n_380),
.A2(n_238),
.B(n_263),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_351),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_403),
.Y(n_415)
);

INVx3_ASAP7_75t_SL g416 ( 
.A(n_397),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_404),
.Y(n_417)
);

AOI211xp5_ASAP7_75t_L g418 ( 
.A1(n_400),
.A2(n_381),
.B(n_393),
.C(n_382),
.Y(n_418)
);

O2A1O1Ixp5_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_181),
.B(n_178),
.C(n_236),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_391),
.Y(n_420)
);

NOR2x2_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_325),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_370),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_392),
.B(n_214),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_395),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_376),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_419),
.A2(n_396),
.B(n_268),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_406),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_353),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_SL g431 ( 
.A1(n_420),
.A2(n_401),
.B(n_239),
.C(n_246),
.Y(n_431)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_408),
.A2(n_230),
.B(n_252),
.C(n_274),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_416),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_424),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_415),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_417),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_425),
.Y(n_437)
);

CKINVDCx11_ASAP7_75t_R g438 ( 
.A(n_433),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_430),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_435),
.Y(n_440)
);

A2O1A1Ixp33_ASAP7_75t_L g441 ( 
.A1(n_434),
.A2(n_411),
.B(n_424),
.C(n_423),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_430),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

AO21x2_ASAP7_75t_L g445 ( 
.A1(n_441),
.A2(n_431),
.B(n_432),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_437),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_442),
.A2(n_426),
.B1(n_290),
.B2(n_303),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_443),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_413),
.C(n_338),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_446),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_376),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_438),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_444),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_453),
.A2(n_312),
.B1(n_448),
.B2(n_450),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_451),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_456),
.B(n_454),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_455),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_456),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_456),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_459),
.B(n_452),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_461),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_457),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_463),
.A2(n_389),
.B1(n_273),
.B2(n_270),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_462),
.Y(n_466)
);

AOI222xp33_ASAP7_75t_L g467 ( 
.A1(n_465),
.A2(n_464),
.B1(n_224),
.B2(n_227),
.C1(n_248),
.C2(n_261),
.Y(n_467)
);

NAND4xp25_ASAP7_75t_L g468 ( 
.A(n_466),
.B(n_262),
.C(n_254),
.D(n_223),
.Y(n_468)
);

AOI211xp5_ASAP7_75t_L g469 ( 
.A1(n_468),
.A2(n_267),
.B(n_421),
.C(n_197),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_467),
.A2(n_191),
.B1(n_195),
.B2(n_182),
.Y(n_470)
);

OAI322xp33_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_338),
.A3(n_356),
.B1(n_398),
.B2(n_210),
.C1(n_280),
.C2(n_220),
.Y(n_471)
);

AOI21xp33_ASAP7_75t_L g472 ( 
.A1(n_471),
.A2(n_469),
.B(n_445),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_157),
.B1(n_428),
.B2(n_412),
.Y(n_473)
);


endmodule