module real_jpeg_14157_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_132)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_5),
.A2(n_74),
.B(n_77),
.C(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_71),
.B1(n_74),
.B2(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_5),
.B(n_82),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_104),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_5),
.A2(n_24),
.B1(n_36),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_5),
.B(n_110),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_71),
.B1(n_74),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_115),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_115),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_115),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_9),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_70),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_70),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_12),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_12),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_13),
.A2(n_65),
.B1(n_71),
.B2(n_74),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_65),
.Y(n_153)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_15),
.A2(n_71),
.B1(n_74),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_81),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_81),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_142),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_117),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_20),
.B(n_117),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_95),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_21),
.B(n_83),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_22),
.B(n_55),
.C(n_68),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_23),
.B(n_39),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_24),
.A2(n_36),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_24),
.A2(n_36),
.B1(n_211),
.B2(n_219),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_24),
.A2(n_86),
.B(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_25),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_25),
.A2(n_30),
.B1(n_32),
.B2(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_25),
.A2(n_35),
.B(n_87),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_25),
.A2(n_30),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_26),
.B(n_41),
.C(n_104),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_26),
.B(n_217),
.Y(n_216)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_36),
.A2(n_88),
.B(n_101),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_36),
.B(n_104),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B(n_49),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_40),
.B(n_51),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_40),
.B(n_104),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_53)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_46),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_45),
.A2(n_58),
.B(n_180),
.C(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_45),
.B(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_46),
.B(n_59),
.C(n_61),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_52),
.A2(n_93),
.B(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_52),
.A2(n_125),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_52),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_52),
.A2(n_92),
.B1(n_187),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_52),
.A2(n_92),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_52),
.A2(n_92),
.B1(n_196),
.B2(n_206),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_68),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_64),
.B(n_66),
.Y(n_55)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_56),
.B(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_56),
.A2(n_107),
.B1(n_110),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_56),
.A2(n_110),
.B1(n_162),
.B2(n_181),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_57),
.A2(n_108),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_62),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_78),
.B(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g181 ( 
.A(n_62),
.B(n_104),
.CON(n_181),
.SN(n_181)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_75),
.B1(n_80),
.B2(n_82),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_69),
.Y(n_116)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_75),
.A2(n_82),
.B1(n_114),
.B2(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_80),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_94),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_92),
.B(n_153),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_95),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.C(n_111),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_96),
.A2(n_97),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_105),
.B(n_111),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_141),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_126),
.B1(n_139),
.B2(n_140),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_171),
.B(n_246),
.C(n_250),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_164),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_154),
.C(n_156),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_146),
.B(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_156),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.C(n_160),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_160),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_241),
.B(n_245),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_197),
.B(n_240),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_192),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_192),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_184),
.C(n_189),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_183),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B(n_188),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.C(n_195),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_195),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_235),
.B(n_239),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_225),
.B(n_234),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_214),
.B(n_224),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_207),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_220),
.B(n_223),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_230),
.C(n_233),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_238),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_244),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_249),
.Y(n_250)
);


endmodule