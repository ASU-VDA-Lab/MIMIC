module fake_jpeg_5822_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_31),
.Y(n_60)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_17),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_66),
.B1(n_19),
.B2(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_18),
.B1(n_25),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_17),
.B1(n_19),
.B2(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_17),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_30),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_18),
.B1(n_29),
.B2(n_28),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_79),
.B1(n_80),
.B2(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_57),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_22),
.B1(n_33),
.B2(n_34),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_22),
.B1(n_33),
.B2(n_34),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_33),
.B1(n_28),
.B2(n_32),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_65),
.B(n_24),
.C(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_28),
.B1(n_20),
.B2(n_30),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_64),
.B1(n_21),
.B2(n_23),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_58),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_30),
.B1(n_20),
.B2(n_32),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_32),
.B1(n_21),
.B2(n_23),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_31),
.B(n_21),
.C(n_37),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_77),
.B(n_73),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_41),
.C(n_36),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_57),
.C(n_47),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_106),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_105),
.C(n_78),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_119),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_85),
.B1(n_94),
.B2(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_118),
.B1(n_69),
.B2(n_75),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_112),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_117),
.Y(n_135)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_109),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_118),
.B1(n_99),
.B2(n_83),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_1),
.Y(n_112)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_49),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_95),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_77),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_58),
.B1(n_21),
.B2(n_27),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_83),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_53),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_141),
.B1(n_147),
.B2(n_103),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_88),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_128),
.A2(n_133),
.B(n_143),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_108),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_139),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_93),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_103),
.C(n_98),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_95),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_151),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_106),
.A3(n_120),
.B1(n_97),
.B2(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_149),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_97),
.A2(n_89),
.B(n_92),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_116),
.B(n_107),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_89),
.B1(n_92),
.B2(n_87),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_84),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_111),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_161),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_176),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_128),
.C(n_152),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_100),
.B1(n_104),
.B2(n_118),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_169),
.B1(n_170),
.B2(n_178),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_173),
.B1(n_130),
.B2(n_129),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_104),
.B1(n_119),
.B2(n_101),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_101),
.B1(n_117),
.B2(n_110),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_181),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_102),
.B1(n_110),
.B2(n_87),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_24),
.B(n_31),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_145),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_128),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_102),
.B1(n_87),
.B2(n_74),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_47),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_140),
.B(n_125),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_177),
.B(n_143),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_171),
.C(n_175),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_142),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_190),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_150),
.B1(n_136),
.B2(n_129),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_191),
.B1(n_202),
.B2(n_170),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_192),
.B(n_208),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_123),
.B(n_138),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_152),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_199),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_206),
.B(n_154),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_143),
.C(n_149),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_151),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_210),
.C(n_154),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_151),
.B1(n_132),
.B2(n_74),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_151),
.B1(n_132),
.B2(n_95),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_209),
.B1(n_153),
.B2(n_163),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_167),
.C(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_157),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_31),
.B(n_24),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_84),
.B1(n_56),
.B2(n_27),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_157),
.B(n_182),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_159),
.B(n_183),
.C(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_219),
.B1(n_227),
.B2(n_229),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_233),
.C(n_190),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_156),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_215),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_228),
.B(n_172),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_161),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

XNOR2x2_ASAP7_75t_SL g255 ( 
.A(n_224),
.B(n_24),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_160),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_226),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_156),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_183),
.B1(n_158),
.B2(n_153),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_174),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_158),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_239),
.C(n_252),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_207),
.C(n_199),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_250),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_184),
.B1(n_206),
.B2(n_193),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_251),
.B1(n_235),
.B2(n_214),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_210),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_255),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_188),
.B1(n_202),
.B2(n_198),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_208),
.C(n_198),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_162),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_254),
.C(n_234),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_41),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_222),
.B1(n_224),
.B2(n_219),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_262),
.B(n_243),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_263),
.C(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_234),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_211),
.C(n_56),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_211),
.C(n_84),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_31),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_11),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_268),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_243),
.B1(n_240),
.B2(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_11),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_23),
.B1(n_3),
.B2(n_5),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_248),
.B1(n_254),
.B2(n_12),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_277),
.B1(n_2),
.B2(n_3),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_245),
.B(n_247),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_280),
.B(n_281),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_31),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_24),
.C(n_3),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_2),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_258),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_264),
.Y(n_285)
);

AOI31xp33_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_290),
.A3(n_282),
.B(n_279),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_288),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_265),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_264),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_285),
.Y(n_302)
);

AOI31xp33_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_265),
.A3(n_283),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_294),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_295),
.C(n_11),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_276),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_304),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_24),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

OAI221xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.C(n_9),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_14),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_13),
.C(n_15),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_6),
.B(n_7),
.Y(n_309)
);

AOI31xp67_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_16),
.A3(n_9),
.B(n_13),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_309),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_291),
.B(n_7),
.C(n_8),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_308),
.B(n_300),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_299),
.B(n_305),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_307),
.B1(n_7),
.B2(n_8),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_7),
.B(n_8),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_8),
.Y(n_317)
);


endmodule