module fake_jpeg_8752_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_39),
.B(n_40),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_18),
.B1(n_35),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_70),
.B1(n_23),
.B2(n_26),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_35),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_26),
.B(n_33),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_18),
.B1(n_25),
.B2(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_71),
.B1(n_15),
.B2(n_14),
.Y(n_116)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_65),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_27),
.C(n_22),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_30),
.C(n_24),
.Y(n_111)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_19),
.B1(n_18),
.B2(n_25),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_34),
.B1(n_33),
.B2(n_20),
.Y(n_71)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_16),
.B1(n_21),
.B2(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_90),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_16),
.B1(n_21),
.B2(n_28),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_16),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_88),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_28),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_48),
.B(n_23),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_111),
.Y(n_140)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_101),
.B(n_1),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_23),
.B1(n_12),
.B2(n_15),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_108),
.B1(n_110),
.B2(n_115),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_114),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_30),
.B1(n_24),
.B2(n_27),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_109),
.B1(n_116),
.B2(n_14),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_69),
.B1(n_50),
.B2(n_73),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_48),
.B(n_27),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_58),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_42),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_42),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_50),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_58),
.A2(n_30),
.B1(n_24),
.B2(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_72),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_80),
.A2(n_42),
.B1(n_38),
.B2(n_48),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_138),
.B1(n_144),
.B2(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_0),
.Y(n_132)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_145),
.B1(n_137),
.B2(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_38),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_0),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_84),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_138)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

NOR2x1p5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_1),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_93),
.B(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_91),
.B(n_1),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_5),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_3),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_155),
.B(n_157),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_165),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_151),
.B(n_153),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_112),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_174),
.C(n_131),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_110),
.B(n_115),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_99),
.B(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_106),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_161),
.B(n_168),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_114),
.B1(n_100),
.B2(n_104),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_134),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_100),
.B1(n_104),
.B2(n_102),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_102),
.B1(n_105),
.B2(n_108),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_171),
.B1(n_182),
.B2(n_126),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_3),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_172),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_96),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_117),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_96),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_146),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_5),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_146),
.B(n_7),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_133),
.A2(n_97),
.B1(n_95),
.B2(n_106),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_144),
.B1(n_134),
.B2(n_143),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_141),
.B1(n_138),
.B2(n_146),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

AOI22x1_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_142),
.B1(n_127),
.B2(n_123),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_183),
.A2(n_211),
.B(n_212),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_120),
.CI(n_124),
.CON(n_184),
.SN(n_184)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_184),
.B(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_202),
.C(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_142),
.B1(n_123),
.B2(n_148),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_209),
.B1(n_177),
.B2(n_168),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_194),
.B1(n_206),
.B2(n_213),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_120),
.B1(n_146),
.B2(n_134),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_196),
.B(n_198),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_207),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_124),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_167),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_120),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_154),
.A2(n_171),
.B1(n_160),
.B2(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_120),
.C(n_139),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_173),
.C(n_158),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_146),
.B1(n_139),
.B2(n_101),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_154),
.A2(n_97),
.B1(n_92),
.B2(n_81),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_143),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_156),
.B(n_6),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_170),
.Y(n_221)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_229),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_156),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_230),
.C(n_233),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_186),
.Y(n_252)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_231),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_178),
.B1(n_181),
.B2(n_173),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_234),
.B1(n_194),
.B2(n_183),
.Y(n_258)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_185),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_158),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_182),
.C(n_165),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_210),
.C(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_198),
.B1(n_200),
.B2(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_251),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_214),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_223),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_263),
.C(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_222),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_266),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_189),
.B1(n_187),
.B2(n_211),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_241),
.A2(n_212),
.B1(n_184),
.B2(n_177),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_184),
.B(n_202),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_201),
.C(n_113),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_216),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_225),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_113),
.B1(n_7),
.B2(n_8),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_271),
.C(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_219),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_262),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_277),
.C(n_281),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_218),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_230),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_233),
.C(n_231),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_258),
.B(n_223),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_280),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_220),
.C(n_221),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_241),
.C(n_242),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_250),
.B(n_217),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_251),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_227),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_284),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_254),
.A2(n_232),
.B1(n_113),
.B2(n_9),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_266),
.B1(n_249),
.B2(n_250),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_254),
.B1(n_256),
.B2(n_264),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_299),
.B1(n_253),
.B2(n_267),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_257),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_296),
.B(n_300),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_294),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_261),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_301),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_245),
.B1(n_256),
.B2(n_259),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_283),
.A2(n_245),
.B1(n_261),
.B2(n_247),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_272),
.C(n_277),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_305),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_271),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_314),
.Y(n_316)
);

AO22x1_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_251),
.B1(n_244),
.B2(n_280),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_310),
.B(n_292),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_273),
.C(n_7),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_287),
.C(n_296),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_290),
.B(n_6),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_6),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_295),
.B(n_10),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_299),
.B1(n_294),
.B2(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_9),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_309),
.A2(n_293),
.B(n_287),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.C(n_307),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_293),
.B1(n_10),
.B2(n_11),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_305),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_328),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_330),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_308),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_319),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_316),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_320),
.Y(n_336)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_329),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_335),
.B1(n_327),
.B2(n_317),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_324),
.B(n_334),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_315),
.B(n_333),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_331),
.B(n_11),
.Y(n_341)
);


endmodule