module fake_jpeg_22049_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_34),
.B(n_36),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_2),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_2),
.B(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_4),
.Y(n_63)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_4),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_52),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_17),
.B1(n_21),
.B2(n_31),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_64),
.B1(n_68),
.B2(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_49),
.A2(n_62),
.B(n_72),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_27),
.B1(n_24),
.B2(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_24),
.B1(n_29),
.B2(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_33),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_25),
.B1(n_23),
.B2(n_7),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_58),
.B1(n_73),
.B2(n_54),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_42),
.B1(n_44),
.B2(n_23),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_96),
.B1(n_100),
.B2(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_86),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_43),
.B(n_44),
.C(n_15),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_91),
.B(n_98),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_89),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_45),
.CI(n_33),
.CON(n_82),
.SN(n_82)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_88),
.CI(n_20),
.CON(n_118),
.SN(n_118)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_5),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_45),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_20),
.CI(n_6),
.CON(n_88),
.SN(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_5),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_5),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_48),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_R g101 ( 
.A1(n_93),
.A2(n_54),
.B(n_20),
.C(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_105),
.Y(n_132)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_107),
.Y(n_129)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_50),
.C(n_74),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_94),
.C(n_76),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_58),
.B(n_50),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_118),
.B(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_73),
.B1(n_20),
.B2(n_74),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_115),
.B1(n_87),
.B2(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_117),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_20),
.B1(n_53),
.B2(n_55),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_121),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_55),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_98),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_85),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_127),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_78),
.C(n_88),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_103),
.C(n_83),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_135),
.B1(n_138),
.B2(n_132),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_136),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_140),
.C(n_122),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_82),
.B1(n_88),
.B2(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_82),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_84),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_143),
.B(n_117),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_83),
.C(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_110),
.B1(n_109),
.B2(n_118),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_149),
.B1(n_123),
.B2(n_135),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_118),
.B1(n_115),
.B2(n_105),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_139),
.C(n_140),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_163),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_131),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_150),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_128),
.C(n_136),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_125),
.B(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_165),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_174),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_172),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_144),
.B1(n_149),
.B2(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_154),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_162),
.A3(n_156),
.B1(n_165),
.B2(n_157),
.C1(n_141),
.C2(n_106),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_167),
.B(n_168),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_106),
.C(n_55),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_173),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_14),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_14),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_181),
.C(n_182),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_182),
.A2(n_176),
.B(n_178),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_184),
.A2(n_87),
.B(n_20),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_179),
.B(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.Y(n_187)
);


endmodule