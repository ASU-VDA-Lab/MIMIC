module real_jpeg_7443_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_2),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_2),
.A2(n_35),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_80),
.B1(n_181),
.B2(n_185),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_80),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_4),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_4),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_4),
.A2(n_148),
.B1(n_197),
.B2(n_281),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_4),
.A2(n_148),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_4),
.A2(n_148),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_5),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_5),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_5),
.A2(n_153),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_5),
.A2(n_153),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_5),
.A2(n_153),
.B1(n_275),
.B2(n_316),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_6),
.A2(n_54),
.B1(n_119),
.B2(n_123),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_6),
.A2(n_54),
.B1(n_271),
.B2(n_275),
.Y(n_270)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_9),
.Y(n_130)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_9),
.Y(n_263)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_11),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_11),
.A2(n_51),
.B1(n_55),
.B2(n_266),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_11),
.B(n_304),
.C(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_11),
.B(n_101),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_11),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_11),
.B(n_86),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_11),
.B(n_256),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_12),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_12),
.Y(n_147)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_12),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_12),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_13),
.A2(n_42),
.B1(n_164),
.B2(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_14),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_14),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_14),
.A2(n_114),
.B1(n_160),
.B2(n_175),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_114),
.B1(n_232),
.B2(n_236),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_14),
.A2(n_114),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_15),
.A2(n_131),
.B1(n_132),
.B2(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_15),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_15),
.A2(n_55),
.B1(n_82),
.B2(n_192),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_15),
.A2(n_192),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_15),
.A2(n_143),
.B1(n_192),
.B2(n_200),
.Y(n_392)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_16),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_240),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_239),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_203),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_20),
.B(n_203),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_156),
.C(n_170),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_21),
.B(n_156),
.CI(n_170),
.CON(n_283),
.SN(n_283)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_87),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_22),
.B(n_88),
.C(n_126),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_23),
.B(n_49),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_38),
.B2(n_41),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_24),
.A2(n_41),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_24),
.A2(n_167),
.B1(n_269),
.B2(n_277),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_24),
.A2(n_309),
.B(n_313),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_24),
.A2(n_266),
.B(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_25),
.A2(n_180),
.B1(n_186),
.B2(n_187),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_25),
.B(n_315),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_25),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_25),
.A2(n_270),
.B1(n_369),
.B2(n_397),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_27),
.Y(n_329)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_27),
.Y(n_346)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_27),
.Y(n_398)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_28),
.Y(n_185)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_31),
.Y(n_186)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_32),
.Y(n_370)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_33),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_34),
.Y(n_274)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_40),
.Y(n_374)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_43),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_48),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B1(n_79),
.B2(n_86),
.Y(n_49)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_50),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_52),
.Y(n_162)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_52),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_53),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_56),
.A2(n_79),
.B1(n_86),
.B2(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_56),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_56),
.A2(n_86),
.B1(n_159),
.B2(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_56),
.B(n_295),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_71),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_64),
.B2(n_68),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_60),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g378 ( 
.A(n_68),
.Y(n_378)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_69),
.Y(n_296)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_71),
.A2(n_173),
.B1(n_174),
.B2(n_178),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_71),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_71),
.A2(n_173),
.B1(n_320),
.B2(n_357),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_71),
.A2(n_174),
.B(n_321),
.Y(n_419)
);

AOI22x1_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_74),
.Y(n_372)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_75),
.Y(n_306)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_82),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_85),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_86),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_126),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_89),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_89),
.A2(n_117),
.B1(n_280),
.B2(n_392),
.Y(n_418)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B1(n_98),
.B2(n_99),
.Y(n_90)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_91),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_97),
.Y(n_259)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_100),
.Y(n_281)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_101),
.A2(n_194),
.B1(n_195),
.B2(n_202),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_101),
.A2(n_194),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_104),
.Y(n_379)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_116),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_117),
.B(n_196),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_117),
.A2(n_392),
.B(n_393),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_119),
.B(n_262),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_145),
.B(n_151),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_127),
.A2(n_138),
.B1(n_145),
.B2(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_128),
.B(n_152),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_128),
.A2(n_413),
.B(n_416),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_138),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_133),
.Y(n_260)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_138),
.B(n_266),
.Y(n_395)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_140),
.Y(n_363)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_151),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_155),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_166),
.B2(n_169),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_166),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_166),
.A2(n_169),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_167),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_167),
.A2(n_333),
.B(n_338),
.Y(n_332)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_189),
.C(n_193),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_171),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_172),
.B(n_179),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_173),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_173),
.A2(n_294),
.B(n_357),
.Y(n_388)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_180),
.Y(n_277)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_185),
.B(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_238),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_193),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_194),
.A2(n_279),
.B(n_282),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_194),
.A2(n_282),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_194),
.B(n_195),
.Y(n_393)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_224),
.B2(n_225),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_216),
.B(n_223),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_284),
.B(n_444),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_283),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_243),
.B(n_283),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.C(n_249),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_248),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_249),
.B(n_434),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_278),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_250),
.A2(n_251),
.B1(n_278),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_253),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_267),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_254),
.A2(n_267),
.B1(n_268),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_254),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_260),
.A3(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_SL g413 ( 
.A1(n_265),
.A2(n_266),
.B(n_414),
.Y(n_413)
);

OAI21xp33_ASAP7_75t_SL g362 ( 
.A1(n_266),
.A2(n_363),
.B(n_364),
.Y(n_362)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_273),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_278),
.Y(n_429)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_283),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_422),
.B(n_441),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_401),
.B(n_421),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_383),
.B(n_400),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_351),
.B(n_382),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_324),
.B(n_350),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_307),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_307),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_292),
.A2(n_299),
.B1(n_300),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_318),
.C(n_323),
.Y(n_352)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_341),
.B(n_349),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_331),
.B(n_340),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_339),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_339),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_338),
.A2(n_368),
.B(n_373),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_347),
.Y(n_349)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_353),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_366),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_360),
.B2(n_361),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_360),
.C(n_366),
.Y(n_384)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AOI32xp33_ASAP7_75t_L g375 ( 
.A1(n_365),
.A2(n_376),
.A3(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_375),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_375),
.Y(n_389)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_384),
.B(n_385),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_390),
.B2(n_399),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_389),
.C(n_399),
.Y(n_402)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_390),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_395),
.C(n_396),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_402),
.B(n_403),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_410),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_405),
.Y(n_409)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_409),
.C(n_410),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_417),
.B2(n_420),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_418),
.C(n_419),
.Y(n_432)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx8_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_417),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_436),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_425),
.A2(n_442),
.B(n_443),
.Y(n_441)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_433),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_433),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.C(n_432),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_430),
.A2(n_431),
.B1(n_432),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_432),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_438),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);


endmodule