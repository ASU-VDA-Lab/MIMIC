module fake_jpeg_15860_n_113 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

NOR3xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_12),
.C(n_15),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_33),
.B(n_12),
.C(n_21),
.Y(n_47)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_25),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_14),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_16),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_42),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_50),
.Y(n_58)
);

AOI32xp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_27),
.A3(n_22),
.B1(n_13),
.B2(n_20),
.Y(n_45)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_11),
.C(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_15),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_21),
.Y(n_57)
);

BUFx24_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_18),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_59),
.B1(n_64),
.B2(n_20),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_25),
.C(n_10),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_66),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_26),
.B1(n_17),
.B2(n_18),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_2),
.B(n_3),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_3),
.B(n_4),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_11),
.C(n_10),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_74),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_40),
.B(n_41),
.C(n_38),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_77),
.B(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_81),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_56),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_58),
.C(n_59),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_86),
.C(n_80),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_68),
.B1(n_60),
.B2(n_57),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_87),
.B1(n_77),
.B2(n_70),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_67),
.C(n_56),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_11),
.B(n_4),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_94),
.B(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_78),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_87),
.Y(n_98)
);

AO221x1_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_62),
.B1(n_53),
.B2(n_51),
.C(n_72),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_96),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_78),
.B(n_92),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_91),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

OAI31xp33_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_99),
.A3(n_62),
.B(n_8),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_105),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_88),
.B1(n_83),
.B2(n_86),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_3),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C1(n_99),
.C2(n_109),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_6),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.C(n_106),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_108),
.Y(n_113)
);


endmodule