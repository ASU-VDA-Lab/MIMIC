module fake_jpeg_26559_n_195 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_195);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_15),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_32),
.Y(n_60)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_11),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_44),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_10),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_31),
.B1(n_18),
.B2(n_30),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_51),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_62),
.B1(n_68),
.B2(n_19),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_29),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_31),
.B(n_21),
.C(n_28),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_60),
.B(n_19),
.Y(n_81)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_32),
.C(n_25),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_65),
.C(n_59),
.Y(n_90)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_16),
.B1(n_28),
.B2(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_32),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_27),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_21),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_27),
.C(n_17),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_34),
.A2(n_16),
.B1(n_24),
.B2(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_85),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_0),
.B(n_1),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_81),
.B(n_3),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_9),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_88),
.Y(n_108)
);

AO21x2_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_23),
.B(n_19),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_53),
.B1(n_57),
.B2(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_9),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_48),
.C(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_2),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_83),
.C(n_69),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_118),
.B(n_87),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_116),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_52),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_56),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_54),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_23),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_79),
.C(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_114),
.B(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_57),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_126),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_84),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_131),
.B(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_87),
.B(n_78),
.C(n_83),
.Y(n_131)
);

NOR4xp25_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_81),
.C(n_83),
.D(n_75),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_102),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_98),
.C(n_117),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_128),
.B(n_131),
.C(n_109),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_142),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_146),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_97),
.B1(n_106),
.B2(n_103),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_97),
.B1(n_126),
.B2(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_108),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_163),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_138),
.C(n_135),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_142),
.C(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_165),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_113),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_153),
.B(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_106),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_120),
.B1(n_149),
.B2(n_124),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_103),
.B1(n_123),
.B2(n_91),
.Y(n_174)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_115),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_153),
.B1(n_145),
.B2(n_143),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_158),
.B1(n_156),
.B2(n_154),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_174),
.B(n_69),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.C(n_173),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_130),
.C(n_116),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_104),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_176),
.B1(n_170),
.B2(n_171),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_115),
.B1(n_155),
.B2(n_113),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_105),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_180),
.A2(n_181),
.B1(n_169),
.B2(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_96),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_180),
.A2(n_70),
.B1(n_93),
.B2(n_105),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_4),
.B(n_5),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_70),
.C(n_63),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_70),
.A3(n_63),
.B1(n_23),
.B2(n_7),
.C1(n_3),
.C2(n_5),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_190),
.C(n_186),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_192),
.B(n_4),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_189),
.B(n_184),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);


endmodule