module fake_jpeg_30288_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_2),
.CON(n_67),
.SN(n_67)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_58),
.Y(n_82)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_60),
.B(n_47),
.C(n_50),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_2),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_54),
.B1(n_61),
.B2(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_83),
.B1(n_57),
.B2(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_4),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_61),
.CON(n_80),
.SN(n_80)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_5),
.Y(n_99)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_80),
.B(n_74),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_57),
.B1(n_54),
.B2(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_97),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_93),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_56),
.C(n_53),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_100),
.C(n_25),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_10),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_28),
.C(n_40),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_26),
.B(n_38),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_29),
.B1(n_11),
.B2(n_13),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_115),
.B1(n_10),
.B2(n_39),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_6),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_27),
.B1(n_37),
.B2(n_36),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_8),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_9),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_121),
.C(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_135),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_35),
.B1(n_15),
.B2(n_16),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_132),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_33),
.B1(n_24),
.B2(n_30),
.Y(n_132)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_23),
.B(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_104),
.B(n_116),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_139),
.B1(n_127),
.B2(n_131),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_122),
.B(n_115),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_113),
.C(n_121),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_133),
.B(n_135),
.C(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_142),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_137),
.C(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_148),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_141),
.B(n_125),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_109),
.C(n_133),
.Y(n_151)
);


endmodule