module fake_netlist_1_11937_n_27 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
OAI21x1_ASAP7_75t_L g15 ( .A1(n_5), .A2(n_7), .B(n_8), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_9), .B(n_10), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
AO21x1_ASAP7_75t_SL g20 ( .A1(n_18), .A2(n_17), .B(n_0), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_14), .Y(n_22) );
O2A1O1Ixp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_19), .B(n_15), .C(n_3), .Y(n_23) );
NAND2xp5_ASAP7_75t_SL g24 ( .A(n_23), .B(n_1), .Y(n_24) );
INVx5_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
OAI22x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_2), .B1(n_6), .B2(n_11), .Y(n_26) );
BUFx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
endmodule