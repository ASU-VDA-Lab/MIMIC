module fake_jpeg_29717_n_425 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_425);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_425;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_50),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_14),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_41),
.Y(n_110)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_13),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_54),
.B(n_76),
.Y(n_136)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_77),
.Y(n_118)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_80),
.Y(n_131)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_9),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_9),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_85),
.Y(n_105)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_86),
.Y(n_119)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_18),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_0),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_90),
.B(n_97),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_22),
.B(n_25),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_93),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_65),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_102),
.B(n_104),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_42),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_117),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_114),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_40),
.B(n_25),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g179 ( 
.A(n_112),
.B(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_66),
.B(n_19),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_70),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_128),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_123),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_67),
.A2(n_19),
.B1(n_39),
.B2(n_36),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_125),
.A2(n_133),
.B1(n_94),
.B2(n_96),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_58),
.A2(n_40),
.B1(n_25),
.B2(n_22),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_74),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_46),
.A2(n_40),
.B1(n_31),
.B2(n_30),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_82),
.B(n_0),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_1),
.C(n_2),
.Y(n_174)
);

OR2x2_ASAP7_75t_SL g135 ( 
.A(n_69),
.B(n_39),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_60),
.B(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_1),
.Y(n_172)
);

OR2x4_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_31),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_135),
.B(n_109),
.C(n_131),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_71),
.A2(n_23),
.B1(n_37),
.B2(n_38),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_123),
.B1(n_126),
.B2(n_23),
.Y(n_162)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_147),
.Y(n_222)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_150),
.A2(n_196),
.B(n_139),
.Y(n_219)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_30),
.B(n_38),
.C(n_37),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_153),
.B(n_156),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_105),
.A2(n_59),
.B1(n_75),
.B2(n_73),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_157),
.A2(n_162),
.B1(n_168),
.B2(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_21),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_170),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_111),
.Y(n_164)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_64),
.B1(n_63),
.B2(n_56),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_165),
.A2(n_166),
.B1(n_175),
.B2(n_180),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_51),
.B1(n_49),
.B2(n_76),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_95),
.A2(n_21),
.B1(n_17),
.B2(n_74),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_17),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_110),
.B(n_17),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_185),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_4),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_118),
.A2(n_4),
.B(n_5),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_181),
.A2(n_115),
.B1(n_116),
.B2(n_137),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_124),
.A2(n_93),
.B(n_99),
.C(n_113),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_186),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_113),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_103),
.B(n_5),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_188),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_107),
.B(n_7),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_113),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_7),
.B1(n_8),
.B2(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_103),
.B(n_8),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_140),
.B1(n_142),
.B2(n_94),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_145),
.B1(n_140),
.B2(n_129),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_130),
.B1(n_108),
.B2(n_127),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_130),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_194),
.B(n_198),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_127),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_139),
.B(n_138),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_150),
.B(n_138),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_227),
.Y(n_240)
);

OAI22x1_ASAP7_75t_SL g213 ( 
.A1(n_173),
.A2(n_179),
.B1(n_162),
.B2(n_182),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g252 ( 
.A1(n_213),
.A2(n_231),
.B(n_208),
.C(n_229),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_137),
.B(n_111),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_217),
.A2(n_231),
.B(n_159),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_225),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_234),
.B1(n_236),
.B2(n_183),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_171),
.B(n_91),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_154),
.B(n_91),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_230),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_167),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_179),
.A2(n_137),
.B(n_108),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_169),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_158),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_164),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_189),
.A2(n_116),
.B1(n_170),
.B2(n_155),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_160),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_243),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_155),
.B1(n_152),
.B2(n_180),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_244),
.B1(n_258),
.B2(n_200),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_188),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_176),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_156),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_249),
.B(n_255),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_SL g287 ( 
.A1(n_252),
.A2(n_272),
.B(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_205),
.Y(n_255)
);

AO22x2_ASAP7_75t_L g257 ( 
.A1(n_213),
.A2(n_180),
.B1(n_153),
.B2(n_187),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_264),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_202),
.A2(n_180),
.B1(n_178),
.B2(n_192),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_230),
.B(n_185),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_186),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_207),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_199),
.B(n_174),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_194),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_215),
.Y(n_274)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_209),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_209),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_273),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_221),
.B(n_151),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_199),
.B(n_197),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_298),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_226),
.B1(n_200),
.B2(n_234),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_280),
.A2(n_283),
.B1(n_295),
.B2(n_224),
.Y(n_326)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_247),
.Y(n_281)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_226),
.B1(n_233),
.B2(n_216),
.Y(n_283)
);

CKINVDCx10_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_285),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_288),
.B1(n_292),
.B2(n_244),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_264),
.A2(n_237),
.B1(n_216),
.B2(n_222),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_SL g292 ( 
.A1(n_272),
.A2(n_204),
.B(n_214),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_240),
.A2(n_252),
.B1(n_244),
.B2(n_257),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_266),
.B(n_206),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_243),
.B(n_239),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_303),
.Y(n_312)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_206),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_256),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_203),
.B(n_211),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_304),
.B(n_315),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_305),
.A2(n_282),
.B(n_289),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_306),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_246),
.C(n_252),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_SL g346 ( 
.A1(n_307),
.A2(n_262),
.A3(n_116),
.B1(n_197),
.B2(n_193),
.C1(n_214),
.C2(n_237),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_274),
.B(n_241),
.C(n_245),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_309),
.C(n_313),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_286),
.C(n_275),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_265),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_248),
.C(n_252),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_276),
.Y(n_314)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

OA21x2_ASAP7_75t_SL g315 ( 
.A1(n_284),
.A2(n_285),
.B(n_275),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_257),
.B1(n_259),
.B2(n_253),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_319),
.B1(n_321),
.B2(n_327),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_257),
.C(n_211),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_290),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_254),
.B1(n_269),
.B2(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_278),
.A2(n_250),
.B1(n_247),
.B2(n_262),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_297),
.B(n_293),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_323),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_250),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_294),
.B1(n_224),
.B2(n_268),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_280),
.B1(n_302),
.B2(n_299),
.Y(n_327)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_312),
.B(n_290),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_334),
.A2(n_344),
.B(n_336),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_335),
.B(n_346),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_296),
.Y(n_336)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_337),
.B(n_204),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_270),
.Y(n_339)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_339),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_340),
.A2(n_330),
.B1(n_319),
.B2(n_320),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_294),
.B(n_203),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_327),
.A2(n_316),
.B1(n_318),
.B2(n_310),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_321),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_313),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_309),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_238),
.Y(n_350)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_235),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_315),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_335),
.B(n_308),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_358),
.Y(n_381)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_322),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_332),
.A2(n_324),
.B1(n_310),
.B2(n_306),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_359),
.A2(n_364),
.B1(n_338),
.B2(n_345),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_357),
.B1(n_360),
.B2(n_362),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_365),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_329),
.C(n_235),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_368),
.C(n_369),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_329),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_367),
.B(n_349),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_147),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_148),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_371),
.C(n_337),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_193),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_343),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_372),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_386),
.Y(n_390)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_375),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_376),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_370),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_331),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_382),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_361),
.A2(n_342),
.B(n_331),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_356),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_350),
.C(n_338),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_384),
.B(n_385),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_347),
.C(n_344),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_349),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_359),
.A2(n_340),
.B1(n_347),
.B2(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_365),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_397),
.Y(n_403)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_381),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_393),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_363),
.C(n_369),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_395),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_382),
.Y(n_407)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_390),
.A2(n_383),
.B(n_378),
.Y(n_400)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_384),
.C(n_385),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_404),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_376),
.Y(n_404)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_396),
.A2(n_379),
.B(n_388),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_389),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_382),
.B(n_373),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_406),
.B(n_407),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_353),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_411),
.Y(n_417)
);

AOI322xp5_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_352),
.A3(n_353),
.B1(n_334),
.B2(n_377),
.C1(n_373),
.C2(n_380),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_399),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_SL g414 ( 
.A1(n_409),
.A2(n_401),
.B(n_368),
.C(n_403),
.Y(n_414)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_414),
.Y(n_419)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_412),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_415),
.A2(n_416),
.B(n_410),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_418),
.B(n_414),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_417),
.A2(n_408),
.B(n_403),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_419),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_421),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_422),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_424),
.Y(n_425)
);


endmodule