module fake_netlist_5_1865_n_151 (n_54, n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_36, n_25, n_53, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_51, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_55, n_14, n_48, n_2, n_31, n_23, n_13, n_50, n_3, n_49, n_52, n_6, n_39, n_151);

input n_54;
input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_36;
input n_25;
input n_53;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_51;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_55;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_50;
input n_3;
input n_49;
input n_52;
input n_6;
input n_39;

output n_151;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_117;
wire n_94;
wire n_113;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_126;
wire n_84;
wire n_130;
wire n_79;
wire n_131;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_99;
wire n_147;
wire n_67;
wire n_121;
wire n_76;
wire n_87;
wire n_150;
wire n_77;
wire n_64;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_104;
wire n_103;
wire n_56;
wire n_63;
wire n_97;
wire n_141;
wire n_145;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_16),
.B1(n_44),
.B2(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_2),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_41),
.B1(n_49),
.B2(n_1),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_12),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_1),
.A2(n_39),
.B1(n_4),
.B2(n_14),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_50),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_15),
.B(n_46),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_22),
.A2(n_38),
.B1(n_40),
.B2(n_33),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_45),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_3),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_R g81 ( 
.A(n_48),
.B(n_0),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_26),
.B(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_8),
.B1(n_13),
.B2(n_21),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_31),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_34),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_37),
.B(n_53),
.C(n_55),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

AND2x6_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_82),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_74),
.B1(n_61),
.B2(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_89),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_86),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_69),
.B1(n_72),
.B2(n_77),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_88),
.B(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

OAI21x1_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_68),
.B(n_85),
.Y(n_115)
);

OAI21x1_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_58),
.B(n_62),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_64),
.B1(n_71),
.B2(n_84),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_69),
.B(n_70),
.C(n_77),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_110),
.B(n_104),
.C(n_108),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_91),
.B(n_111),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_100),
.B1(n_92),
.B2(n_102),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_90),
.B1(n_95),
.B2(n_98),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_106),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_98),
.B1(n_111),
.B2(n_99),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_96),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_114),
.Y(n_130)
);

OR2x6_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_101),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_96),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_118),
.B1(n_120),
.B2(n_96),
.C(n_116),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_116),
.Y(n_139)
);

OAI321xp33_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_131),
.A3(n_130),
.B1(n_128),
.B2(n_118),
.C(n_126),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_131),
.B1(n_115),
.B2(n_112),
.Y(n_141)
);

AOI221xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_128),
.B1(n_96),
.B2(n_125),
.C(n_99),
.Y(n_142)
);

NAND4xp25_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_125),
.C(n_98),
.D(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_141),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_139),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_145),
.A2(n_140),
.B1(n_99),
.B2(n_142),
.Y(n_148)
);

OAI31xp33_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_137),
.A3(n_145),
.B(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

AO221x1_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_148),
.B1(n_149),
.B2(n_137),
.C(n_99),
.Y(n_151)
);


endmodule