module real_jpeg_18108_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_351),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_0),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_1),
.B(n_39),
.Y(n_38)
);

NAND2x1_ASAP7_75t_SL g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

NAND2x1_ASAP7_75t_L g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_1),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_1),
.B(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_4),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_5),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_39),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_5),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_6),
.Y(n_120)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_6),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_7),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_7),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_7),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_7),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_7),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_8),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_8),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_8),
.B(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_8),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_8),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_8),
.B(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_9),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_11),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_166),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_164),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_141),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_19),
.B(n_141),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_R g19 ( 
.A(n_20),
.B(n_65),
.C(n_106),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_20),
.B(n_65),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_21),
.B(n_41),
.C(n_52),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_23),
.B(n_32),
.C(n_38),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_23),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_23),
.A2(n_212),
.B(n_213),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

OR2x4_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_35),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_24),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_29),
.Y(n_198)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_32),
.B(n_119),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_32),
.B(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_32),
.B(n_305),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_32),
.A2(n_33),
.B1(n_49),
.B2(n_105),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp5_ASAP7_75t_L g180 ( 
.A1(n_33),
.A2(n_49),
.B(n_181),
.C(n_186),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_33),
.B(n_72),
.C(n_119),
.Y(n_192)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_35),
.Y(n_136)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_36),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_54),
.C(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_37),
.B(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_37),
.A2(n_38),
.B1(n_132),
.B2(n_210),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_38),
.A2(n_69),
.B(n_93),
.Y(n_92)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_69),
.Y(n_93)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_39),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_52),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.C(n_49),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_42),
.A2(n_43),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_42),
.B(n_192),
.C(n_194),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_42),
.A2(n_43),
.B1(n_84),
.B2(n_124),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_43),
.B(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_43),
.B(n_124),
.C(n_269),
.Y(n_293)
);

AO22x1_ASAP7_75t_L g104 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_49),
.A2(n_105),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_50),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_54),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_53),
.B(n_58),
.C(n_62),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_53),
.A2(n_54),
.B1(n_194),
.B2(n_195),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_54),
.B(n_93),
.C(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_61),
.A2(n_62),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_81),
.C(n_84),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_62),
.B(n_75),
.C(n_220),
.Y(n_326)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_90),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_78),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_67),
.B(n_78),
.C(n_90),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_68),
.B(n_72),
.C(n_75),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_69),
.B(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_97),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_97),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_69),
.A2(n_111),
.B1(n_272),
.B2(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_72),
.A2(n_77),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_72),
.A2(n_77),
.B1(n_162),
.B2(n_163),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_79),
.C(n_87),
.Y(n_78)
);

AOI22x1_ASAP7_75t_SL g224 ( 
.A1(n_74),
.A2(n_75),
.B1(n_135),
.B2(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_127),
.C(n_135),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_87),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_75),
.B(n_176),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_80),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_84),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_81),
.A2(n_97),
.B1(n_112),
.B2(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_81),
.B(n_97),
.C(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_114),
.B(n_121),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_84),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_84),
.B(n_115),
.Y(n_201)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_87),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_128),
.C(n_132),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_103),
.Y(n_90)
);

XOR2x1_ASAP7_75t_L g253 ( 
.A(n_91),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_92),
.A2(n_94),
.B1(n_187),
.B2(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_93),
.B(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_94),
.A2(n_187),
.B(n_281),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_95),
.B(n_103),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_96),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_97),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_97),
.A2(n_112),
.B1(n_282),
.B2(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_106),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_126),
.C(n_137),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_107),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.C(n_122),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_113),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_116),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_119),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_118),
.A2(n_119),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_118),
.A2(n_119),
.B1(n_187),
.B2(n_286),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_187),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_SL g296 ( 
.A1(n_119),
.A2(n_186),
.B(n_187),
.C(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_126),
.A2(n_137),
.B1(n_138),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_126),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_127),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_128),
.A2(n_132),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_132),
.Y(n_210)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_155),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_153),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI321xp33_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_244),
.A3(n_261),
.B1(n_344),
.B2(n_345),
.C(n_350),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI31xp33_ASAP7_75t_L g345 ( 
.A1(n_170),
.A2(n_257),
.A3(n_346),
.B(n_349),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_233),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_171),
.B(n_233),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_203),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_172),
.B(n_204),
.C(n_229),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_191),
.C(n_199),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_179),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_174),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_178),
.B(n_180),
.Y(n_336)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_181),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_181),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_181),
.A2(n_269),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_187),
.Y(n_286)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_199),
.B1(n_200),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_228),
.B2(n_229),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_221),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.C(n_219),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_210),
.B(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_210),
.A2(n_271),
.B(n_272),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_212),
.B1(n_219),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_251),
.C(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_234),
.B(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_237),
.B(n_240),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_241),
.B(n_243),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_242),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_257),
.Y(n_244)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_245),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_255),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_246),
.B(n_255),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_253),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_253),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g349 ( 
.A(n_258),
.B(n_260),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_340),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_330),
.B(n_339),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_313),
.B(n_329),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_294),
.B(n_312),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_278),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_278),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.C(n_275),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_271),
.A2(n_275),
.B1(n_276),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_288),
.C(n_293),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_285),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_304),
.B(n_306),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_302),
.B(n_311),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_299),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_308),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_307),
.B(n_310),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_315),
.Y(n_329)
);

XOR2x2_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_319),
.C(n_320),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_325),
.C(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_332),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_335),
.C(n_337),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_342),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);


endmodule