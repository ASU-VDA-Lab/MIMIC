module real_aes_7360_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_1), .A2(n_149), .B(n_154), .C(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_2), .A2(n_144), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g461 ( .A(n_3), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_4), .B(n_168), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_5), .A2(n_15), .B1(n_723), .B2(n_724), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_5), .Y(n_724) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_6), .A2(n_144), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g149 ( .A(n_7), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g178 ( .A(n_8), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_9), .B(n_43), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_9), .B(n_43), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_10), .A2(n_256), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_11), .B(n_159), .Y(n_195) );
INVx1_ASAP7_75t_L g483 ( .A(n_12), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_13), .B(n_158), .Y(n_531) );
INVx1_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_15), .Y(n_723) );
INVx1_ASAP7_75t_L g543 ( .A(n_16), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_17), .A2(n_179), .B(n_204), .C(n_206), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_18), .B(n_168), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_19), .B(n_472), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_20), .B(n_144), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_21), .B(n_264), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_22), .A2(n_158), .B(n_160), .C(n_164), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_23), .B(n_168), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_24), .B(n_159), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_25), .A2(n_162), .B(n_206), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_26), .B(n_159), .Y(n_240) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_27), .Y(n_224) );
INVx1_ASAP7_75t_L g238 ( .A(n_28), .Y(n_238) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_29), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_30), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_31), .B(n_159), .Y(n_462) );
INVx1_ASAP7_75t_L g261 ( .A(n_32), .Y(n_261) );
INVx1_ASAP7_75t_L g496 ( .A(n_33), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_34), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g147 ( .A(n_35), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_36), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_37), .A2(n_158), .B(n_217), .C(n_219), .Y(n_216) );
INVxp67_ASAP7_75t_L g262 ( .A(n_38), .Y(n_262) );
CKINVDCx14_ASAP7_75t_R g215 ( .A(n_39), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_40), .A2(n_154), .B(n_237), .C(n_243), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_41), .A2(n_149), .B(n_154), .C(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_42), .A2(n_92), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_42), .Y(n_128) );
INVx1_ASAP7_75t_L g495 ( .A(n_44), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_45), .A2(n_176), .B(n_177), .C(n_180), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_46), .B(n_159), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_47), .A2(n_125), .B1(n_437), .B2(n_438), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_47), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_48), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_49), .Y(n_258) );
INVx1_ASAP7_75t_L g152 ( .A(n_50), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_51), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_52), .B(n_144), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_53), .A2(n_154), .B1(n_164), .B2(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_54), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_55), .Y(n_458) );
CKINVDCx14_ASAP7_75t_R g174 ( .A(n_56), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_57), .A2(n_176), .B(n_219), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_58), .Y(n_524) );
INVx1_ASAP7_75t_L g480 ( .A(n_59), .Y(n_480) );
INVx1_ASAP7_75t_L g150 ( .A(n_60), .Y(n_150) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
INVx1_ASAP7_75t_SL g218 ( .A(n_62), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_63), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_64), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g227 ( .A(n_65), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_SL g471 ( .A1(n_66), .A2(n_219), .B(n_472), .C(n_473), .Y(n_471) );
INVxp67_ASAP7_75t_L g474 ( .A(n_67), .Y(n_474) );
INVx1_ASAP7_75t_L g116 ( .A(n_68), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_69), .A2(n_144), .B(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_70), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_71), .A2(n_144), .B(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_72), .Y(n_499) );
INVx1_ASAP7_75t_L g518 ( .A(n_73), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_74), .A2(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g202 ( .A(n_75), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_76), .Y(n_235) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_77), .A2(n_449), .B1(n_720), .B2(n_726), .C1(n_730), .C2(n_731), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_78), .A2(n_149), .B(n_154), .C(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_79), .A2(n_144), .B(n_151), .Y(n_143) );
INVx1_ASAP7_75t_L g205 ( .A(n_80), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_81), .B(n_239), .Y(n_512) );
INVx2_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
INVx1_ASAP7_75t_L g192 ( .A(n_83), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_84), .B(n_472), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_85), .A2(n_149), .B(n_154), .C(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g113 ( .A(n_86), .Y(n_113) );
OR2x2_ASAP7_75t_L g441 ( .A(n_86), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g719 ( .A(n_86), .B(n_443), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_87), .A2(n_154), .B(n_226), .C(n_229), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_88), .A2(n_104), .B1(n_117), .B2(n_735), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_89), .A2(n_721), .B1(n_722), .B2(n_725), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_89), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_90), .B(n_171), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_91), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_92), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_93), .A2(n_149), .B(n_154), .C(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_94), .Y(n_535) );
INVx1_ASAP7_75t_L g470 ( .A(n_95), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_96), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_97), .B(n_239), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_98), .B(n_137), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_99), .B(n_137), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g161 ( .A(n_101), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_102), .A2(n_144), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g736 ( .A(n_107), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g443 ( .A(n_112), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g718 ( .A(n_113), .B(n_443), .Y(n_718) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_113), .B(n_442), .Y(n_733) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_447), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g734 ( .A(n_120), .Y(n_734) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_439), .B(n_445), .Y(n_123) );
INVx1_ASAP7_75t_L g438 ( .A(n_125), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_435), .B2(n_436), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_126), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_129), .A2(n_718), .B1(n_727), .B2(n_728), .Y(n_726) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g436 ( .A(n_130), .Y(n_436) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_361), .Y(n_130) );
NOR4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_303), .C(n_333), .D(n_343), .Y(n_131) );
OAI211xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_208), .B(n_266), .C(n_293), .Y(n_132) );
OAI222xp33_ASAP7_75t_L g388 ( .A1(n_133), .A2(n_308), .B1(n_389), .B2(n_390), .C1(n_391), .C2(n_392), .Y(n_388) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_183), .Y(n_133) );
AOI33xp33_ASAP7_75t_L g314 ( .A1(n_134), .A2(n_301), .A3(n_302), .B1(n_315), .B2(n_320), .B3(n_322), .Y(n_314) );
OAI211xp5_ASAP7_75t_SL g371 ( .A1(n_134), .A2(n_372), .B(n_374), .C(n_376), .Y(n_371) );
OR2x2_ASAP7_75t_L g387 ( .A(n_134), .B(n_373), .Y(n_387) );
INVx1_ASAP7_75t_L g420 ( .A(n_134), .Y(n_420) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_170), .Y(n_134) );
INVx2_ASAP7_75t_L g297 ( .A(n_135), .Y(n_297) );
AND2x2_ASAP7_75t_L g313 ( .A(n_135), .B(n_199), .Y(n_313) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_135), .Y(n_348) );
AND2x2_ASAP7_75t_L g377 ( .A(n_135), .B(n_170), .Y(n_377) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_167), .Y(n_135) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_136), .A2(n_200), .B(n_207), .Y(n_199) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_136), .A2(n_213), .B(n_221), .Y(n_212) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx4_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_137), .A2(n_468), .B(n_475), .Y(n_467) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g254 ( .A(n_138), .Y(n_254) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_139), .B(n_140), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx2_ASAP7_75t_L g256 ( .A(n_144), .Y(n_256) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_145), .B(n_149), .Y(n_189) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g242 ( .A(n_146), .Y(n_242) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
INVx1_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
INVx3_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx1_ASAP7_75t_L g472 ( .A(n_148), .Y(n_472) );
INVx4_ASAP7_75t_SL g166 ( .A(n_149), .Y(n_166) );
BUFx3_ASAP7_75t_L g243 ( .A(n_149), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_153), .B(n_157), .C(n_166), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_153), .A2(n_166), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_153), .A2(n_166), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_153), .A2(n_166), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_153), .A2(n_166), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_153), .A2(n_166), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_153), .A2(n_166), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_153), .A2(n_166), .B(n_540), .C(n_541), .Y(n_539) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx3_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_158), .B(n_218), .Y(n_217) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_162), .B(n_205), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_162), .A2(n_239), .B1(n_261), .B2(n_262), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_162), .B(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_163), .A2(n_194), .B1(n_495), .B2(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g463 ( .A(n_164), .Y(n_463) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_166), .A2(n_189), .B1(n_493), .B2(n_497), .Y(n_492) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_168), .A2(n_478), .B(n_484), .Y(n_477) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_169), .B(n_198), .Y(n_197) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_169), .A2(n_223), .B(n_230), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_169), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_SL g514 ( .A(n_169), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g277 ( .A(n_170), .Y(n_277) );
BUFx3_ASAP7_75t_L g285 ( .A(n_170), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_170), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g296 ( .A(n_170), .B(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_170), .B(n_184), .Y(n_325) );
AND2x2_ASAP7_75t_L g394 ( .A(n_170), .B(n_328), .Y(n_394) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_182), .Y(n_170) );
INVx1_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
INVx2_ASAP7_75t_L g232 ( .A(n_171), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_171), .A2(n_189), .B(n_235), .C(n_236), .Y(n_234) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_171), .A2(n_538), .B(n_544), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx5_ASAP7_75t_L g239 ( .A(n_179), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_179), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_179), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g196 ( .A(n_180), .Y(n_196) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g206 ( .A(n_181), .Y(n_206) );
INVx2_ASAP7_75t_SL g288 ( .A(n_183), .Y(n_288) );
OR2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_199), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_184), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g330 ( .A(n_184), .Y(n_330) );
AND2x2_ASAP7_75t_L g341 ( .A(n_184), .B(n_297), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_184), .B(n_326), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_184), .B(n_328), .Y(n_373) );
AND2x2_ASAP7_75t_L g432 ( .A(n_184), .B(n_377), .Y(n_432) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g302 ( .A(n_185), .B(n_199), .Y(n_302) );
AND2x2_ASAP7_75t_L g312 ( .A(n_185), .B(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g334 ( .A(n_185), .Y(n_334) );
AND3x2_ASAP7_75t_L g393 ( .A(n_185), .B(n_394), .C(n_395), .Y(n_393) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_197), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_186), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_186), .B(n_524), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_186), .B(n_535), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_189), .A2(n_224), .B(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_189), .A2(n_458), .B(n_459), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_189), .A2(n_518), .B(n_519), .Y(n_517) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .C(n_196), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_193), .A2(n_196), .B(n_227), .C(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_196), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_196), .A2(n_521), .B(n_522), .Y(n_520) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
INVx1_ASAP7_75t_SL g328 ( .A(n_199), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_199), .B(n_277), .C(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_246), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_209), .A2(n_312), .B(n_364), .C(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_211), .B(n_233), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_211), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g380 ( .A(n_211), .Y(n_380) );
AND2x2_ASAP7_75t_L g401 ( .A(n_211), .B(n_248), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_211), .B(n_310), .Y(n_429) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AND2x2_ASAP7_75t_L g274 ( .A(n_212), .B(n_265), .Y(n_274) );
INVx2_ASAP7_75t_L g281 ( .A(n_212), .Y(n_281) );
AND2x2_ASAP7_75t_L g301 ( .A(n_212), .B(n_248), .Y(n_301) );
AND2x2_ASAP7_75t_L g351 ( .A(n_212), .B(n_233), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_212), .Y(n_355) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_220), .Y(n_532) );
INVx2_ASAP7_75t_SL g265 ( .A(n_222), .Y(n_265) );
BUFx2_ASAP7_75t_L g291 ( .A(n_222), .Y(n_291) );
AND2x2_ASAP7_75t_L g418 ( .A(n_222), .B(n_233), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g264 ( .A(n_232), .Y(n_264) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_232), .A2(n_527), .B(n_534), .Y(n_526) );
INVx3_ASAP7_75t_SL g248 ( .A(n_233), .Y(n_248) );
AND2x2_ASAP7_75t_L g273 ( .A(n_233), .B(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g280 ( .A(n_233), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g310 ( .A(n_233), .B(n_270), .Y(n_310) );
OR2x2_ASAP7_75t_L g319 ( .A(n_233), .B(n_265), .Y(n_319) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
AND2x2_ASAP7_75t_L g342 ( .A(n_233), .B(n_295), .Y(n_342) );
AND2x2_ASAP7_75t_L g370 ( .A(n_233), .B(n_250), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_233), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g408 ( .A(n_233), .B(n_249), .Y(n_408) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_244), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .C(n_241), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_239), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_242), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_L g332 ( .A(n_248), .B(n_281), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_248), .B(n_274), .Y(n_360) );
AND2x2_ASAP7_75t_L g378 ( .A(n_248), .B(n_295), .Y(n_378) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_265), .Y(n_249) );
AND2x2_ASAP7_75t_L g279 ( .A(n_250), .B(n_265), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_250), .B(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g317 ( .A(n_250), .Y(n_317) );
OR2x2_ASAP7_75t_L g365 ( .A(n_250), .B(n_285), .Y(n_365) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_255), .B(n_263), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_252), .A2(n_271), .B(n_272), .Y(n_270) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_252), .A2(n_517), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI21xp5_ASAP7_75t_SL g508 ( .A1(n_253), .A2(n_509), .B(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_254), .A2(n_457), .B(n_464), .Y(n_456) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_254), .A2(n_492), .B(n_498), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_254), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_263), .Y(n_272) );
AND2x2_ASAP7_75t_L g300 ( .A(n_265), .B(n_270), .Y(n_300) );
INVx1_ASAP7_75t_L g308 ( .A(n_265), .Y(n_308) );
AND2x2_ASAP7_75t_L g403 ( .A(n_265), .B(n_281), .Y(n_403) );
AOI222xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_275), .B1(n_278), .B2(n_282), .C1(n_286), .C2(n_289), .Y(n_266) );
INVx1_ASAP7_75t_L g398 ( .A(n_267), .Y(n_398) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_273), .Y(n_267) );
AND2x2_ASAP7_75t_L g294 ( .A(n_268), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g305 ( .A(n_268), .B(n_274), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_268), .B(n_296), .Y(n_321) );
OAI222xp33_ASAP7_75t_L g343 ( .A1(n_268), .A2(n_344), .B1(n_349), .B2(n_350), .C1(n_358), .C2(n_360), .Y(n_343) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g331 ( .A(n_270), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_270), .B(n_351), .Y(n_391) );
AND2x2_ASAP7_75t_L g402 ( .A(n_270), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g410 ( .A(n_273), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_275), .B(n_326), .Y(n_389) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_277), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g347 ( .A(n_277), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx3_ASAP7_75t_L g292 ( .A(n_280), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_280), .A2(n_383), .B(n_386), .C(n_388), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_280), .B(n_317), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_280), .B(n_300), .Y(n_422) );
AND2x2_ASAP7_75t_L g295 ( .A(n_281), .B(n_291), .Y(n_295) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_285), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g374 ( .A(n_285), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g413 ( .A(n_285), .B(n_313), .Y(n_413) );
INVx1_ASAP7_75t_L g425 ( .A(n_285), .Y(n_425) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_288), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g406 ( .A(n_291), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B(n_298), .C(n_302), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_294), .A2(n_324), .B1(n_339), .B2(n_342), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_295), .B(n_309), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_295), .B(n_317), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_296), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g359 ( .A(n_296), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_296), .B(n_346), .Y(n_366) );
INVx2_ASAP7_75t_L g327 ( .A(n_297), .Y(n_327) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NOR4xp25_ASAP7_75t_L g304 ( .A(n_301), .B(n_305), .C(n_306), .D(n_309), .Y(n_304) );
INVx1_ASAP7_75t_SL g375 ( .A(n_302), .Y(n_375) );
AND2x2_ASAP7_75t_L g419 ( .A(n_302), .B(n_420), .Y(n_419) );
OAI211xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_311), .B(n_314), .C(n_323), .Y(n_303) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_310), .B(n_380), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_312), .A2(n_431), .B1(n_432), .B2(n_433), .Y(n_430) );
INVx1_ASAP7_75t_SL g385 ( .A(n_313), .Y(n_385) );
AND2x2_ASAP7_75t_L g424 ( .A(n_313), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_317), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_321), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_322), .B(n_347), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_329), .B(n_331), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g399 ( .A(n_326), .Y(n_399) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g427 ( .A(n_327), .Y(n_427) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_328), .Y(n_354) );
OAI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B(n_338), .Y(n_333) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_334), .Y(n_346) );
OR2x2_ASAP7_75t_L g384 ( .A(n_334), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI21xp33_ASAP7_75t_SL g379 ( .A1(n_337), .A2(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_341), .A2(n_368), .B1(n_371), .B2(n_378), .C(n_379), .Y(n_367) );
INVx1_ASAP7_75t_SL g411 ( .A(n_342), .Y(n_411) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OR2x2_ASAP7_75t_L g358 ( .A(n_346), .B(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_355), .B2(n_356), .Y(n_350) );
INVx1_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_354), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_396), .C(n_409), .D(n_421), .Y(n_361) );
NAND3xp33_ASAP7_75t_SL g362 ( .A(n_363), .B(n_367), .C(n_382), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_365), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_372), .B(n_377), .Y(n_381) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g409 ( .A1(n_384), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_409) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_386), .A2(n_401), .B(n_402), .C(n_404), .Y(n_400) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_387), .A2(n_405), .B1(n_407), .B2(n_408), .Y(n_404) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_399), .C(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g415 ( .A(n_408), .Y(n_415) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_419), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_423), .B1(n_426), .B2(n_428), .C(n_430), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_436), .A2(n_450), .B1(n_718), .B2(n_719), .Y(n_449) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g446 ( .A(n_441), .Y(n_446) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI21xp33_ASAP7_75t_SL g447 ( .A1(n_445), .A2(n_448), .B(n_734), .Y(n_447) );
INVx1_ASAP7_75t_L g727 ( .A(n_450), .Y(n_727) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_634), .Y(n_450) );
NOR5xp2_ASAP7_75t_L g451 ( .A(n_452), .B(n_557), .C(n_589), .D(n_604), .E(n_621), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_485), .B(n_504), .C(n_545), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_466), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_454), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_454), .B(n_609), .Y(n_672) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_455), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_455), .B(n_501), .Y(n_558) );
AND2x2_ASAP7_75t_L g599 ( .A(n_455), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_455), .B(n_568), .Y(n_603) );
OR2x2_ASAP7_75t_L g640 ( .A(n_455), .B(n_491), .Y(n_640) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g490 ( .A(n_456), .B(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g548 ( .A(n_456), .Y(n_548) );
OR2x2_ASAP7_75t_L g711 ( .A(n_456), .B(n_551), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_466), .A2(n_614), .B1(n_615), .B2(n_618), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_466), .B(n_548), .Y(n_697) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
AND2x2_ASAP7_75t_L g503 ( .A(n_467), .B(n_491), .Y(n_503) );
AND2x2_ASAP7_75t_L g550 ( .A(n_467), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g555 ( .A(n_467), .Y(n_555) );
INVx3_ASAP7_75t_L g568 ( .A(n_467), .Y(n_568) );
OR2x2_ASAP7_75t_L g588 ( .A(n_467), .B(n_551), .Y(n_588) );
AND2x2_ASAP7_75t_L g607 ( .A(n_467), .B(n_477), .Y(n_607) );
BUFx2_ASAP7_75t_L g639 ( .A(n_467), .Y(n_639) );
AND2x4_ASAP7_75t_L g554 ( .A(n_476), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g489 ( .A(n_477), .Y(n_489) );
INVx2_ASAP7_75t_L g502 ( .A(n_477), .Y(n_502) );
OR2x2_ASAP7_75t_L g570 ( .A(n_477), .B(n_551), .Y(n_570) );
AND2x2_ASAP7_75t_L g600 ( .A(n_477), .B(n_491), .Y(n_600) );
AND2x2_ASAP7_75t_L g617 ( .A(n_477), .B(n_548), .Y(n_617) );
AND2x2_ASAP7_75t_L g657 ( .A(n_477), .B(n_568), .Y(n_657) );
AND2x2_ASAP7_75t_SL g693 ( .A(n_477), .B(n_503), .Y(n_693) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp33_ASAP7_75t_SL g486 ( .A(n_487), .B(n_500), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_488), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_489), .A2(n_503), .B(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_489), .B(n_491), .Y(n_687) );
AND2x2_ASAP7_75t_L g623 ( .A(n_490), .B(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_491), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_500), .B(n_548), .Y(n_716) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_501), .A2(n_659), .B1(n_660), .B2(n_665), .Y(n_658) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AND2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g587 ( .A(n_502), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g624 ( .A(n_502), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_503), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g678 ( .A(n_503), .Y(n_678) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_525), .Y(n_505) );
INVx4_ASAP7_75t_L g564 ( .A(n_506), .Y(n_564) );
AND2x2_ASAP7_75t_L g642 ( .A(n_506), .B(n_609), .Y(n_642) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
INVx3_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
AND2x2_ASAP7_75t_L g575 ( .A(n_507), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g579 ( .A(n_507), .Y(n_579) );
INVx2_ASAP7_75t_L g593 ( .A(n_507), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_507), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g650 ( .A(n_507), .B(n_645), .Y(n_650) );
AND2x2_ASAP7_75t_L g715 ( .A(n_507), .B(n_685), .Y(n_715) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
AND2x2_ASAP7_75t_L g556 ( .A(n_516), .B(n_537), .Y(n_556) );
INVx2_ASAP7_75t_L g576 ( .A(n_516), .Y(n_576) );
INVx1_ASAP7_75t_L g581 ( .A(n_525), .Y(n_581) );
AND2x2_ASAP7_75t_L g627 ( .A(n_525), .B(n_575), .Y(n_627) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_536), .Y(n_525) );
INVx2_ASAP7_75t_L g566 ( .A(n_526), .Y(n_566) );
INVx1_ASAP7_75t_L g574 ( .A(n_526), .Y(n_574) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_526), .B(n_576), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
AND2x2_ASAP7_75t_L g609 ( .A(n_536), .B(n_566), .Y(n_609) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g562 ( .A(n_537), .Y(n_562) );
AND2x2_ASAP7_75t_L g645 ( .A(n_537), .B(n_576), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_552), .B(n_556), .Y(n_545) );
INVx1_ASAP7_75t_SL g590 ( .A(n_546), .Y(n_590) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_547), .B(n_554), .Y(n_647) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g596 ( .A(n_548), .B(n_551), .Y(n_596) );
AND2x2_ASAP7_75t_L g625 ( .A(n_548), .B(n_569), .Y(n_625) );
OR2x2_ASAP7_75t_L g628 ( .A(n_548), .B(n_588), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_549), .A2(n_641), .B1(n_693), .B2(n_694), .C1(n_696), .C2(n_698), .Y(n_692) );
BUFx2_ASAP7_75t_L g606 ( .A(n_551), .Y(n_606) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g595 ( .A(n_554), .B(n_596), .Y(n_595) );
INVx3_ASAP7_75t_SL g612 ( .A(n_554), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_554), .B(n_606), .Y(n_666) );
AND2x2_ASAP7_75t_L g601 ( .A(n_556), .B(n_561), .Y(n_601) );
INVx1_ASAP7_75t_L g620 ( .A(n_556), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_559), .B1(n_563), .B2(n_567), .C(n_571), .Y(n_557) );
OR2x2_ASAP7_75t_L g629 ( .A(n_559), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g614 ( .A(n_561), .B(n_584), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_561), .B(n_574), .Y(n_654) );
AND2x2_ASAP7_75t_L g659 ( .A(n_561), .B(n_609), .Y(n_659) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_561), .Y(n_669) );
NAND2x1_ASAP7_75t_SL g680 ( .A(n_561), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g565 ( .A(n_562), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g585 ( .A(n_562), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_562), .B(n_580), .Y(n_611) );
INVx1_ASAP7_75t_L g677 ( .A(n_562), .Y(n_677) );
INVx1_ASAP7_75t_L g652 ( .A(n_563), .Y(n_652) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g664 ( .A(n_564), .Y(n_664) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_564), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g681 ( .A(n_565), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_565), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g584 ( .A(n_566), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_566), .B(n_576), .Y(n_597) );
INVx1_ASAP7_75t_L g663 ( .A(n_566), .Y(n_663) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI21xp5_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_577), .B(n_586), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g717 ( .A(n_573), .B(n_650), .Y(n_717) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g685 ( .A(n_574), .B(n_645), .Y(n_685) );
AOI32xp33_ASAP7_75t_L g598 ( .A1(n_575), .A2(n_581), .A3(n_599), .B1(n_601), .B2(n_602), .Y(n_598) );
AOI322xp5_ASAP7_75t_L g700 ( .A1(n_575), .A2(n_607), .A3(n_690), .B1(n_701), .B2(n_702), .C1(n_703), .C2(n_705), .Y(n_700) );
INVx2_ASAP7_75t_L g580 ( .A(n_576), .Y(n_580) );
INVx1_ASAP7_75t_L g690 ( .A(n_576), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_578), .B(n_584), .Y(n_633) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_579), .B(n_645), .Y(n_695) );
INVx1_ASAP7_75t_L g582 ( .A(n_580), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_580), .B(n_609), .Y(n_699) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_588), .B(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_591), .B1(n_594), .B2(n_597), .C(n_598), .Y(n_589) );
OR2x2_ASAP7_75t_L g610 ( .A(n_591), .B(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g619 ( .A(n_591), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g644 ( .A(n_592), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g648 ( .A(n_602), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_608), .B1(n_610), .B2(n_612), .C(n_613), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_606), .A2(n_637), .B1(n_641), .B2(n_642), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_607), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g712 ( .A(n_607), .Y(n_712) );
INVx1_ASAP7_75t_L g706 ( .A(n_609), .Y(n_706) );
INVx1_ASAP7_75t_SL g641 ( .A(n_610), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_612), .B(n_640), .Y(n_702) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_617), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g683 ( .A(n_617), .Y(n_683) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_626), .B1(n_628), .B2(n_629), .C(n_631), .Y(n_621) );
NOR2xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_623), .A2(n_641), .B1(n_687), .B2(n_688), .Y(n_686) );
CKINVDCx14_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_628), .A2(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_667), .C(n_691), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_636), .B(n_643), .C(n_651), .D(n_658), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g714 ( .A(n_639), .Y(n_714) );
INVx3_ASAP7_75t_SL g708 ( .A(n_640), .Y(n_708) );
OR2x2_ASAP7_75t_L g713 ( .A(n_640), .B(n_714), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B1(n_648), .B2(n_650), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_645), .B(n_663), .Y(n_704) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_655), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_670), .B(n_673), .C(n_686), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g701 ( .A(n_672), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_678), .B1(n_679), .B2(n_682), .C1(n_684), .C2(n_685), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND4xp25_ASAP7_75t_SL g710 ( .A(n_683), .B(n_711), .C(n_712), .D(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_700), .C(n_709), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_709) );
INVx1_ASAP7_75t_L g729 ( .A(n_719), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_720), .Y(n_730) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
endmodule