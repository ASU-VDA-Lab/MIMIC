module real_aes_7341_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g103 ( .A(n_0), .Y(n_103) );
INVx1_ASAP7_75t_L g478 ( .A(n_1), .Y(n_478) );
INVx1_ASAP7_75t_L g192 ( .A(n_2), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_3), .A2(n_37), .B1(n_153), .B2(n_508), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g160 ( .A1(n_4), .A2(n_134), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_5), .B(n_127), .Y(n_491) );
AND2x6_ASAP7_75t_L g139 ( .A(n_6), .B(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_7), .A2(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_8), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_8), .B(n_38), .Y(n_448) );
INVx1_ASAP7_75t_L g167 ( .A(n_9), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_10), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g132 ( .A(n_11), .Y(n_132) );
INVx1_ASAP7_75t_L g472 ( .A(n_12), .Y(n_472) );
INVx1_ASAP7_75t_L g248 ( .A(n_13), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_14), .B(n_175), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_15), .B(n_128), .Y(n_549) );
AO32x2_ASAP7_75t_L g521 ( .A1(n_16), .A2(n_127), .A3(n_172), .B1(n_500), .B2(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_17), .A2(n_117), .B1(n_118), .B2(n_443), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_17), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_18), .B(n_153), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_19), .B(n_148), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_20), .B(n_128), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_21), .A2(n_49), .B1(n_153), .B2(n_508), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_22), .B(n_134), .Y(n_204) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_23), .A2(n_75), .B1(n_153), .B2(n_175), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_24), .B(n_153), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_25), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_26), .A2(n_246), .B(n_247), .C(n_249), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_27), .Y(n_451) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_28), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_29), .B(n_169), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_30), .B(n_165), .Y(n_194) );
INVx1_ASAP7_75t_L g181 ( .A(n_31), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_32), .B(n_169), .Y(n_538) );
INVx2_ASAP7_75t_L g137 ( .A(n_33), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_34), .B(n_153), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_35), .B(n_169), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_36), .A2(n_139), .B(n_143), .C(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g109 ( .A(n_38), .Y(n_109) );
INVx1_ASAP7_75t_L g179 ( .A(n_39), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_40), .B(n_165), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_41), .B(n_153), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_42), .A2(n_85), .B1(n_211), .B2(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_43), .B(n_153), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_44), .B(n_153), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_45), .Y(n_182) );
OAI222xp33_ASAP7_75t_L g453 ( .A1(n_46), .A2(n_454), .B1(n_751), .B2(n_752), .C1(n_757), .C2(n_761), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g751 ( .A(n_46), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_47), .B(n_477), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_48), .B(n_134), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_50), .A2(n_59), .B1(n_153), .B2(n_175), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_51), .A2(n_143), .B1(n_175), .B2(n_177), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_52), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_53), .B(n_153), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_54), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_55), .B(n_153), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_56), .A2(n_152), .B(n_164), .C(n_166), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_57), .Y(n_224) );
INVx1_ASAP7_75t_L g162 ( .A(n_58), .Y(n_162) );
INVx1_ASAP7_75t_L g140 ( .A(n_60), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_61), .B(n_153), .Y(n_479) );
INVx1_ASAP7_75t_L g131 ( .A(n_62), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_63), .Y(n_114) );
AO32x2_ASAP7_75t_L g505 ( .A1(n_64), .A2(n_127), .A3(n_228), .B1(n_500), .B2(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g498 ( .A(n_65), .Y(n_498) );
INVx1_ASAP7_75t_L g533 ( .A(n_66), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_67), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_SL g147 ( .A1(n_68), .A2(n_148), .B(n_149), .C(n_152), .Y(n_147) );
INVxp67_ASAP7_75t_L g150 ( .A(n_69), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_70), .B(n_175), .Y(n_534) );
INVx1_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_72), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_73), .A2(n_100), .B1(n_110), .B2(n_764), .Y(n_99) );
INVx1_ASAP7_75t_L g217 ( .A(n_74), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_76), .A2(n_139), .B(n_143), .C(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_77), .B(n_508), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_78), .B(n_175), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_79), .B(n_193), .Y(n_207) );
INVx2_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_81), .B(n_148), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_82), .B(n_175), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_83), .A2(n_139), .B(n_143), .C(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g104 ( .A(n_84), .Y(n_104) );
OR2x2_ASAP7_75t_L g445 ( .A(n_84), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g456 ( .A(n_84), .B(n_447), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_86), .A2(n_98), .B1(n_175), .B2(n_176), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_87), .B(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_88), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_89), .A2(n_139), .B(n_143), .C(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_90), .Y(n_238) );
INVx1_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_92), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_93), .B(n_193), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_94), .B(n_175), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_95), .B(n_127), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_96), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_97), .A2(n_134), .B(n_141), .Y(n_133) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g765 ( .A(n_101), .Y(n_765) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_108), .Y(n_101) );
NAND3xp33_ASAP7_75t_SL g102 ( .A(n_103), .B(n_104), .C(n_105), .Y(n_102) );
AND2x2_ASAP7_75t_L g447 ( .A(n_103), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g459 ( .A(n_104), .B(n_447), .Y(n_459) );
NOR2x2_ASAP7_75t_L g760 ( .A(n_104), .B(n_446), .Y(n_760) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_115), .B(n_452), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g763 ( .A(n_113), .Y(n_763) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_444), .B(n_449), .Y(n_115) );
INVx2_ASAP7_75t_L g443 ( .A(n_118), .Y(n_443) );
INVx1_ASAP7_75t_SL g457 ( .A(n_118), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_118), .A2(n_753), .B1(n_755), .B2(n_756), .Y(n_752) );
INVx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND4x1_ASAP7_75t_L g119 ( .A(n_120), .B(n_361), .C(n_408), .D(n_428), .Y(n_119) );
NOR3xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_291), .C(n_316), .Y(n_120) );
OAI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_199), .B(n_251), .C(n_281), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_170), .Y(n_123) );
INVx3_ASAP7_75t_SL g333 ( .A(n_124), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_124), .B(n_264), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_124), .B(n_186), .Y(n_414) );
AND2x2_ASAP7_75t_L g437 ( .A(n_124), .B(n_303), .Y(n_437) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_158), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g255 ( .A(n_126), .B(n_159), .Y(n_255) );
INVx3_ASAP7_75t_L g268 ( .A(n_126), .Y(n_268) );
AND2x2_ASAP7_75t_L g273 ( .A(n_126), .B(n_158), .Y(n_273) );
OR2x2_ASAP7_75t_L g324 ( .A(n_126), .B(n_265), .Y(n_324) );
BUFx2_ASAP7_75t_L g344 ( .A(n_126), .Y(n_344) );
AND2x2_ASAP7_75t_L g354 ( .A(n_126), .B(n_265), .Y(n_354) );
AND2x2_ASAP7_75t_L g360 ( .A(n_126), .B(n_171), .Y(n_360) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_133), .B(n_155), .Y(n_126) );
INVx4_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_127), .A2(n_484), .B(n_491), .Y(n_483) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_129), .B(n_130), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
BUFx2_ASAP7_75t_L g242 ( .A(n_134), .Y(n_242) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_135), .B(n_139), .Y(n_183) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g477 ( .A(n_136), .Y(n_477) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
INVx1_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
INVx1_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx1_ASAP7_75t_L g148 ( .A(n_138), .Y(n_148) );
INVx3_ASAP7_75t_L g151 ( .A(n_138), .Y(n_151) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
INVx4_ASAP7_75t_SL g154 ( .A(n_139), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_139), .A2(n_471), .B(n_475), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_139), .A2(n_485), .B(n_488), .Y(n_484) );
BUFx3_ASAP7_75t_L g500 ( .A(n_139), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_139), .A2(n_513), .B(n_517), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_139), .A2(n_532), .B(n_535), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_147), .C(n_154), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_142), .A2(n_154), .B(n_162), .C(n_163), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_142), .A2(n_154), .B(n_244), .C(n_245), .Y(n_243) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
BUFx3_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
INVx1_ASAP7_75t_L g508 ( .A(n_144), .Y(n_508) );
INVx1_ASAP7_75t_L g516 ( .A(n_148), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_151), .B(n_167), .Y(n_166) );
INVx5_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g506 ( .A1(n_151), .A2(n_165), .B1(n_507), .B2(n_509), .Y(n_506) );
O2A1O1Ixp5_ASAP7_75t_SL g532 ( .A1(n_152), .A2(n_193), .B(n_533), .C(n_534), .Y(n_532) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_153), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_154), .A2(n_174), .B1(n_182), .B2(n_183), .Y(n_173) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_156), .A2(n_160), .B(n_168), .Y(n_159) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_157), .B(n_214), .Y(n_213) );
AO21x1_ASAP7_75t_L g544 ( .A1(n_157), .A2(n_545), .B(n_548), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_157), .B(n_500), .C(n_545), .Y(n_563) );
INVx1_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_159), .B(n_265), .Y(n_279) );
INVx2_ASAP7_75t_L g289 ( .A(n_159), .Y(n_289) );
AND2x2_ASAP7_75t_L g302 ( .A(n_159), .B(n_268), .Y(n_302) );
OR2x2_ASAP7_75t_L g313 ( .A(n_159), .B(n_265), .Y(n_313) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_159), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g371 ( .A(n_159), .Y(n_371) );
AND2x2_ASAP7_75t_L g417 ( .A(n_159), .B(n_171), .Y(n_417) );
O2A1O1Ixp5_ASAP7_75t_L g497 ( .A1(n_164), .A2(n_476), .B(n_498), .C(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_164), .A2(n_518), .B(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx4_ASAP7_75t_L g234 ( .A(n_165), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_165), .A2(n_480), .B1(n_523), .B2(n_524), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_165), .A2(n_480), .B1(n_546), .B2(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g198 ( .A(n_169), .Y(n_198) );
INVx2_ASAP7_75t_L g228 ( .A(n_169), .Y(n_228) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_169), .A2(n_241), .B(n_250), .Y(n_240) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_169), .A2(n_512), .B(n_520), .Y(n_511) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_169), .A2(n_531), .B(n_538), .Y(n_530) );
INVx3_ASAP7_75t_SL g290 ( .A(n_170), .Y(n_290) );
OR2x2_ASAP7_75t_L g343 ( .A(n_170), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_186), .Y(n_170) );
INVx3_ASAP7_75t_L g265 ( .A(n_171), .Y(n_265) );
AND2x2_ASAP7_75t_L g332 ( .A(n_171), .B(n_187), .Y(n_332) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_171), .Y(n_400) );
AOI33xp33_ASAP7_75t_L g404 ( .A1(n_171), .A2(n_333), .A3(n_340), .B1(n_349), .B2(n_405), .B3(n_406), .Y(n_404) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_184), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_172), .B(n_185), .Y(n_184) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_172), .A2(n_188), .B(n_196), .Y(n_187) );
INVx2_ASAP7_75t_L g212 ( .A(n_172), .Y(n_212) );
INVx2_ASAP7_75t_L g195 ( .A(n_175), .Y(n_195) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_177) );
INVx2_ASAP7_75t_L g180 ( .A(n_178), .Y(n_180) );
INVx4_ASAP7_75t_L g246 ( .A(n_178), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_183), .A2(n_189), .B(n_190), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_183), .A2(n_217), .B(n_218), .Y(n_216) );
INVx1_ASAP7_75t_L g253 ( .A(n_186), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_186), .B(n_268), .Y(n_267) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_186), .B(n_328), .C(n_330), .Y(n_327) );
AND2x2_ASAP7_75t_L g353 ( .A(n_186), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_186), .B(n_360), .Y(n_363) );
AND2x2_ASAP7_75t_L g416 ( .A(n_186), .B(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx3_ASAP7_75t_L g272 ( .A(n_187), .Y(n_272) );
OR2x2_ASAP7_75t_L g366 ( .A(n_187), .B(n_265), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .C(n_195), .Y(n_191) );
INVx2_ASAP7_75t_L g480 ( .A(n_193), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_193), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_193), .A2(n_495), .B(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_195), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_198), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_198), .B(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_225), .Y(n_199) );
AOI32xp33_ASAP7_75t_L g317 ( .A1(n_200), .A2(n_318), .A3(n_320), .B1(n_322), .B2(n_325), .Y(n_317) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_200), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g420 ( .A(n_200), .Y(n_420) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g352 ( .A(n_201), .B(n_336), .Y(n_352) );
AND2x2_ASAP7_75t_L g372 ( .A(n_201), .B(n_298), .Y(n_372) );
AND2x2_ASAP7_75t_L g440 ( .A(n_201), .B(n_358), .Y(n_440) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_215), .Y(n_201) );
INVx3_ASAP7_75t_L g261 ( .A(n_202), .Y(n_261) );
AND2x2_ASAP7_75t_L g275 ( .A(n_202), .B(n_259), .Y(n_275) );
OR2x2_ASAP7_75t_L g280 ( .A(n_202), .B(n_258), .Y(n_280) );
INVx1_ASAP7_75t_L g287 ( .A(n_202), .Y(n_287) );
AND2x2_ASAP7_75t_L g295 ( .A(n_202), .B(n_269), .Y(n_295) );
AND2x2_ASAP7_75t_L g297 ( .A(n_202), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_202), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g350 ( .A(n_202), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_202), .B(n_435), .Y(n_434) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
AOI21xp5_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_205), .B(n_212), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_209), .A2(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
INVx1_ASAP7_75t_L g222 ( .A(n_212), .Y(n_222) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_212), .A2(n_470), .B(n_481), .Y(n_469) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_212), .A2(n_493), .B(n_501), .Y(n_492) );
INVx2_ASAP7_75t_L g259 ( .A(n_215), .Y(n_259) );
AND2x2_ASAP7_75t_L g305 ( .A(n_215), .B(n_226), .Y(n_305) );
AND2x2_ASAP7_75t_L g315 ( .A(n_215), .B(n_240), .Y(n_315) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_222), .B(n_223), .Y(n_215) );
INVx2_ASAP7_75t_L g435 ( .A(n_225), .Y(n_435) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_226), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g276 ( .A(n_226), .Y(n_276) );
AND2x2_ASAP7_75t_L g320 ( .A(n_226), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g336 ( .A(n_226), .B(n_299), .Y(n_336) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g284 ( .A(n_227), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_227), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g349 ( .A(n_227), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_227), .B(n_259), .Y(n_381) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_235), .Y(n_231) );
AND2x2_ASAP7_75t_L g260 ( .A(n_239), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g321 ( .A(n_239), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_239), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g358 ( .A(n_239), .Y(n_358) );
INVx1_ASAP7_75t_L g391 ( .A(n_239), .Y(n_391) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g269 ( .A(n_240), .B(n_259), .Y(n_269) );
INVx1_ASAP7_75t_L g299 ( .A(n_240), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_246), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g474 ( .A(n_246), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_246), .A2(n_536), .B(n_537), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_256), .B1(n_262), .B2(n_269), .C(n_270), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_253), .B(n_273), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_253), .B(n_336), .Y(n_413) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_255), .B(n_303), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_255), .B(n_264), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_255), .B(n_278), .Y(n_407) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g329 ( .A(n_259), .Y(n_329) );
AND2x2_ASAP7_75t_L g304 ( .A(n_260), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g382 ( .A(n_260), .Y(n_382) );
AND2x2_ASAP7_75t_L g314 ( .A(n_261), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_261), .B(n_284), .Y(n_330) );
AND2x2_ASAP7_75t_L g394 ( .A(n_261), .B(n_320), .Y(n_394) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g303 ( .A(n_265), .B(n_272), .Y(n_303) );
AND2x2_ASAP7_75t_L g399 ( .A(n_266), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_268), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_269), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_269), .B(n_276), .Y(n_364) );
AND2x2_ASAP7_75t_L g384 ( .A(n_269), .B(n_284), .Y(n_384) );
AND2x2_ASAP7_75t_L g405 ( .A(n_269), .B(n_349), .Y(n_405) );
OAI32xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .A3(n_276), .B1(n_277), .B2(n_280), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_SL g278 ( .A(n_272), .Y(n_278) );
NAND2x1_ASAP7_75t_L g319 ( .A(n_272), .B(n_302), .Y(n_319) );
OR2x2_ASAP7_75t_L g323 ( .A(n_272), .B(n_324), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_272), .B(n_371), .Y(n_424) );
INVx1_ASAP7_75t_L g292 ( .A(n_273), .Y(n_292) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_274), .A2(n_365), .B1(n_411), .B2(n_414), .C(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g282 ( .A(n_275), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g325 ( .A(n_275), .B(n_298), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_275), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g403 ( .A(n_275), .B(n_336), .Y(n_403) );
INVxp67_ASAP7_75t_L g339 ( .A(n_276), .Y(n_339) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g409 ( .A(n_278), .B(n_396), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_278), .B(n_359), .Y(n_432) );
INVx1_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_280), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g425 ( .A(n_280), .B(n_426), .Y(n_425) );
OAI21xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_285), .B(n_288), .Y(n_281) );
AND2x2_ASAP7_75t_L g294 ( .A(n_283), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g378 ( .A(n_287), .B(n_298), .Y(n_378) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g396 ( .A(n_289), .B(n_354), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_289), .B(n_353), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_290), .B(n_302), .Y(n_376) );
OAI211xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_296), .C(n_306), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_292), .A2(n_327), .B1(n_331), .B2(n_334), .C(n_337), .Y(n_326) );
AOI31xp33_ASAP7_75t_L g421 ( .A1(n_292), .A2(n_422), .A3(n_423), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .B1(n_302), .B2(n_304), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g422 ( .A(n_302), .Y(n_422) );
INVx1_ASAP7_75t_L g385 ( .A(n_303), .Y(n_385) );
O2A1O1Ixp33_ASAP7_75t_L g428 ( .A1(n_305), .A2(n_429), .B(n_431), .C(n_433), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_310), .B2(n_314), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_311), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_313), .A2(n_347), .B1(n_366), .B2(n_402), .C(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g397 ( .A(n_314), .Y(n_397) );
INVx1_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
NAND3xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_326), .C(n_341), .Y(n_316) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_318), .A2(n_368), .B(n_372), .Y(n_367) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_320), .B(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g427 ( .A(n_321), .Y(n_427) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g365 ( .A(n_328), .B(n_348), .Y(n_365) );
INVx1_ASAP7_75t_L g340 ( .A(n_329), .Y(n_340) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g338 ( .A(n_332), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_332), .B(n_370), .Y(n_369) );
NOR4xp25_ASAP7_75t_L g337 ( .A(n_333), .B(n_338), .C(n_339), .D(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI222xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_346), .B1(n_352), .B2(n_353), .C1(n_355), .C2(n_359), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g439 ( .A(n_343), .Y(n_439) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_355), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_360), .A2(n_416), .B(n_418), .Y(n_415) );
NOR4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_373), .C(n_386), .D(n_401), .Y(n_361) );
OAI221xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_364), .B1(n_365), .B2(n_366), .C(n_367), .Y(n_362) );
INVx1_ASAP7_75t_L g442 ( .A(n_363), .Y(n_442) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_370), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OAI222xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_379), .B2(n_380), .C1(n_383), .C2(n_385), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI211xp5_ASAP7_75t_L g408 ( .A1(n_378), .A2(n_409), .B(n_410), .C(n_421), .Y(n_408) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
OAI222xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_392), .B1(n_393), .B2(n_395), .C1(n_397), .C2(n_398), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_403), .A2(n_406), .B1(n_439), .B2(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_436), .B(n_438), .C(n_441), .Y(n_433) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_445), .Y(n_450) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g452 ( .A1(n_449), .A2(n_453), .B(n_762), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_457), .B1(n_458), .B2(n_460), .Y(n_454) );
INVx2_ASAP7_75t_L g754 ( .A(n_455), .Y(n_754) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx6_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g755 ( .A(n_459), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_460), .Y(n_756) );
AND2x2_ASAP7_75t_SL g460 ( .A(n_461), .B(n_717), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_621), .C(n_705), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_564), .C(n_586), .D(n_602), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_502), .B1(n_525), .B2(n_543), .C(n_550), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_482), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_466), .B(n_543), .Y(n_576) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_466), .B(n_604), .C(n_617), .D(n_619), .Y(n_616) );
INVxp67_ASAP7_75t_L g733 ( .A(n_466), .Y(n_733) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g615 ( .A(n_467), .B(n_553), .Y(n_615) );
AND2x2_ASAP7_75t_L g639 ( .A(n_467), .B(n_482), .Y(n_639) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g606 ( .A(n_468), .B(n_542), .Y(n_606) );
AND2x2_ASAP7_75t_L g646 ( .A(n_468), .B(n_627), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_468), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_468), .B(n_483), .Y(n_687) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g541 ( .A(n_469), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g558 ( .A(n_469), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g570 ( .A(n_469), .B(n_483), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_469), .B(n_492), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_478), .B(n_479), .C(n_480), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_480), .A2(n_489), .B(n_490), .Y(n_488) );
AND2x2_ASAP7_75t_L g573 ( .A(n_482), .B(n_574), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_482), .A2(n_623), .B1(n_626), .B2(n_628), .C(n_632), .Y(n_622) );
AND2x2_ASAP7_75t_L g681 ( .A(n_482), .B(n_646), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_482), .B(n_663), .Y(n_715) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
INVx3_ASAP7_75t_L g542 ( .A(n_483), .Y(n_542) );
AND2x2_ASAP7_75t_L g590 ( .A(n_483), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g644 ( .A(n_483), .B(n_559), .Y(n_644) );
AND2x2_ASAP7_75t_L g702 ( .A(n_483), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g543 ( .A(n_492), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g614 ( .A(n_492), .Y(n_614) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_492), .Y(n_620) );
AND2x2_ASAP7_75t_L g665 ( .A(n_492), .B(n_542), .Y(n_665) );
OR2x2_ASAP7_75t_L g704 ( .A(n_492), .B(n_544), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_497), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_502), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
AND2x2_ASAP7_75t_L g700 ( .A(n_503), .B(n_697), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_503), .B(n_682), .Y(n_732) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g631 ( .A(n_504), .B(n_555), .Y(n_631) );
AND2x2_ASAP7_75t_L g680 ( .A(n_504), .B(n_528), .Y(n_680) );
INVx1_ASAP7_75t_L g726 ( .A(n_504), .Y(n_726) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_505), .Y(n_540) );
AND2x2_ASAP7_75t_L g581 ( .A(n_505), .B(n_555), .Y(n_581) );
INVx1_ASAP7_75t_L g598 ( .A(n_505), .Y(n_598) );
AND2x2_ASAP7_75t_L g604 ( .A(n_505), .B(n_521), .Y(n_604) );
AND2x2_ASAP7_75t_L g672 ( .A(n_510), .B(n_580), .Y(n_672) );
INVx2_ASAP7_75t_L g737 ( .A(n_510), .Y(n_737) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
AND2x2_ASAP7_75t_L g554 ( .A(n_511), .B(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g567 ( .A(n_511), .B(n_529), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_511), .B(n_528), .Y(n_595) );
INVx1_ASAP7_75t_L g601 ( .A(n_511), .Y(n_601) );
INVx1_ASAP7_75t_L g618 ( .A(n_511), .Y(n_618) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_511), .Y(n_630) );
INVx2_ASAP7_75t_L g698 ( .A(n_511), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g555 ( .A(n_521), .Y(n_555) );
BUFx2_ASAP7_75t_L g652 ( .A(n_521), .Y(n_652) );
AND2x2_ASAP7_75t_L g697 ( .A(n_521), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_539), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_527), .B(n_634), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_527), .A2(n_696), .B(n_710), .Y(n_720) );
AND2x2_ASAP7_75t_L g745 ( .A(n_527), .B(n_631), .Y(n_745) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g667 ( .A(n_529), .Y(n_667) );
AND2x2_ASAP7_75t_L g696 ( .A(n_529), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_530), .Y(n_580) );
INVx2_ASAP7_75t_L g599 ( .A(n_530), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g553 ( .A(n_540), .Y(n_553) );
OR2x2_ASAP7_75t_L g566 ( .A(n_540), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g634 ( .A(n_540), .B(n_630), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_540), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g735 ( .A(n_540), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_540), .B(n_672), .Y(n_747) );
AND2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g649 ( .A(n_541), .B(n_543), .Y(n_649) );
INVx2_ASAP7_75t_L g561 ( .A(n_542), .Y(n_561) );
AND2x2_ASAP7_75t_L g589 ( .A(n_542), .B(n_562), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_542), .B(n_614), .Y(n_670) );
AND2x2_ASAP7_75t_L g584 ( .A(n_543), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g731 ( .A(n_543), .Y(n_731) );
AND2x2_ASAP7_75t_L g743 ( .A(n_543), .B(n_606), .Y(n_743) );
AND2x2_ASAP7_75t_L g569 ( .A(n_544), .B(n_559), .Y(n_569) );
INVx1_ASAP7_75t_L g664 ( .A(n_544), .Y(n_664) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g562 ( .A(n_549), .B(n_563), .Y(n_562) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_553), .B(n_600), .Y(n_609) );
OR2x2_ASAP7_75t_L g741 ( .A(n_553), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g658 ( .A(n_554), .B(n_599), .Y(n_658) );
AND2x2_ASAP7_75t_L g666 ( .A(n_554), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g725 ( .A(n_554), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g749 ( .A(n_554), .B(n_596), .Y(n_749) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_555), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g736 ( .A(n_555), .B(n_599), .Y(n_736) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
AND2x2_ASAP7_75t_L g588 ( .A(n_558), .B(n_589), .Y(n_588) );
INVxp67_ASAP7_75t_L g750 ( .A(n_558), .Y(n_750) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g585 ( .A(n_561), .Y(n_585) );
AND2x2_ASAP7_75t_L g636 ( .A(n_561), .B(n_569), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_561), .B(n_704), .Y(n_730) );
INVx2_ASAP7_75t_L g575 ( .A(n_562), .Y(n_575) );
INVx3_ASAP7_75t_L g627 ( .A(n_562), .Y(n_627) );
OR2x2_ASAP7_75t_L g655 ( .A(n_562), .B(n_656), .Y(n_655) );
AOI311xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .A3(n_570), .B(n_571), .C(n_582), .Y(n_564) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_565), .A2(n_603), .B(n_605), .C(n_607), .Y(n_602) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g587 ( .A(n_567), .Y(n_587) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g605 ( .A(n_569), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_569), .B(n_585), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_569), .B(n_570), .Y(n_738) );
AND2x2_ASAP7_75t_L g660 ( .A(n_570), .B(n_574), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g718 ( .A(n_574), .B(n_606), .Y(n_718) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_575), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g603 ( .A(n_579), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g648 ( .A(n_581), .Y(n_648) );
AND2x4_ASAP7_75t_L g710 ( .A(n_581), .B(n_679), .Y(n_710) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_584), .A2(n_650), .B1(n_662), .B2(n_666), .C1(n_668), .C2(n_672), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_590), .C(n_593), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_587), .B(n_631), .Y(n_654) );
INVx1_ASAP7_75t_L g676 ( .A(n_589), .Y(n_676) );
INVx1_ASAP7_75t_L g610 ( .A(n_591), .Y(n_610) );
OR2x2_ASAP7_75t_L g675 ( .A(n_592), .B(n_676), .Y(n_675) );
OAI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B(n_600), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_594), .B(n_612), .C(n_613), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_594), .A2(n_631), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_598), .Y(n_651) );
AND2x2_ASAP7_75t_SL g617 ( .A(n_599), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g708 ( .A(n_599), .Y(n_708) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_599), .Y(n_724) );
INVx2_ASAP7_75t_L g682 ( .A(n_600), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_604), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g656 ( .A(n_606), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_611), .B2(n_615), .C(n_616), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_610), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g744 ( .A(n_610), .Y(n_744) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g625 ( .A(n_617), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_617), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g683 ( .A(n_617), .B(n_631), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_617), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g716 ( .A(n_617), .B(n_651), .Y(n_716) );
BUFx3_ASAP7_75t_L g679 ( .A(n_618), .Y(n_679) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND5xp2_ASAP7_75t_L g621 ( .A(n_622), .B(n_640), .C(n_661), .D(n_673), .E(n_688), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g713 ( .A1(n_625), .A2(n_652), .A3(n_668), .B1(n_714), .B2(n_716), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_627), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g637 ( .A(n_631), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B1(n_637), .B2(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_647), .B1(n_649), .B2(n_650), .C(n_653), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g712 ( .A(n_644), .B(n_663), .Y(n_712) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_649), .A2(n_710), .B1(n_728), .B2(n_733), .C(n_734), .Y(n_727) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx2_ASAP7_75t_L g693 ( .A(n_652), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_657), .B2(n_659), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g671 ( .A(n_663), .Y(n_671) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B1(n_681), .B2(n_682), .C1(n_683), .C2(n_684), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_682), .A2(n_729), .B1(n_731), .B2(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_694), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_699), .B(n_701), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g742 ( .A(n_697), .Y(n_742) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_711), .C(n_713), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI211xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B(n_721), .C(n_746), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g722 ( .A(n_718), .Y(n_722) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_727), .C(n_739), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B(n_738), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
endmodule