module fake_jpeg_5254_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_27),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_63),
.B1(n_64),
.B2(n_29),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_28),
.B1(n_22),
.B2(n_20),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_68),
.B1(n_24),
.B2(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_36),
.B1(n_24),
.B2(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_33),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_42),
.B1(n_28),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_79),
.Y(n_106)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_93),
.Y(n_110)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_94),
.B1(n_52),
.B2(n_63),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_39),
.B(n_38),
.C(n_23),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_92),
.B(n_67),
.C(n_52),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_23),
.B(n_39),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_87),
.C(n_93),
.Y(n_101)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_28),
.B(n_39),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_28),
.B1(n_39),
.B2(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_74),
.B1(n_88),
.B2(n_84),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_103),
.B(n_113),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_69),
.B1(n_55),
.B2(n_56),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_75),
.B1(n_95),
.B2(n_83),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_65),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_54),
.B1(n_47),
.B2(n_60),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_118),
.B1(n_94),
.B2(n_88),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_66),
.B1(n_22),
.B2(n_38),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_119),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_65),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_80),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_130),
.B1(n_100),
.B2(n_99),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_139),
.B1(n_141),
.B2(n_146),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_85),
.B1(n_74),
.B2(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_90),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_40),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_108),
.B(n_1),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_144),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_71),
.C(n_73),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_99),
.C(n_116),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_148),
.B1(n_81),
.B2(n_89),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_80),
.B1(n_64),
.B2(n_71),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_80),
.B(n_96),
.C(n_65),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_33),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_118),
.B1(n_114),
.B2(n_122),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_145),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_104),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_105),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_51),
.B1(n_47),
.B2(n_45),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_81),
.B1(n_75),
.B2(n_51),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_75),
.B1(n_66),
.B2(n_28),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_150),
.B1(n_123),
.B2(n_98),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_46),
.B1(n_30),
.B2(n_44),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_176),
.C(n_178),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_162),
.B1(n_128),
.B2(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_103),
.B(n_119),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_163),
.B(n_167),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_165),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_107),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_177),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_120),
.B1(n_112),
.B2(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_173),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_108),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_137),
.B(n_130),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_174),
.B1(n_179),
.B2(n_128),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_139),
.B1(n_140),
.B2(n_132),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_37),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_124),
.A2(n_98),
.B1(n_121),
.B2(n_29),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_180),
.B(n_183),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_126),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_184),
.C(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_126),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_166),
.CI(n_154),
.CON(n_215),
.SN(n_215)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_200),
.B1(n_202),
.B2(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_89),
.B1(n_111),
.B2(n_151),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_40),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_162),
.A2(n_111),
.B1(n_44),
.B2(n_59),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_177),
.B1(n_175),
.B2(n_168),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_158),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_166),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_214),
.B(n_215),
.Y(n_245)
);

AO22x2_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_167),
.B1(n_164),
.B2(n_173),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_185),
.B1(n_183),
.B2(n_188),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_179),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_231),
.B1(n_206),
.B2(n_189),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_157),
.C(n_156),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_225),
.C(n_226),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_40),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_227),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_40),
.C(n_37),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_37),
.C(n_147),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_37),
.C(n_147),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_105),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_233),
.CI(n_196),
.CON(n_238),
.SN(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_59),
.C(n_117),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_206),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_18),
.B1(n_17),
.B2(n_44),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_200),
.B1(n_202),
.B2(n_191),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_207),
.B1(n_217),
.B2(n_205),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_26),
.Y(n_233)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_255),
.B1(n_256),
.B2(n_2),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_240),
.Y(n_267)
);

NAND4xp25_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_199),
.C(n_211),
.D(n_195),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_192),
.B1(n_198),
.B2(n_17),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_249),
.B1(n_210),
.B2(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_246),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_227),
.A2(n_17),
.B1(n_26),
.B2(n_18),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_226),
.B1(n_225),
.B2(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_252),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_212),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_R g253 ( 
.A1(n_217),
.A2(n_26),
.B(n_27),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_214),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_26),
.B(n_1),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_0),
.B(n_2),
.Y(n_268)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_220),
.C(n_223),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_260),
.C(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_248),
.C(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_215),
.B1(n_17),
.B2(n_26),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_262),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_26),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_0),
.C(n_2),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_240),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_0),
.B(n_2),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_271),
.B(n_274),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_243),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_4),
.C(n_5),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.C(n_234),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_4),
.C(n_5),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_273),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_234),
.B1(n_238),
.B2(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_282),
.B(n_7),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_291),
.C(n_268),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_271),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_267),
.B(n_265),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_238),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_SL g297 ( 
.A1(n_289),
.A2(n_259),
.B(n_266),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_261),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_246),
.C(n_8),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_298),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_297),
.B(n_306),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_262),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_289),
.B1(n_282),
.B2(n_292),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_269),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_280),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_315),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_279),
.B(n_289),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_309),
.C(n_314),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_277),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_316),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_291),
.B(n_277),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_293),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_7),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_11),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_13),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_322),
.B(n_323),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_324),
.C(n_326),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_304),
.B(n_12),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_12),
.C(n_14),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_307),
.B(n_10),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_15),
.B(n_8),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_13),
.C(n_14),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_327),
.A2(n_15),
.B(n_8),
.C(n_9),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_15),
.C(n_8),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_331),
.B(n_332),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_7),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_330),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_335),
.B(n_9),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.Y(n_339)
);


endmodule