module fake_netlist_5_1471_n_1527 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_403, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_409, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_411, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1527);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_403;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1527;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

BUFx3_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

BUFx10_ASAP7_75t_L g415 ( 
.A(n_255),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_82),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_270),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_249),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_268),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_271),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_84),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_119),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_30),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_160),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_130),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_344),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_201),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_191),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_239),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_225),
.Y(n_433)
);

BUFx8_ASAP7_75t_SL g434 ( 
.A(n_79),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_281),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_244),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_145),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_71),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_220),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_228),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_150),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_284),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_93),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_262),
.B(n_299),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_15),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_29),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_305),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_44),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_153),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_331),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_303),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_113),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_102),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_186),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_411),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_44),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_219),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_89),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_137),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_177),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_157),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_223),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_66),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_0),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_178),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_43),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_26),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_320),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_162),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_277),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_333),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_51),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_232),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_348),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_5),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_396),
.Y(n_478)
);

BUFx8_ASAP7_75t_SL g479 ( 
.A(n_31),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_237),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_315),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_92),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_183),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_4),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_407),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_374),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_358),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_7),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_240),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_82),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_242),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_9),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_336),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_318),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_84),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_104),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_256),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_115),
.Y(n_499)
);

BUFx10_ASAP7_75t_L g500 ( 
.A(n_38),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_234),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_12),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_72),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_19),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_27),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_111),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_125),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_340),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_321),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_18),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_400),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_347),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_149),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_304),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_182),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_48),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_250),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_248),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_138),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_283),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_383),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_253),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_342),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_93),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_139),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_5),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_46),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_52),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_307),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_62),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_203),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_363),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_156),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_38),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_88),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_98),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_152),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_127),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_230),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_29),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_94),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_213),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_193),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_369),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_98),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_69),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_212),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_236),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_365),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_259),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_110),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_26),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_293),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_184),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_395),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_126),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_155),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_187),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_317),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_325),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_224),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_18),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_200),
.B(n_141),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_180),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_408),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_329),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_261),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_294),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_377),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_196),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_159),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_332),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_3),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_207),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_290),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_389),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_121),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_188),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_47),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_274),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_50),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_273),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_108),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_25),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_129),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_103),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_349),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_231),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_370),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_106),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_402),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_210),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_433),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_433),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_500),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_415),
.Y(n_598)
);

OA21x2_ASAP7_75t_L g599 ( 
.A1(n_524),
.A2(n_555),
.B(n_550),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_415),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_581),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_488),
.B(n_0),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_433),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_413),
.B(n_1),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_525),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_434),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_417),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_430),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_609)
);

BUFx8_ASAP7_75t_L g610 ( 
.A(n_501),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_413),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_581),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_424),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_529),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_581),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_424),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_587),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_430),
.A2(n_492),
.B1(n_416),
.B2(n_425),
.Y(n_618)
);

AND2x6_ASAP7_75t_L g619 ( 
.A(n_550),
.B(n_105),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_529),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_587),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_555),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_438),
.Y(n_623)
);

OA21x2_ASAP7_75t_L g624 ( 
.A1(n_585),
.A2(n_2),
.B(n_4),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_582),
.B(n_6),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_585),
.B(n_6),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_446),
.Y(n_627)
);

BUFx12f_ASAP7_75t_L g628 ( 
.A(n_417),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_457),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_459),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_504),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_414),
.Y(n_632)
);

AOI22x1_ASAP7_75t_SL g633 ( 
.A1(n_466),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_633)
);

BUFx12f_ASAP7_75t_L g634 ( 
.A(n_421),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_420),
.B(n_10),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_422),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_426),
.B(n_10),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_465),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_428),
.B(n_11),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_432),
.B(n_11),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_468),
.Y(n_641)
);

BUFx12f_ASAP7_75t_L g642 ( 
.A(n_421),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_444),
.Y(n_643)
);

NOR2x1_ASAP7_75t_L g644 ( 
.A(n_565),
.B(n_107),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_502),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_423),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_497),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_479),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_497),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_451),
.B(n_453),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_504),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_455),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_586),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_461),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_440),
.B(n_16),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_462),
.B(n_17),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_491),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_471),
.B(n_20),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_472),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_498),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_475),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_445),
.B(n_109),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_476),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_485),
.B(n_20),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_443),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_494),
.B(n_495),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_512),
.B(n_21),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_498),
.B(n_21),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_447),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_516),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_523),
.B(n_22),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_572),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_674),
.B(n_530),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_625),
.B(n_449),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_R g678 ( 
.A(n_667),
.B(n_469),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_602),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_598),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_R g681 ( 
.A(n_606),
.B(n_431),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_612),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_628),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_610),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_634),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_642),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_610),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_612),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_649),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_607),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_597),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_601),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_608),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_R g694 ( 
.A(n_662),
.B(n_478),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_609),
.A2(n_564),
.B1(n_482),
.B2(n_484),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_648),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_662),
.B(n_480),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_622),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_650),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_674),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

CKINVDCx16_ASAP7_75t_R g703 ( 
.A(n_618),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_605),
.B(n_429),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_674),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_671),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_622),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_613),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_613),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_644),
.B(n_594),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_595),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_616),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_596),
.B(n_531),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_626),
.B(n_593),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_595),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_616),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_616),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_617),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_617),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_670),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_611),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_617),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_621),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_R g724 ( 
.A(n_603),
.B(n_511),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_621),
.Y(n_725)
);

OA21x2_ASAP7_75t_L g726 ( 
.A1(n_668),
.A2(n_539),
.B(n_534),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_611),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_695),
.B(n_656),
.C(n_640),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_704),
.B(n_596),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_727),
.B(n_605),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_678),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_703),
.B(n_651),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_704),
.B(n_596),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_708),
.B(n_651),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_715),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_714),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_714),
.B(n_614),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_714),
.B(n_614),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_694),
.B(n_626),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_714),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_697),
.B(n_572),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_717),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_709),
.B(n_577),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_712),
.B(n_614),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_711),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_680),
.B(n_620),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_719),
.B(n_620),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_699),
.B(n_620),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_722),
.B(n_639),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_707),
.B(n_635),
.Y(n_750)
);

BUFx6f_ASAP7_75t_SL g751 ( 
.A(n_690),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_723),
.B(n_657),
.Y(n_752)
);

BUFx6f_ASAP7_75t_SL g753 ( 
.A(n_690),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_681),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_692),
.B(n_666),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_716),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_693),
.B(n_669),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_L g758 ( 
.A(n_710),
.B(n_619),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_682),
.B(n_635),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_718),
.Y(n_760)
);

BUFx8_ASAP7_75t_L g761 ( 
.A(n_725),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_701),
.B(n_418),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_688),
.B(n_726),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_677),
.B(n_647),
.C(n_558),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_711),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_702),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_726),
.B(n_637),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_706),
.B(n_514),
.C(n_517),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_710),
.B(n_637),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_696),
.B(n_700),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_675),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_L g772 ( 
.A(n_679),
.B(n_599),
.C(n_624),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_676),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_710),
.B(n_660),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_713),
.Y(n_775)
);

NOR3xp33_ASAP7_75t_L g776 ( 
.A(n_691),
.B(n_542),
.C(n_538),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_721),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_705),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_724),
.B(n_720),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_683),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_685),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_686),
.B(n_673),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_689),
.B(n_673),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_684),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_687),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_SL g786 ( 
.A(n_695),
.B(n_520),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_695),
.B(n_554),
.C(n_543),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_711),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_698),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_727),
.B(n_632),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_717),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_704),
.B(n_595),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_717),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_695),
.B(n_583),
.C(n_575),
.Y(n_794)
);

NOR3xp33_ASAP7_75t_L g795 ( 
.A(n_695),
.B(n_489),
.C(n_474),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_704),
.B(n_604),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_708),
.B(n_631),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_727),
.B(n_588),
.Y(n_798)
);

AND2x6_ASAP7_75t_SL g799 ( 
.A(n_783),
.B(n_623),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_792),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_749),
.B(n_599),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_754),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_627),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_791),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_796),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_728),
.A2(n_767),
.B1(n_763),
.B2(n_787),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_752),
.B(n_619),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_755),
.B(n_619),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_771),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_797),
.B(n_731),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_770),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_757),
.B(n_535),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_769),
.A2(n_556),
.B1(n_562),
.B2(n_544),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_732),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_794),
.A2(n_764),
.B1(n_795),
.B2(n_664),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_773),
.B(n_790),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_739),
.B(n_573),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_786),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_786),
.B(n_493),
.Y(n_819)
);

INVx8_ASAP7_75t_L g820 ( 
.A(n_785),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_793),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_750),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_785),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_735),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_774),
.B(n_540),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_734),
.B(n_419),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_780),
.B(n_630),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_788),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_772),
.A2(n_664),
.B1(n_624),
.B2(n_552),
.Y(n_829)
);

INVx5_ASAP7_75t_L g830 ( 
.A(n_736),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_745),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_729),
.B(n_545),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_765),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_772),
.A2(n_664),
.B1(n_560),
.B2(n_563),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_733),
.B(n_553),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_741),
.B(n_658),
.C(n_646),
.Y(n_837)
);

AND2x2_ASAP7_75t_SL g838 ( 
.A(n_768),
.B(n_776),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_SL g839 ( 
.A(n_779),
.B(n_505),
.C(n_503),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_777),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_730),
.B(n_427),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_759),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_756),
.Y(n_843)
);

AOI22x1_ASAP7_75t_L g844 ( 
.A1(n_789),
.A2(n_645),
.B1(n_571),
.B2(n_574),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_760),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_748),
.Y(n_846)
);

BUFx4f_ASAP7_75t_L g847 ( 
.A(n_778),
.Y(n_847)
);

BUFx5_ASAP7_75t_L g848 ( 
.A(n_775),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_737),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_738),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_743),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_744),
.B(n_568),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_781),
.B(n_629),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_747),
.B(n_580),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_761),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_782),
.B(n_746),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_761),
.Y(n_857)
);

OR2x2_ASAP7_75t_SL g858 ( 
.A(n_798),
.B(n_633),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_762),
.A2(n_590),
.B1(n_592),
.B2(n_584),
.Y(n_859)
);

AND2x6_ASAP7_75t_SL g860 ( 
.A(n_784),
.B(n_659),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_751),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_758),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_740),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_751),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_753),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_753),
.Y(n_866)
);

INVx5_ASAP7_75t_L g867 ( 
.A(n_788),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_792),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_749),
.B(n_664),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_791),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_791),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_792),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_742),
.B(n_638),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_731),
.B(n_435),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_728),
.A2(n_636),
.B1(n_643),
.B2(n_632),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_792),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_754),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_749),
.B(n_636),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_731),
.B(n_510),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_767),
.A2(n_641),
.B(n_437),
.C(n_439),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_792),
.Y(n_881)
);

OR2x4_ASAP7_75t_L g882 ( 
.A(n_732),
.B(n_652),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_788),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_749),
.B(n_636),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_792),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_728),
.A2(n_441),
.B1(n_442),
.B2(n_436),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_728),
.A2(n_653),
.B1(n_655),
.B2(n_643),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_731),
.B(n_448),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_731),
.B(n_450),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_SL g890 ( 
.A1(n_786),
.A2(n_633),
.B1(n_589),
.B2(n_588),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_SL g891 ( 
.A(n_786),
.B(n_528),
.C(n_527),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_749),
.B(n_643),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_783),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_792),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_749),
.B(n_653),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_749),
.B(n_653),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_749),
.B(n_655),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_766),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_749),
.B(n_655),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_728),
.A2(n_454),
.B1(n_456),
.B2(n_452),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_731),
.B(n_458),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_792),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_731),
.B(n_532),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_791),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_822),
.B(n_460),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_811),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_812),
.B(n_536),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_836),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_806),
.A2(n_464),
.B1(n_467),
.B2(n_463),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_800),
.B(n_805),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_818),
.A2(n_473),
.B1(n_481),
.B2(n_470),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_868),
.B(n_483),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_813),
.B(n_537),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_810),
.B(n_879),
.Y(n_914)
);

OAI21xp33_ASAP7_75t_L g915 ( 
.A1(n_819),
.A2(n_548),
.B(n_547),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_821),
.B(n_870),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_904),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_903),
.A2(n_487),
.B(n_490),
.C(n_486),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_872),
.B(n_499),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_820),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_804),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_801),
.A2(n_507),
.B(n_506),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_876),
.B(n_508),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_SL g924 ( 
.A(n_839),
.B(n_509),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_836),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_881),
.B(n_513),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_893),
.B(n_515),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_898),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_862),
.A2(n_519),
.B1(n_521),
.B2(n_518),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_L g930 ( 
.A(n_836),
.B(n_522),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_885),
.B(n_526),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_804),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_891),
.A2(n_661),
.B1(n_665),
.B2(n_663),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_804),
.B(n_631),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_863),
.A2(n_807),
.B(n_829),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_842),
.B(n_654),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_845),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_847),
.B(n_803),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_825),
.A2(n_541),
.B(n_546),
.C(n_533),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_817),
.B(n_549),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_894),
.B(n_902),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_849),
.A2(n_557),
.B(n_551),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_L g943 ( 
.A(n_802),
.B(n_877),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_815),
.A2(n_561),
.B1(n_566),
.B2(n_559),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_874),
.B(n_567),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_808),
.A2(n_570),
.B(n_569),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_850),
.A2(n_578),
.B(n_576),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_878),
.B(n_579),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_884),
.B(n_892),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_871),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_823),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_824),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_820),
.B(n_661),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_895),
.B(n_591),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_856),
.B(n_672),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_896),
.B(n_22),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_897),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_882),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_888),
.A2(n_27),
.B(n_23),
.C(n_24),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_830),
.B(n_112),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_873),
.B(n_28),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_SL g962 ( 
.A(n_841),
.B(n_28),
.C(n_31),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_889),
.B(n_32),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_901),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_853),
.Y(n_965)
);

OAI22x1_ASAP7_75t_L g966 ( 
.A1(n_844),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_L g967 ( 
.A(n_830),
.B(n_114),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_814),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_899),
.B(n_35),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_851),
.B(n_116),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_890),
.B(n_36),
.C(n_37),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_R g972 ( 
.A(n_864),
.B(n_117),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_840),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_833),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_834),
.A2(n_120),
.B1(n_122),
.B2(n_118),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_848),
.B(n_846),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_SL g977 ( 
.A(n_826),
.B(n_866),
.C(n_865),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_848),
.B(n_37),
.Y(n_978)
);

BUFx12f_ASAP7_75t_L g979 ( 
.A(n_860),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_886),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_SL g981 ( 
.A1(n_838),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_832),
.A2(n_124),
.B(n_123),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_900),
.A2(n_45),
.B(n_42),
.C(n_43),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_835),
.A2(n_46),
.B(n_42),
.C(n_45),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_843),
.B(n_47),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_855),
.B(n_857),
.Y(n_986)
);

INVx3_ASAP7_75t_SL g987 ( 
.A(n_871),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_SL g988 ( 
.A1(n_875),
.A2(n_48),
.B(n_49),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_848),
.B(n_128),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_887),
.A2(n_132),
.B1(n_133),
.B2(n_131),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_852),
.A2(n_135),
.B1(n_136),
.B2(n_134),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_848),
.B(n_49),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_SL g993 ( 
.A(n_837),
.B(n_50),
.C(n_51),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_854),
.B(n_52),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_853),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_799),
.Y(n_996)
);

NOR2xp67_ASAP7_75t_L g997 ( 
.A(n_861),
.B(n_140),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_831),
.B(n_53),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_859),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_828),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_828),
.B(n_142),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_867),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_827),
.A2(n_883),
.B(n_144),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_883),
.A2(n_146),
.B1(n_147),
.B2(n_143),
.Y(n_1004)
);

CKINVDCx6p67_ASAP7_75t_R g1005 ( 
.A(n_883),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_858),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_893),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_822),
.B(n_56),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_SL g1009 ( 
.A1(n_880),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1009)
);

AO22x1_ASAP7_75t_L g1010 ( 
.A1(n_819),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_821),
.B(n_148),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_809),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_819),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_809),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_SL g1015 ( 
.A1(n_806),
.A2(n_154),
.B(n_158),
.C(n_151),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_819),
.A2(n_64),
.B1(n_61),
.B2(n_63),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_818),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_818),
.A2(n_163),
.B1(n_164),
.B2(n_161),
.Y(n_1018)
);

O2A1O1Ixp5_ASAP7_75t_L g1019 ( 
.A1(n_808),
.A2(n_166),
.B(n_167),
.C(n_165),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_809),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_836),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_804),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_SL g1023 ( 
.A1(n_880),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_819),
.A2(n_67),
.B(n_68),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_822),
.B(n_68),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_814),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_818),
.A2(n_169),
.B1(n_170),
.B2(n_168),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_819),
.B(n_70),
.C(n_71),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_816),
.B(n_171),
.Y(n_1029)
);

AND2x4_ASAP7_75t_SL g1030 ( 
.A(n_823),
.B(n_172),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_821),
.B(n_173),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_836),
.B(n_174),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_804),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_819),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_869),
.A2(n_176),
.B(n_175),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_819),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_836),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_818),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_811),
.B(n_78),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_822),
.B(n_78),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_SL g1041 ( 
.A1(n_880),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_819),
.A2(n_83),
.B(n_80),
.C(n_81),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_821),
.B(n_179),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_893),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_810),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_SL g1046 ( 
.A(n_839),
.B(n_85),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_819),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_811),
.B(n_86),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_935),
.A2(n_185),
.B(n_181),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_906),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_949),
.A2(n_969),
.B(n_956),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_928),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_910),
.B(n_87),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_908),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_976),
.A2(n_190),
.B(n_189),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_986),
.B(n_88),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_1026),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1045),
.B(n_936),
.Y(n_1058)
);

OA21x2_ASAP7_75t_L g1059 ( 
.A1(n_978),
.A2(n_992),
.B(n_1019),
.Y(n_1059)
);

CKINVDCx11_ASAP7_75t_R g1060 ( 
.A(n_979),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_925),
.Y(n_1061)
);

BUFx8_ASAP7_75t_L g1062 ( 
.A(n_950),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_987),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_922),
.A2(n_194),
.B(n_192),
.Y(n_1064)
);

OR2x6_ASAP7_75t_L g1065 ( 
.A(n_986),
.B(n_89),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_989),
.A2(n_197),
.B(n_195),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_941),
.A2(n_199),
.B(n_198),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_1022),
.B(n_202),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_914),
.B(n_90),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_921),
.B(n_204),
.Y(n_1070)
);

BUFx2_ASAP7_75t_R g1071 ( 
.A(n_951),
.Y(n_1071)
);

AOI22x1_ASAP7_75t_L g1072 ( 
.A1(n_966),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_932),
.B(n_205),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1008),
.A2(n_208),
.B(n_206),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_937),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_952),
.Y(n_1076)
);

AO21x2_ASAP7_75t_L g1077 ( 
.A1(n_1029),
.A2(n_211),
.B(n_209),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_968),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1012),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_955),
.B(n_1025),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1014),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_925),
.Y(n_1082)
);

NAND2x1p5_ASAP7_75t_L g1083 ( 
.A(n_1033),
.B(n_214),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_SL g1084 ( 
.A(n_917),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_982),
.A2(n_216),
.B(n_215),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1003),
.A2(n_218),
.B(n_217),
.Y(n_1086)
);

AO21x2_ASAP7_75t_L g1087 ( 
.A1(n_1015),
.A2(n_222),
.B(n_221),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1020),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_943),
.B(n_91),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_958),
.Y(n_1090)
);

BUFx2_ASAP7_75t_R g1091 ( 
.A(n_938),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_925),
.Y(n_1092)
);

INVx5_ASAP7_75t_L g1093 ( 
.A(n_1021),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1021),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_950),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_916),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1007),
.B(n_94),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_916),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_920),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_960),
.A2(n_227),
.B(n_226),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1044),
.B(n_95),
.Y(n_1101)
);

AO21x2_ASAP7_75t_L g1102 ( 
.A1(n_948),
.A2(n_233),
.B(n_229),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_973),
.B(n_95),
.Y(n_1103)
);

AO21x2_ASAP7_75t_L g1104 ( 
.A1(n_954),
.A2(n_238),
.B(n_235),
.Y(n_1104)
);

AND2x6_ASAP7_75t_SL g1105 ( 
.A(n_1039),
.B(n_96),
.Y(n_1105)
);

INVx3_ASAP7_75t_SL g1106 ( 
.A(n_996),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_974),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1021),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_907),
.A2(n_96),
.B(n_97),
.C(n_99),
.Y(n_1109)
);

CKINVDCx11_ASAP7_75t_R g1110 ( 
.A(n_953),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_1037),
.B(n_241),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_913),
.B(n_97),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_953),
.B(n_99),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_1037),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1002),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1002),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_1002),
.Y(n_1117)
);

BUFx2_ASAP7_75t_SL g1118 ( 
.A(n_1011),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_961),
.Y(n_1119)
);

INVx6_ASAP7_75t_L g1120 ( 
.A(n_996),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_946),
.A2(n_918),
.B(n_1035),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_SL g1122 ( 
.A1(n_1048),
.A2(n_100),
.B1(n_101),
.B2(n_243),
.Y(n_1122)
);

INVx6_ASAP7_75t_SL g1123 ( 
.A(n_1011),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_1031),
.B(n_245),
.Y(n_1124)
);

INVx5_ASAP7_75t_L g1125 ( 
.A(n_1031),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1005),
.Y(n_1126)
);

BUFx2_ASAP7_75t_R g1127 ( 
.A(n_1000),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1040),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_965),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1043),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_934),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_994),
.A2(n_327),
.B(n_409),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_988),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_998),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1032),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1030),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_985),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_996),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_912),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_919),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_923),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_905),
.A2(n_326),
.B(n_404),
.Y(n_1142)
);

BUFx2_ASAP7_75t_SL g1143 ( 
.A(n_997),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_967),
.A2(n_324),
.B(n_401),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_927),
.B(n_100),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_963),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_926),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_945),
.A2(n_334),
.B(n_246),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1009),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_975),
.A2(n_335),
.B(n_247),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_931),
.B(n_995),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_970),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_924),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1023),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_939),
.A2(n_1004),
.B(n_991),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_977),
.B(n_251),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1041),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1028),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_940),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_957),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_972),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_990),
.A2(n_337),
.B(n_252),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1010),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_942),
.A2(n_338),
.B(n_254),
.Y(n_1164)
);

BUFx12f_ASAP7_75t_L g1165 ( 
.A(n_1046),
.Y(n_1165)
);

INVx5_ASAP7_75t_L g1166 ( 
.A(n_1001),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_947),
.A2(n_341),
.B(n_257),
.Y(n_1167)
);

INVx2_ASAP7_75t_R g1168 ( 
.A(n_1018),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1024),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_959),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_911),
.Y(n_1171)
);

BUFx2_ASAP7_75t_SL g1172 ( 
.A(n_1027),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_909),
.A2(n_1047),
.B(n_1042),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_929),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_971),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_930),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_993),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_964),
.A2(n_933),
.B(n_944),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_915),
.A2(n_343),
.B(n_258),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_962),
.B(n_981),
.Y(n_1180)
);

BUFx2_ASAP7_75t_SL g1181 ( 
.A(n_980),
.Y(n_1181)
);

AO21x2_ASAP7_75t_L g1182 ( 
.A1(n_1013),
.A2(n_1034),
.B(n_983),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1006),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_984),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1016),
.Y(n_1185)
);

BUFx2_ASAP7_75t_R g1186 ( 
.A(n_1017),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1036),
.A2(n_345),
.B(n_260),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_999),
.A2(n_346),
.B(n_263),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1187),
.A2(n_1145),
.B1(n_1181),
.B2(n_1185),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1078),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1177),
.A2(n_1181),
.B1(n_1180),
.B2(n_1168),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1088),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1058),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1146),
.B(n_1038),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1054),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1128),
.B(n_101),
.Y(n_1196)
);

BUFx12f_ASAP7_75t_L g1197 ( 
.A(n_1110),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1175),
.B(n_264),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1172),
.A2(n_1125),
.B1(n_1128),
.B2(n_1133),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1183),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1063),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1141),
.B(n_269),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1172),
.A2(n_272),
.B1(n_275),
.B2(n_276),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1117),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1090),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1139),
.B(n_278),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1117),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1075),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1079),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1081),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1057),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1054),
.Y(n_1213)
);

AOI222xp33_ASAP7_75t_L g1214 ( 
.A1(n_1177),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.C1(n_285),
.C2(n_286),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1119),
.B(n_287),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1177),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1076),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1052),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1107),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1125),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1169),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1140),
.B(n_297),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1053),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1069),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1099),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1049),
.A2(n_298),
.B(n_300),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1125),
.B(n_412),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1159),
.B(n_301),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1057),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1133),
.A2(n_302),
.B1(n_306),
.B2(n_308),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1062),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1093),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1137),
.B(n_399),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1062),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1149),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1064),
.A2(n_309),
.B(n_310),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1149),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1120),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1126),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_SL g1240 ( 
.A(n_1123),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1112),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_1241)
);

NOR2x1_ASAP7_75t_R g1242 ( 
.A(n_1050),
.B(n_314),
.Y(n_1242)
);

AO21x1_ASAP7_75t_L g1243 ( 
.A1(n_1154),
.A2(n_1157),
.B(n_1179),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_SL g1244 ( 
.A(n_1123),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1060),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1098),
.B(n_316),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1129),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1130),
.B(n_398),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1118),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1157),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1118),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1097),
.B(n_353),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1158),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1184),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1134),
.Y(n_1255)
);

BUFx2_ASAP7_75t_R g1256 ( 
.A(n_1106),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1116),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1160),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1115),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1070),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1120),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1073),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1115),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1163),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1132),
.A2(n_362),
.B(n_364),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1092),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1101),
.B(n_366),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1061),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1094),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1130),
.A2(n_367),
.B1(n_368),
.B2(n_371),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1130),
.A2(n_372),
.B1(n_373),
.B2(n_376),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1108),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1080),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1096),
.B(n_1147),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1126),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1174),
.A2(n_1173),
.B1(n_1182),
.B2(n_1122),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1071),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1170),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1093),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1072),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1136),
.Y(n_1281)
);

OAI22x1_ASAP7_75t_L g1282 ( 
.A1(n_1072),
.A2(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1152),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1171),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1091),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1095),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1153),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1165),
.A2(n_388),
.B1(n_390),
.B2(n_391),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1151),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1114),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1105),
.Y(n_1291)
);

BUFx2_ASAP7_75t_R g1292 ( 
.A(n_1138),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1061),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1051),
.B(n_397),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1082),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1190),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1195),
.Y(n_1297)
);

NOR3xp33_ASAP7_75t_SL g1298 ( 
.A(n_1277),
.B(n_1109),
.C(n_1103),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1195),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1193),
.B(n_1161),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1225),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1205),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1193),
.B(n_1161),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1189),
.A2(n_1156),
.B1(n_1074),
.B2(n_1142),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1274),
.B(n_1161),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1235),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1273),
.B(n_1166),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1201),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1289),
.B(n_1135),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1229),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1236),
.A2(n_1089),
.B1(n_1067),
.B2(n_1113),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1237),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1247),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1194),
.B(n_1089),
.Y(n_1314)
);

NOR3xp33_ASAP7_75t_SL g1315 ( 
.A(n_1228),
.B(n_1055),
.C(n_1100),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1260),
.B(n_1131),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1289),
.B(n_1198),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1212),
.Y(n_1318)
);

CKINVDCx6p67_ASAP7_75t_R g1319 ( 
.A(n_1197),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1295),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1195),
.Y(n_1321)
);

CKINVDCx16_ASAP7_75t_R g1322 ( 
.A(n_1245),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1239),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1287),
.Y(n_1324)
);

INVx4_ASAP7_75t_L g1325 ( 
.A(n_1213),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1236),
.A2(n_1214),
.B1(n_1191),
.B2(n_1223),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1234),
.B(n_1056),
.Y(n_1327)
);

NAND3xp33_ASAP7_75t_SL g1328 ( 
.A(n_1214),
.B(n_1124),
.C(n_1186),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1224),
.B(n_1166),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1192),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1252),
.B(n_1065),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1233),
.A2(n_1176),
.B1(n_1084),
.B2(n_1143),
.Y(n_1332)
);

OR2x2_ASAP7_75t_SL g1333 ( 
.A(n_1239),
.B(n_1196),
.Y(n_1333)
);

NOR3xp33_ASAP7_75t_SL g1334 ( 
.A(n_1241),
.B(n_1127),
.C(n_1113),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1243),
.A2(n_1176),
.B1(n_1143),
.B2(n_1135),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1275),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_R g1337 ( 
.A(n_1227),
.B(n_1065),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1256),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1255),
.B(n_1166),
.Y(n_1339)
);

NOR3xp33_ASAP7_75t_SL g1340 ( 
.A(n_1202),
.B(n_1056),
.C(n_1135),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1267),
.B(n_1215),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_SL g1342 ( 
.A(n_1238),
.B(n_1261),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1292),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1211),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1213),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1294),
.A2(n_1178),
.B(n_1155),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1209),
.B(n_1210),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1268),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1221),
.B(n_1111),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1199),
.A2(n_1068),
.B1(n_1083),
.B2(n_1059),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1262),
.B(n_1148),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1250),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1240),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1285),
.A2(n_1246),
.B1(n_1276),
.B2(n_1206),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1232),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1244),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1203),
.A2(n_1144),
.B1(n_1162),
.B2(n_1150),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1281),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1285),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1265),
.A2(n_1087),
.A3(n_1121),
.B(n_1188),
.Y(n_1360)
);

CKINVDCx16_ASAP7_75t_R g1361 ( 
.A(n_1231),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1254),
.B(n_1077),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1290),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_SL g1364 ( 
.A(n_1222),
.B(n_1104),
.C(n_1102),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1217),
.B(n_1066),
.Y(n_1365)
);

XOR2x2_ASAP7_75t_SL g1366 ( 
.A(n_1291),
.B(n_392),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1286),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_R g1368 ( 
.A(n_1204),
.B(n_394),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1203),
.A2(n_1167),
.B1(n_1086),
.B2(n_1164),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1293),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1219),
.B(n_1085),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1258),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_R g1373 ( 
.A(n_1207),
.B(n_1259),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1279),
.Y(n_1374)
);

AND2x2_ASAP7_75t_SL g1375 ( 
.A(n_1226),
.B(n_1216),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1280),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1283),
.B(n_1208),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1263),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1359),
.B(n_1242),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1306),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1328),
.A2(n_1264),
.B1(n_1278),
.B2(n_1230),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1312),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1372),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1312),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1352),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1352),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1296),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1318),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1351),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1330),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1371),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1323),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1376),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1333),
.B(n_1218),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1363),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1377),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1347),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1317),
.B(n_1282),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1341),
.B(n_1266),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1308),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1362),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1302),
.B(n_1248),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1320),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1365),
.B(n_1272),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1346),
.B(n_1257),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1370),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1349),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1313),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_1309),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1326),
.B(n_1269),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1307),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1360),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1348),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1373),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1311),
.A2(n_1253),
.B1(n_1200),
.B2(n_1284),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1360),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1314),
.B(n_1305),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1339),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1354),
.B(n_1251),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1389),
.B(n_1375),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1389),
.B(n_1360),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1388),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1391),
.B(n_1335),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1380),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1383),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1380),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1409),
.B(n_1300),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1391),
.B(n_1303),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1384),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1391),
.B(n_1401),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1397),
.B(n_1329),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1401),
.B(n_1304),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1392),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1385),
.B(n_1364),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1415),
.B(n_1298),
.C(n_1315),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1395),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1395),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1400),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1407),
.B(n_1332),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1411),
.B(n_1331),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1382),
.B(n_1357),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1396),
.B(n_1340),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1381),
.A2(n_1334),
.B1(n_1327),
.B2(n_1200),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1403),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1390),
.B(n_1350),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1400),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1405),
.B(n_1369),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1424),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1440),
.B(n_1379),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1437),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1426),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1438),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1430),
.B(n_1416),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1421),
.B(n_1412),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1434),
.B(n_1393),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1420),
.B(n_1417),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1429),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1425),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1420),
.B(n_1417),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_SL g1461 ( 
.A(n_1435),
.B(n_1393),
.Y(n_1461)
);

AND2x4_ASAP7_75t_SL g1462 ( 
.A(n_1428),
.B(n_1404),
.Y(n_1462)
);

NOR3xp33_ASAP7_75t_L g1463 ( 
.A(n_1436),
.B(n_1419),
.C(n_1418),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1435),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1448),
.B(n_1405),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1422),
.B(n_1406),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1443),
.B(n_1408),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1421),
.B(n_1398),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1447),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1450),
.A2(n_1444),
.B1(n_1419),
.B2(n_1439),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1458),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1463),
.A2(n_1432),
.B1(n_1337),
.B2(n_1442),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1458),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1449),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1469),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1456),
.B(n_1428),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1465),
.B(n_1445),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1467),
.B(n_1433),
.Y(n_1478)
);

O2A1O1Ixp33_ASAP7_75t_SL g1479 ( 
.A1(n_1466),
.A2(n_1414),
.B(n_1441),
.C(n_1431),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1465),
.B(n_1432),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1452),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1464),
.A2(n_1249),
.B1(n_1251),
.B2(n_1410),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1459),
.Y(n_1483)
);

OAI32xp33_ASAP7_75t_L g1484 ( 
.A1(n_1455),
.A2(n_1454),
.A3(n_1394),
.B1(n_1451),
.B2(n_1427),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1457),
.B(n_1446),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1483),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_SL g1487 ( 
.A(n_1472),
.B(n_1453),
.C(n_1394),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1470),
.B(n_1446),
.C(n_1453),
.Y(n_1488)
);

NOR3xp33_ASAP7_75t_L g1489 ( 
.A(n_1479),
.B(n_1402),
.C(n_1322),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1482),
.A2(n_1428),
.B1(n_1398),
.B2(n_1423),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1476),
.Y(n_1491)
);

OAI21xp33_ASAP7_75t_L g1492 ( 
.A1(n_1482),
.A2(n_1460),
.B(n_1457),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1480),
.A2(n_1469),
.B1(n_1462),
.B2(n_1468),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1489),
.A2(n_1477),
.B1(n_1478),
.B2(n_1475),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1486),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1492),
.B(n_1319),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1491),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1487),
.A2(n_1288),
.B(n_1414),
.Y(n_1498)
);

NOR3xp33_ASAP7_75t_L g1499 ( 
.A(n_1496),
.B(n_1488),
.C(n_1361),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1494),
.A2(n_1490),
.B(n_1484),
.C(n_1493),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1498),
.A2(n_1461),
.B(n_1301),
.Y(n_1501)
);

NOR2xp67_ASAP7_75t_L g1502 ( 
.A(n_1497),
.B(n_1476),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1495),
.A2(n_1481),
.B(n_1474),
.Y(n_1503)
);

XNOR2xp5_ASAP7_75t_L g1504 ( 
.A(n_1494),
.B(n_1310),
.Y(n_1504)
);

OA22x2_ASAP7_75t_L g1505 ( 
.A1(n_1504),
.A2(n_1327),
.B1(n_1462),
.B2(n_1387),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1500),
.B(n_1485),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1501),
.A2(n_1342),
.B(n_1242),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1506),
.A2(n_1502),
.B1(n_1499),
.B2(n_1503),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_SL g1509 ( 
.A1(n_1507),
.A2(n_1356),
.B(n_1324),
.C(n_1358),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1508),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1510),
.A2(n_1509),
.B1(n_1505),
.B2(n_1336),
.C(n_1338),
.Y(n_1511)
);

AOI32xp33_ASAP7_75t_L g1512 ( 
.A1(n_1511),
.A2(n_1408),
.A3(n_1353),
.B1(n_1343),
.B2(n_1392),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1511),
.Y(n_1513)
);

INVx3_ASAP7_75t_SL g1514 ( 
.A(n_1513),
.Y(n_1514)
);

NOR3xp33_ASAP7_75t_L g1515 ( 
.A(n_1512),
.B(n_1367),
.C(n_1344),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1515),
.A2(n_1413),
.B1(n_1378),
.B2(n_1399),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1514),
.B(n_1471),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1516),
.A2(n_1413),
.B1(n_1399),
.B2(n_1297),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1517),
.Y(n_1519)
);

OAI22x1_ASAP7_75t_L g1520 ( 
.A1(n_1519),
.A2(n_1366),
.B1(n_1325),
.B2(n_1374),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1518),
.A2(n_1473),
.B1(n_1297),
.B2(n_1299),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1520),
.A2(n_1249),
.B(n_1270),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1521),
.B(n_1316),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1523),
.A2(n_1297),
.B1(n_1321),
.B2(n_1325),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1522),
.A2(n_1345),
.B1(n_1355),
.B2(n_1374),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1524),
.A2(n_1220),
.B1(n_1271),
.B2(n_1270),
.C(n_1368),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1526),
.A2(n_1525),
.B1(n_1345),
.B2(n_1355),
.Y(n_1527)
);


endmodule