module fake_netlist_1_8362_n_1724 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_381, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1724);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_381;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1724;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_1671;
wire n_646;
wire n_1334;
wire n_1627;
wire n_1698;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_1646;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_1667;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_1663;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_1714;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1672;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_1661;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1683;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_1656;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_1654;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1718;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1620;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_1707;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_1693;
wire n_1690;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1703;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1711;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_1716;
wire n_1662;
wire n_790;
wire n_761;
wire n_1660;
wire n_1287;
wire n_472;
wire n_1100;
wire n_1648;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_1695;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1682;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_1694;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_753;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1681;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_1675;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1709;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1670;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1643;
wire n_1687;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_1710;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1647;
wire n_1621;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1668;
wire n_1692;
wire n_1153;
wire n_1657;
wire n_1655;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_1665;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1696;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1645;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1626;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1577;
wire n_1719;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_1705;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1697;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_1720;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1679;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_1688;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1653;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1658;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1659;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1701;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1704;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1609;
wire n_1576;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1684;
wire n_1089;
wire n_1717;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1706;
wire n_1473;
wire n_1678;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1674;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1712;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_1700;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1722;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_584;
wire n_1130;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1689;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_1699;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_1713;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_1676;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_1708;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1204;
wire n_1094;
wire n_1666;
wire n_392;
wire n_1169;
wire n_975;
wire n_1721;
wire n_1081;
wire n_1680;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_1669;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1673;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_1664;
wire n_682;
wire n_1607;
wire n_906;
wire n_1650;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1702;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1685;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1677;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1649;
wire n_1143;
wire n_629;
wire n_1723;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_1691;
wire n_1715;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_1686;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1651;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_1652;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g383 ( .A(n_309), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_41), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_265), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_305), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_178), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_365), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_7), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_261), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_213), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_159), .Y(n_392) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_41), .B(n_314), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_146), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_343), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_167), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_81), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_315), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_43), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_97), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_258), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_229), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_102), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_316), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_12), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_235), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_101), .B(n_230), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_295), .Y(n_409) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_162), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_350), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_21), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_220), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_2), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_224), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_311), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_202), .Y(n_417) );
CKINVDCx14_ASAP7_75t_R g418 ( .A(n_344), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_160), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_32), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_267), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_274), .B(n_328), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_143), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_114), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_308), .Y(n_425) );
INVxp33_ASAP7_75t_SL g426 ( .A(n_158), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_243), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_183), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_368), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_133), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_155), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_307), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_374), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_359), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_372), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_2), .Y(n_436) );
BUFx2_ASAP7_75t_SL g437 ( .A(n_166), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_44), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_245), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_114), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_289), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_35), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_67), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_214), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_152), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_250), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_278), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_340), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_244), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_341), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_312), .B(n_140), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g452 ( .A(n_130), .B(n_110), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_163), .B(n_58), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_53), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_347), .Y(n_455) );
INVxp33_ASAP7_75t_SL g456 ( .A(n_285), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_141), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_182), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_326), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_241), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_331), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_248), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_358), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_266), .Y(n_464) );
INVxp33_ASAP7_75t_SL g465 ( .A(n_24), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_171), .Y(n_466) );
INVxp33_ASAP7_75t_SL g467 ( .A(n_318), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_67), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_209), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_349), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_193), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_128), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_256), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_102), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_299), .Y(n_475) );
INVxp33_ASAP7_75t_SL g476 ( .A(n_303), .Y(n_476) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_112), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_354), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_16), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_255), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_217), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_123), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_119), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_100), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_98), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_324), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_63), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_154), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_283), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_281), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_84), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_323), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_177), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_17), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_16), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_168), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_313), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_237), .Y(n_498) );
BUFx8_ASAP7_75t_SL g499 ( .A(n_101), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_173), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_290), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_271), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_26), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_132), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_9), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_197), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_139), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_76), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_126), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_221), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_57), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_275), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_29), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_227), .Y(n_514) );
BUFx3_ASAP7_75t_L g515 ( .A(n_280), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_117), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_175), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_153), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_79), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_273), .Y(n_520) );
CKINVDCx14_ASAP7_75t_R g521 ( .A(n_23), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_77), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_367), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_56), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_124), .Y(n_525) );
BUFx8_ASAP7_75t_SL g526 ( .A(n_251), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_376), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_46), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_30), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_26), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_306), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_96), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_262), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_34), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_284), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_40), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_72), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_296), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_18), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_94), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_233), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_38), .Y(n_542) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_66), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_74), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_236), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_117), .B(n_20), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_77), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_83), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_106), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_302), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_17), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_14), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_179), .Y(n_553) );
CKINVDCx14_ASAP7_75t_R g554 ( .A(n_27), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_379), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_49), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_165), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_211), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_357), .Y(n_559) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_34), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_188), .B(n_147), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_109), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_161), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_184), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_198), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_362), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_27), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_361), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_144), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_320), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_135), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_112), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_0), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_304), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_330), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_346), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_404), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_388), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_404), .Y(n_579) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_388), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_521), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_436), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_516), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_433), .B(n_0), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_526), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_521), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_436), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_388), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_443), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_443), .B(n_1), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_388), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_420), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_420), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_498), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_498), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_526), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_395), .B(n_1), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_498), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_536), .Y(n_599) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_498), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_416), .Y(n_601) );
AND2x6_ASAP7_75t_L g602 ( .A(n_478), .B(n_121), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_554), .Y(n_603) );
AND2x6_ASAP7_75t_L g604 ( .A(n_478), .B(n_122), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_446), .B(n_3), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_421), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_495), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_536), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_495), .B(n_3), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_556), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_458), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_556), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_515), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_397), .B(n_4), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_464), .B(n_497), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_573), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_554), .B(n_4), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_505), .Y(n_619) );
AND2x6_ASAP7_75t_L g620 ( .A(n_609), .B(n_515), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_601), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_581), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_586), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_601), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_609), .A2(n_401), .B1(n_406), .B2(n_399), .Y(n_625) );
INVx5_ASAP7_75t_L g626 ( .A(n_602), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_601), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_587), .B(n_416), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_607), .Y(n_629) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_578), .Y(n_630) );
INVx5_ASAP7_75t_L g631 ( .A(n_602), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_609), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_586), .B(n_418), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_587), .B(n_505), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_603), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_587), .B(n_461), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_603), .B(n_500), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_585), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_587), .B(n_418), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_589), .B(n_461), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_607), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_589), .B(n_414), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_615), .B(n_386), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_617), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_583), .B(n_387), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_589), .B(n_386), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_609), .Y(n_647) );
NOR2xp33_ASAP7_75t_SL g648 ( .A(n_602), .B(n_394), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_589), .B(n_396), .Y(n_649) );
INVx4_ASAP7_75t_L g650 ( .A(n_602), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_578), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_578), .Y(n_652) );
OAI22xp5_ASAP7_75t_SL g653 ( .A1(n_596), .A2(n_384), .B1(n_487), .B2(n_442), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_617), .Y(n_654) );
AO21x2_ASAP7_75t_L g655 ( .A1(n_614), .A2(n_422), .B(n_385), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_577), .B(n_402), .Y(n_656) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_590), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_577), .B(n_492), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_597), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_579), .B(n_396), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_607), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_578), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_578), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_607), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_588), .Y(n_665) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_578), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_613), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_657), .B(n_615), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_657), .Y(n_669) );
INVx5_ASAP7_75t_L g670 ( .A(n_620), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_659), .A2(n_611), .B1(n_606), .B2(n_597), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_659), .B(n_584), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_646), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_650), .B(n_383), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_633), .A2(n_654), .B1(n_623), .B2(n_644), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_623), .B(n_412), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_633), .A2(n_605), .B1(n_465), .B2(n_403), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_629), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_646), .Y(n_679) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_637), .B(n_590), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_646), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_633), .A2(n_465), .B1(n_403), .B2(n_449), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_649), .B(n_660), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_649), .B(n_579), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_649), .Y(n_685) );
BUFx8_ASAP7_75t_L g686 ( .A(n_644), .Y(n_686) );
INVx3_ASAP7_75t_L g687 ( .A(n_632), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_634), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_660), .B(n_582), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_660), .B(n_582), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_629), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_620), .A2(n_614), .B1(n_619), .B2(n_426), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_639), .B(n_592), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_645), .B(n_426), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_620), .A2(n_619), .B1(n_467), .B2(n_476), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_641), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_639), .B(n_592), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_641), .Y(n_698) );
HB1xp67_ASAP7_75t_SL g699 ( .A(n_638), .Y(n_699) );
NOR3xp33_ASAP7_75t_SL g700 ( .A(n_653), .B(n_454), .C(n_412), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_654), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_632), .A2(n_509), .B(n_490), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_635), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_634), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_661), .Y(n_705) );
INVx3_ASAP7_75t_L g706 ( .A(n_632), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_661), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_634), .Y(n_708) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_648), .B(n_408), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_634), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_664), .Y(n_711) );
INVx2_ASAP7_75t_SL g712 ( .A(n_639), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_650), .B(n_390), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_634), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_642), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_650), .B(n_391), .Y(n_716) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_650), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_626), .B(n_392), .Y(n_718) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_626), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_626), .B(n_398), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_626), .B(n_400), .Y(n_721) );
O2A1O1Ixp5_ASAP7_75t_L g722 ( .A1(n_632), .A2(n_429), .B(n_473), .C(n_410), .Y(n_722) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_643), .B(n_394), .Y(n_723) );
NAND2x1p5_ASAP7_75t_L g724 ( .A(n_642), .B(n_546), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_625), .B(n_454), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_642), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_626), .B(n_405), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_664), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_655), .B(n_419), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_620), .A2(n_467), .B1(n_476), .B2(n_456), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_653), .B(n_534), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_626), .B(n_407), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_655), .B(n_419), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_620), .A2(n_456), .B1(n_604), .B2(n_602), .Y(n_734) );
INVx2_ASAP7_75t_SL g735 ( .A(n_620), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_642), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_620), .A2(n_604), .B1(n_602), .B2(n_438), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_626), .B(n_409), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_665), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_655), .B(n_504), .Y(n_740) );
BUFx2_ASAP7_75t_L g741 ( .A(n_620), .Y(n_741) );
INVx1_ASAP7_75t_SL g742 ( .A(n_622), .Y(n_742) );
INVx3_ASAP7_75t_L g743 ( .A(n_647), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_665), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_642), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_648), .A2(n_442), .B1(n_487), .B2(n_384), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_625), .B(n_389), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_631), .B(n_411), .Y(n_748) );
BUFx12f_ASAP7_75t_L g749 ( .A(n_620), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_647), .A2(n_604), .B1(n_602), .B2(n_440), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_647), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_647), .B(n_593), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_655), .B(n_504), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_658), .A2(n_449), .B1(n_550), .B2(n_471), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_658), .B(n_531), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_621), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_667), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_621), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_624), .Y(n_759) );
BUFx3_ASAP7_75t_L g760 ( .A(n_631), .Y(n_760) );
INVxp67_ASAP7_75t_L g761 ( .A(n_656), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_631), .B(n_413), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_628), .B(n_593), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_667), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_683), .B(n_628), .Y(n_765) );
INVx1_ASAP7_75t_SL g766 ( .A(n_701), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_687), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_703), .Y(n_768) );
OAI22xp5_ASAP7_75t_SL g769 ( .A1(n_746), .A2(n_508), .B1(n_532), .B2(n_491), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_676), .B(n_491), .Y(n_770) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_749), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_669), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_754), .A2(n_508), .B1(n_552), .B2(n_532), .Y(n_773) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_749), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_687), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_687), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_699), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_673), .B(n_636), .Y(n_778) );
BUFx4f_ASAP7_75t_L g779 ( .A(n_724), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_706), .Y(n_780) );
BUFx4f_ASAP7_75t_L g781 ( .A(n_724), .Y(n_781) );
INVx1_ASAP7_75t_SL g782 ( .A(n_759), .Y(n_782) );
NOR2xp33_ASAP7_75t_SL g783 ( .A(n_670), .B(n_631), .Y(n_783) );
BUFx4f_ASAP7_75t_L g784 ( .A(n_688), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_674), .A2(n_631), .B(n_636), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_674), .A2(n_631), .B(n_640), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_686), .A2(n_552), .B1(n_471), .B2(n_550), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_709), .A2(n_640), .B1(n_627), .B2(n_624), .Y(n_788) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_670), .Y(n_789) );
INVx2_ASAP7_75t_SL g790 ( .A(n_686), .Y(n_790) );
AOI21xp33_ASAP7_75t_L g791 ( .A1(n_709), .A2(n_627), .B(n_561), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_715), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_673), .B(n_424), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_726), .Y(n_794) );
INVx3_ASAP7_75t_SL g795 ( .A(n_742), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_706), .Y(n_796) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_670), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_679), .A2(n_604), .B1(n_602), .B2(n_479), .Y(n_798) );
O2A1O1Ixp33_ASAP7_75t_SL g799 ( .A1(n_713), .A2(n_716), .B(n_720), .C(n_718), .Y(n_799) );
BUFx4f_ASAP7_75t_SL g800 ( .A(n_686), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_706), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_684), .B(n_543), .Y(n_802) );
BUFx2_ASAP7_75t_L g803 ( .A(n_682), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_681), .A2(n_483), .B1(n_484), .B2(n_474), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_745), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_684), .B(n_560), .Y(n_806) );
AOI21xp33_ASAP7_75t_L g807 ( .A1(n_685), .A2(n_486), .B(n_417), .Y(n_807) );
OAI22x1_ASAP7_75t_L g808 ( .A1(n_677), .A2(n_499), .B1(n_547), .B2(n_533), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_725), .A2(n_533), .B1(n_535), .B2(n_531), .Y(n_809) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_747), .A2(n_494), .B1(n_511), .B2(n_503), .C(n_485), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_684), .Y(n_811) );
AND2x4_ASAP7_75t_L g812 ( .A(n_680), .B(n_712), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_693), .B(n_535), .Y(n_813) );
BUFx8_ASAP7_75t_SL g814 ( .A(n_741), .Y(n_814) );
INVx4_ASAP7_75t_L g815 ( .A(n_670), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_722), .A2(n_513), .B(n_522), .C(n_519), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_692), .A2(n_528), .B1(n_529), .B2(n_524), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_704), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_763), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_671), .B(n_499), .Y(n_820) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_763), .Y(n_821) );
INVx4_ASAP7_75t_L g822 ( .A(n_693), .Y(n_822) );
O2A1O1Ixp5_ASAP7_75t_L g823 ( .A1(n_713), .A2(n_667), .B(n_453), .C(n_451), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_675), .B(n_599), .Y(n_824) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_717), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_694), .A2(n_555), .B1(n_530), .B2(n_539), .Y(n_826) );
OAI33xp33_ASAP7_75t_L g827 ( .A1(n_672), .A2(n_612), .A3(n_608), .B1(n_616), .B2(n_610), .B3(n_599), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_708), .Y(n_828) );
BUFx2_ASAP7_75t_L g829 ( .A(n_668), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_743), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_710), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_731), .A2(n_555), .B1(n_437), .B2(n_604), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_761), .B(n_537), .Y(n_833) );
INVx3_ASAP7_75t_L g834 ( .A(n_743), .Y(n_834) );
NOR2xp33_ASAP7_75t_SL g835 ( .A(n_735), .B(n_604), .Y(n_835) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_736), .Y(n_836) );
INVx2_ASAP7_75t_SL g837 ( .A(n_693), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_694), .B(n_608), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_729), .A2(n_423), .B(n_415), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_714), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_752), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_689), .A2(n_542), .B1(n_544), .B2(n_540), .Y(n_842) );
INVx3_ASAP7_75t_L g843 ( .A(n_743), .Y(n_843) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_733), .A2(n_428), .B(n_425), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_752), .Y(n_845) );
AO21x2_ASAP7_75t_L g846 ( .A1(n_740), .A2(n_431), .B(n_430), .Y(n_846) );
INVx3_ASAP7_75t_L g847 ( .A(n_751), .Y(n_847) );
AOI21xp5_ASAP7_75t_L g848 ( .A1(n_753), .A2(n_439), .B(n_435), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_751), .Y(n_849) );
OR2x6_ASAP7_75t_SL g850 ( .A(n_700), .B(n_434), .Y(n_850) );
NOR2xp33_ASAP7_75t_SL g851 ( .A(n_735), .B(n_604), .Y(n_851) );
BUFx6f_ASAP7_75t_L g852 ( .A(n_717), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_690), .B(n_548), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_697), .B(n_549), .Y(n_854) );
INVx1_ASAP7_75t_SL g855 ( .A(n_697), .Y(n_855) );
INVx4_ASAP7_75t_L g856 ( .A(n_697), .Y(n_856) );
OAI221xp5_ASAP7_75t_L g857 ( .A1(n_730), .A2(n_567), .B1(n_572), .B2(n_562), .C(n_551), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_751), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_702), .A2(n_444), .B(n_441), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_695), .B(n_610), .Y(n_860) );
A2O1A1Ixp33_ASAP7_75t_L g861 ( .A1(n_756), .A2(n_453), .B(n_452), .C(n_393), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_723), .B(n_612), .Y(n_862) );
INVx5_ASAP7_75t_L g863 ( .A(n_752), .Y(n_863) );
INVx3_ASAP7_75t_L g864 ( .A(n_678), .Y(n_864) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_717), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_678), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_758), .A2(n_618), .B1(n_616), .B2(n_447), .Y(n_867) );
CKINVDCx6p67_ASAP7_75t_R g868 ( .A(n_755), .Y(n_868) );
NAND2xp5_ASAP7_75t_SL g869 ( .A(n_717), .B(n_469), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_691), .B(n_618), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_734), .A2(n_448), .B1(n_450), .B2(n_445), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_691), .B(n_496), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g873 ( .A1(n_696), .A2(n_457), .B(n_455), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_696), .A2(n_460), .B(n_459), .Y(n_874) );
CKINVDCx16_ASAP7_75t_R g875 ( .A(n_760), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_737), .A2(n_463), .B1(n_466), .B2(n_462), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_698), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_705), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_705), .B(n_559), .Y(n_879) );
NOR2xp33_ASAP7_75t_R g880 ( .A(n_750), .B(n_475), .Y(n_880) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_739), .Y(n_881) );
BUFx2_ASAP7_75t_L g882 ( .A(n_739), .Y(n_882) );
OA21x2_ASAP7_75t_L g883 ( .A1(n_707), .A2(n_509), .B(n_490), .Y(n_883) );
OR2x6_ASAP7_75t_L g884 ( .A(n_707), .B(n_468), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_711), .B(n_427), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_711), .A2(n_604), .B(n_472), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_728), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_744), .B(n_520), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_744), .A2(n_468), .B1(n_477), .B2(n_557), .Y(n_889) );
INVx3_ASAP7_75t_L g890 ( .A(n_760), .Y(n_890) );
INVx3_ASAP7_75t_L g891 ( .A(n_719), .Y(n_891) );
INVx3_ASAP7_75t_L g892 ( .A(n_719), .Y(n_892) );
A2O1A1Ixp33_ASAP7_75t_SL g893 ( .A1(n_757), .A2(n_451), .B(n_591), .C(n_588), .Y(n_893) );
BUFx3_ASAP7_75t_L g894 ( .A(n_764), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_764), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_718), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_720), .A2(n_470), .B1(n_481), .B2(n_480), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_721), .Y(n_898) );
INVx3_ASAP7_75t_L g899 ( .A(n_719), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_721), .Y(n_900) );
INVxp67_ASAP7_75t_L g901 ( .A(n_727), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_727), .Y(n_902) );
BUFx2_ASAP7_75t_L g903 ( .A(n_719), .Y(n_903) );
BUFx2_ASAP7_75t_L g904 ( .A(n_732), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_732), .B(n_432), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_738), .B(n_514), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_738), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_748), .B(n_468), .Y(n_908) );
INVx4_ASAP7_75t_L g909 ( .A(n_748), .Y(n_909) );
O2A1O1Ixp33_ASAP7_75t_L g910 ( .A1(n_762), .A2(n_488), .B(n_489), .C(n_482), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_762), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g912 ( .A(n_722), .B(n_613), .C(n_477), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_683), .B(n_477), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_709), .A2(n_477), .B1(n_613), .B2(n_501), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_674), .A2(n_502), .B(n_493), .Y(n_915) );
AO31x2_ASAP7_75t_L g916 ( .A1(n_788), .A2(n_861), .A3(n_867), .B(n_816), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_772), .Y(n_917) );
OA21x2_ASAP7_75t_L g918 ( .A1(n_886), .A2(n_570), .B(n_563), .Y(n_918) );
NAND2x1p5_ASAP7_75t_L g919 ( .A(n_779), .B(n_506), .Y(n_919) );
OAI21xp33_ASAP7_75t_L g920 ( .A1(n_833), .A2(n_510), .B(n_507), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_819), .B(n_512), .Y(n_921) );
NAND2xp5_ASAP7_75t_SL g922 ( .A(n_825), .B(n_613), .Y(n_922) );
A2O1A1Ixp33_ASAP7_75t_L g923 ( .A1(n_791), .A2(n_570), .B(n_576), .C(n_563), .Y(n_923) );
CKINVDCx16_ASAP7_75t_R g924 ( .A(n_769), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_882), .Y(n_925) );
NAND2x1p5_ASAP7_75t_L g926 ( .A(n_779), .B(n_517), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_821), .A2(n_824), .B1(n_803), .B2(n_827), .Y(n_927) );
OAI21x1_ASAP7_75t_L g928 ( .A1(n_883), .A2(n_576), .B(n_523), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_766), .Y(n_929) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_912), .A2(n_525), .B(n_518), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_766), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_800), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_765), .B(n_527), .Y(n_933) );
O2A1O1Ixp33_ASAP7_75t_SL g934 ( .A1(n_893), .A2(n_541), .B(n_545), .C(n_538), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_788), .A2(n_844), .B(n_839), .Y(n_935) );
A2O1A1Ixp33_ASAP7_75t_L g936 ( .A1(n_791), .A2(n_558), .B(n_564), .C(n_553), .Y(n_936) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_912), .A2(n_566), .B(n_565), .Y(n_937) );
INVx6_ASAP7_75t_L g938 ( .A(n_863), .Y(n_938) );
AND2x4_ASAP7_75t_L g939 ( .A(n_782), .B(n_568), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_793), .Y(n_940) );
BUFx12f_ASAP7_75t_L g941 ( .A(n_777), .Y(n_941) );
INVx3_ASAP7_75t_L g942 ( .A(n_863), .Y(n_942) );
BUFx3_ASAP7_75t_L g943 ( .A(n_781), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_793), .A2(n_613), .B1(n_571), .B2(n_574), .Y(n_944) );
OA21x2_ASAP7_75t_L g945 ( .A1(n_886), .A2(n_575), .B(n_569), .Y(n_945) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_795), .Y(n_946) );
OAI21x1_ASAP7_75t_L g947 ( .A1(n_883), .A2(n_652), .B(n_651), .Y(n_947) );
OA21x2_ASAP7_75t_L g948 ( .A1(n_823), .A2(n_652), .B(n_651), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_782), .B(n_5), .Y(n_949) );
OA21x2_ASAP7_75t_L g950 ( .A1(n_914), .A2(n_662), .B(n_591), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_854), .Y(n_951) );
AO21x2_ASAP7_75t_L g952 ( .A1(n_846), .A2(n_594), .B(n_588), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_817), .A2(n_613), .B1(n_594), .B2(n_598), .Y(n_953) );
NOR4xp25_ASAP7_75t_L g954 ( .A(n_857), .B(n_595), .C(n_598), .D(n_594), .Y(n_954) );
CKINVDCx14_ASAP7_75t_R g955 ( .A(n_781), .Y(n_955) );
AO32x2_ASAP7_75t_L g956 ( .A1(n_871), .A2(n_580), .A3(n_600), .B1(n_598), .B2(n_595), .Y(n_956) );
OR2x2_ASAP7_75t_L g957 ( .A(n_770), .B(n_5), .Y(n_957) );
INVx2_ASAP7_75t_SL g958 ( .A(n_790), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_864), .Y(n_959) );
OA21x2_ASAP7_75t_L g960 ( .A1(n_848), .A2(n_662), .B(n_595), .Y(n_960) );
INVx3_ASAP7_75t_SL g961 ( .A(n_875), .Y(n_961) );
INVx2_ASAP7_75t_SL g962 ( .A(n_768), .Y(n_962) );
OAI21x1_ASAP7_75t_SL g963 ( .A1(n_778), .A2(n_6), .B(n_7), .Y(n_963) );
A2O1A1Ixp33_ASAP7_75t_L g964 ( .A1(n_853), .A2(n_600), .B(n_580), .C(n_630), .Y(n_964) );
OAI21x1_ASAP7_75t_L g965 ( .A1(n_913), .A2(n_600), .B(n_580), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_787), .Y(n_966) );
OA21x2_ASAP7_75t_L g967 ( .A1(n_859), .A2(n_600), .B(n_580), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_811), .Y(n_968) );
OAI21x1_ASAP7_75t_L g969 ( .A1(n_877), .A2(n_127), .B(n_125), .Y(n_969) );
OA21x2_ASAP7_75t_L g970 ( .A1(n_798), .A2(n_663), .B(n_630), .Y(n_970) );
OR2x2_ASAP7_75t_L g971 ( .A(n_773), .B(n_6), .Y(n_971) );
OAI21x1_ASAP7_75t_SL g972 ( .A1(n_878), .A2(n_8), .B(n_9), .Y(n_972) );
INVx8_ASAP7_75t_L g973 ( .A(n_863), .Y(n_973) );
NOR2x1_ASAP7_75t_SL g974 ( .A(n_884), .B(n_8), .Y(n_974) );
OA21x2_ASAP7_75t_L g975 ( .A1(n_908), .A2(n_874), .B(n_873), .Y(n_975) );
OAI21x1_ASAP7_75t_L g976 ( .A1(n_870), .A2(n_131), .B(n_129), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g977 ( .A1(n_855), .A2(n_12), .B1(n_10), .B2(n_11), .Y(n_977) );
NAND2xp33_ASAP7_75t_SL g978 ( .A(n_881), .B(n_10), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_806), .Y(n_979) );
OAI21x1_ASAP7_75t_L g980 ( .A1(n_891), .A2(n_136), .B(n_134), .Y(n_980) );
OAI21x1_ASAP7_75t_L g981 ( .A1(n_891), .A2(n_138), .B(n_137), .Y(n_981) );
OAI21x1_ASAP7_75t_L g982 ( .A1(n_892), .A2(n_145), .B(n_142), .Y(n_982) );
CKINVDCx14_ASAP7_75t_R g983 ( .A(n_769), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_817), .A2(n_663), .B1(n_666), .B2(n_630), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_866), .Y(n_985) );
OA21x2_ASAP7_75t_L g986 ( .A1(n_915), .A2(n_663), .B(n_630), .Y(n_986) );
AO21x2_ASAP7_75t_L g987 ( .A1(n_846), .A2(n_666), .B(n_663), .Y(n_987) );
OAI21x1_ASAP7_75t_L g988 ( .A1(n_892), .A2(n_149), .B(n_148), .Y(n_988) );
NAND2x1p5_ASAP7_75t_L g989 ( .A(n_822), .B(n_11), .Y(n_989) );
AND2x4_ASAP7_75t_L g990 ( .A(n_822), .B(n_13), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_802), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_838), .B(n_13), .Y(n_992) );
NAND2x1p5_ASAP7_75t_L g993 ( .A(n_856), .B(n_14), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_855), .A2(n_663), .B1(n_666), .B2(n_630), .Y(n_994) );
OAI21x1_ASAP7_75t_L g995 ( .A1(n_899), .A2(n_151), .B(n_150), .Y(n_995) );
OA21x2_ASAP7_75t_L g996 ( .A1(n_887), .A2(n_663), .B(n_630), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_802), .Y(n_997) );
OAI21x1_ASAP7_75t_L g998 ( .A1(n_785), .A2(n_157), .B(n_156), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_814), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_841), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1001 ( .A(n_784), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_856), .B(n_15), .Y(n_1002) );
AOI21xp5_ASAP7_75t_L g1003 ( .A1(n_786), .A2(n_663), .B(n_630), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_845), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_818), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_828), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_862), .A2(n_666), .B1(n_19), .B2(n_15), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_850), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_884), .A2(n_666), .B1(n_20), .B2(n_18), .Y(n_1009) );
INVx2_ASAP7_75t_L g1010 ( .A(n_792), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_837), .B(n_19), .Y(n_1011) );
OAI21x1_ASAP7_75t_L g1012 ( .A1(n_895), .A2(n_169), .B(n_164), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_868), .B(n_21), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_831), .Y(n_1014) );
AO21x2_ASAP7_75t_L g1015 ( .A1(n_876), .A2(n_666), .B(n_172), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_862), .A2(n_666), .B1(n_24), .B2(n_22), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_810), .A2(n_25), .B1(n_22), .B2(n_23), .Y(n_1017) );
OAI21x1_ASAP7_75t_L g1018 ( .A1(n_896), .A2(n_174), .B(n_170), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_840), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_794), .Y(n_1020) );
INVx1_ASAP7_75t_SL g1021 ( .A(n_879), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_835), .A2(n_180), .B(n_176), .Y(n_1022) );
INVx2_ASAP7_75t_L g1023 ( .A(n_805), .Y(n_1023) );
OAI21x1_ASAP7_75t_L g1024 ( .A1(n_898), .A2(n_185), .B(n_181), .Y(n_1024) );
OAI21x1_ASAP7_75t_L g1025 ( .A1(n_900), .A2(n_187), .B(n_186), .Y(n_1025) );
NAND2xp5_ASAP7_75t_SL g1026 ( .A(n_825), .B(n_189), .Y(n_1026) );
INVx3_ASAP7_75t_L g1027 ( .A(n_815), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_879), .Y(n_1028) );
OAI21xp5_ASAP7_75t_L g1029 ( .A1(n_871), .A2(n_25), .B(n_28), .Y(n_1029) );
AO21x2_ASAP7_75t_L g1030 ( .A1(n_876), .A2(n_191), .B(n_190), .Y(n_1030) );
OAI21x1_ASAP7_75t_L g1031 ( .A1(n_902), .A2(n_194), .B(n_192), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_829), .B(n_28), .Y(n_1032) );
OA21x2_ASAP7_75t_L g1033 ( .A1(n_860), .A2(n_196), .B(n_195), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_884), .Y(n_1034) );
OAI22xp33_ASAP7_75t_L g1035 ( .A1(n_867), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_812), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_812), .Y(n_1037) );
OAI21xp5_ASAP7_75t_L g1038 ( .A1(n_807), .A2(n_31), .B(n_32), .Y(n_1038) );
OAI21xp5_ASAP7_75t_L g1039 ( .A1(n_807), .A2(n_33), .B(n_35), .Y(n_1039) );
AO31x2_ASAP7_75t_L g1040 ( .A1(n_842), .A2(n_33), .A3(n_36), .B(n_37), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_809), .B(n_820), .Y(n_1041) );
OAI21x1_ASAP7_75t_L g1042 ( .A1(n_907), .A2(n_200), .B(n_199), .Y(n_1042) );
OAI21x1_ASAP7_75t_L g1043 ( .A1(n_890), .A2(n_203), .B(n_201), .Y(n_1043) );
OAI21x1_ASAP7_75t_L g1044 ( .A1(n_890), .A2(n_205), .B(n_204), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_842), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_1045) );
AO21x2_ASAP7_75t_L g1046 ( .A1(n_889), .A2(n_207), .B(n_206), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g1047 ( .A1(n_804), .A2(n_39), .B1(n_40), .B2(n_42), .Y(n_1047) );
BUFx4_ASAP7_75t_SL g1048 ( .A(n_911), .Y(n_1048) );
OAI21x1_ASAP7_75t_L g1049 ( .A1(n_767), .A2(n_210), .B(n_208), .Y(n_1049) );
OA21x2_ASAP7_75t_L g1050 ( .A1(n_885), .A2(n_215), .B(n_212), .Y(n_1050) );
AND2x4_ASAP7_75t_L g1051 ( .A(n_771), .B(n_39), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_872), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_804), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_826), .B(n_45), .Y(n_1054) );
OAI21x1_ASAP7_75t_L g1055 ( .A1(n_775), .A2(n_218), .B(n_216), .Y(n_1055) );
OAI21x1_ASAP7_75t_L g1056 ( .A1(n_776), .A2(n_222), .B(n_219), .Y(n_1056) );
OAI21x1_ASAP7_75t_L g1057 ( .A1(n_780), .A2(n_225), .B(n_223), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_813), .Y(n_1058) );
OAI21x1_ASAP7_75t_L g1059 ( .A1(n_801), .A2(n_228), .B(n_226), .Y(n_1059) );
OA21x2_ASAP7_75t_L g1060 ( .A1(n_888), .A2(n_232), .B(n_231), .Y(n_1060) );
AOI21x1_ASAP7_75t_L g1061 ( .A1(n_869), .A2(n_238), .B(n_234), .Y(n_1061) );
OAI21x1_ASAP7_75t_L g1062 ( .A1(n_830), .A2(n_240), .B(n_239), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_836), .Y(n_1063) );
A2O1A1Ixp33_ASAP7_75t_L g1064 ( .A1(n_910), .A2(n_45), .B(n_46), .C(n_47), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_825), .Y(n_1065) );
OAI21x1_ASAP7_75t_L g1066 ( .A1(n_849), .A2(n_246), .B(n_242), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_808), .B(n_47), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_858), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_796), .Y(n_1069) );
OA21x2_ASAP7_75t_L g1070 ( .A1(n_897), .A2(n_249), .B(n_247), .Y(n_1070) );
O2A1O1Ixp33_ASAP7_75t_SL g1071 ( .A1(n_901), .A2(n_252), .B(n_381), .C(n_378), .Y(n_1071) );
AOI21xp5_ASAP7_75t_SL g1072 ( .A1(n_852), .A2(n_382), .B(n_254), .Y(n_1072) );
OAI21x1_ASAP7_75t_L g1073 ( .A1(n_796), .A2(n_377), .B(n_375), .Y(n_1073) );
OR2x6_ASAP7_75t_L g1074 ( .A(n_771), .B(n_48), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_894), .Y(n_1075) );
OAI21x1_ASAP7_75t_L g1076 ( .A1(n_834), .A2(n_373), .B(n_371), .Y(n_1076) );
INVx1_ASAP7_75t_SL g1077 ( .A(n_903), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_834), .B(n_48), .Y(n_1078) );
INVx4_ASAP7_75t_L g1079 ( .A(n_771), .Y(n_1079) );
INVx4_ASAP7_75t_L g1080 ( .A(n_774), .Y(n_1080) );
INVx2_ASAP7_75t_SL g1081 ( .A(n_784), .Y(n_1081) );
AOI21x1_ASAP7_75t_L g1082 ( .A1(n_904), .A2(n_370), .B(n_369), .Y(n_1082) );
NAND2x1p5_ASAP7_75t_L g1083 ( .A(n_774), .B(n_49), .Y(n_1083) );
AO21x2_ASAP7_75t_L g1084 ( .A1(n_799), .A2(n_366), .B(n_364), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_843), .Y(n_1085) );
A2O1A1Ixp33_ASAP7_75t_L g1086 ( .A1(n_905), .A2(n_50), .B(n_51), .C(n_52), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1087 ( .A1(n_906), .A2(n_50), .B1(n_51), .B2(n_52), .C(n_53), .Y(n_1087) );
OAI21xp5_ASAP7_75t_L g1088 ( .A1(n_832), .A2(n_54), .B(n_55), .Y(n_1088) );
AO31x2_ASAP7_75t_L g1089 ( .A1(n_909), .A2(n_54), .A3(n_55), .B(n_56), .Y(n_1089) );
NAND2x1p5_ASAP7_75t_L g1090 ( .A(n_774), .B(n_57), .Y(n_1090) );
NAND2xp33_ASAP7_75t_R g1091 ( .A(n_880), .B(n_58), .Y(n_1091) );
OA21x2_ASAP7_75t_L g1092 ( .A1(n_865), .A2(n_363), .B(n_360), .Y(n_1092) );
OAI21x1_ASAP7_75t_L g1093 ( .A1(n_947), .A2(n_847), .B(n_843), .Y(n_1093) );
AOI22xp33_ASAP7_75t_SL g1094 ( .A1(n_983), .A2(n_835), .B1(n_851), .B2(n_847), .Y(n_1094) );
OR2x6_ASAP7_75t_L g1095 ( .A(n_943), .B(n_815), .Y(n_1095) );
AOI221xp5_ASAP7_75t_L g1096 ( .A1(n_1052), .A2(n_909), .B1(n_852), .B2(n_797), .C(n_789), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_955), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_983), .A2(n_852), .B1(n_797), .B2(n_789), .Y(n_1098) );
AOI222xp33_ASAP7_75t_L g1099 ( .A1(n_966), .A2(n_851), .B1(n_797), .B2(n_789), .C1(n_783), .C2(n_63), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g1100 ( .A1(n_1058), .A2(n_783), .B1(n_60), .B2(n_61), .C(n_62), .Y(n_1100) );
NAND2xp5_ASAP7_75t_SL g1101 ( .A(n_919), .B(n_59), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_927), .B(n_59), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_929), .Y(n_1103) );
OAI21x1_ASAP7_75t_L g1104 ( .A1(n_965), .A2(n_356), .B(n_355), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_931), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_917), .Y(n_1106) );
NAND2x1p5_ASAP7_75t_L g1107 ( .A(n_943), .B(n_60), .Y(n_1107) );
AOI221xp5_ASAP7_75t_L g1108 ( .A1(n_951), .A2(n_61), .B1(n_62), .B2(n_64), .C(n_65), .Y(n_1108) );
OAI211xp5_ASAP7_75t_L g1109 ( .A1(n_1017), .A2(n_64), .B(n_65), .C(n_66), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_1041), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_955), .B(n_68), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_924), .A2(n_69), .B1(n_70), .B2(n_71), .Y(n_1112) );
OAI21xp5_ASAP7_75t_L g1113 ( .A1(n_935), .A2(n_71), .B(n_72), .Y(n_1113) );
OAI221xp5_ASAP7_75t_L g1114 ( .A1(n_957), .A2(n_73), .B1(n_74), .B2(n_75), .C(n_76), .Y(n_1114) );
OAI221xp5_ASAP7_75t_L g1115 ( .A1(n_927), .A2(n_73), .B1(n_75), .B2(n_78), .C(n_79), .Y(n_1115) );
AOI21xp5_ASAP7_75t_L g1116 ( .A1(n_935), .A2(n_263), .B(n_352), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_925), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_1091), .A2(n_78), .B1(n_80), .B2(n_81), .Y(n_1118) );
AO21x2_ASAP7_75t_L g1119 ( .A1(n_964), .A2(n_264), .B(n_351), .Y(n_1119) );
OAI211xp5_ASAP7_75t_L g1120 ( .A1(n_1017), .A2(n_80), .B(n_82), .C(n_83), .Y(n_1120) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_1003), .A2(n_268), .B(n_348), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g1122 ( .A1(n_1091), .A2(n_82), .B1(n_84), .B2(n_85), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_1021), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g1124 ( .A(n_973), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_978), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_971), .A2(n_88), .B1(n_89), .B2(n_90), .Y(n_1126) );
AND2x4_ASAP7_75t_SL g1127 ( .A(n_932), .B(n_89), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_979), .B(n_90), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1028), .B(n_91), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1130 ( .A1(n_948), .A2(n_276), .B(n_345), .Y(n_1130) );
AOI22xp5_ASAP7_75t_L g1131 ( .A1(n_949), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_940), .B(n_92), .Y(n_1132) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1010), .Y(n_1133) );
CKINVDCx8_ASAP7_75t_R g1134 ( .A(n_946), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1020), .Y(n_1135) );
OA21x2_ASAP7_75t_L g1136 ( .A1(n_928), .A2(n_277), .B(n_342), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_991), .B(n_93), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_978), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_997), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1023), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_949), .A2(n_939), .B1(n_1002), .B2(n_990), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1005), .B(n_95), .Y(n_1142) );
A2O1A1Ixp33_ASAP7_75t_L g1143 ( .A1(n_1088), .A2(n_97), .B(n_98), .C(n_99), .Y(n_1143) );
AOI22xp33_ASAP7_75t_SL g1144 ( .A1(n_1074), .A2(n_99), .B1(n_100), .B2(n_103), .Y(n_1144) );
OAI221xp5_ASAP7_75t_SL g1145 ( .A1(n_1053), .A2(n_103), .B1(n_104), .B2(n_105), .C(n_106), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_962), .B(n_961), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_919), .B(n_104), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_989), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_1029), .A2(n_105), .B1(n_107), .B2(n_108), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_990), .A2(n_107), .B1(n_108), .B2(n_109), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_989), .Y(n_1151) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_1074), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_926), .B(n_110), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1006), .B(n_111), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_993), .Y(n_1155) );
OAI22xp33_ASAP7_75t_L g1156 ( .A1(n_1074), .A2(n_111), .B1(n_113), .B2(n_115), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_1002), .A2(n_113), .B1(n_115), .B2(n_116), .Y(n_1157) );
NOR2x1_ASAP7_75t_SL g1158 ( .A(n_1079), .B(n_116), .Y(n_1158) );
A2O1A1Ixp33_ASAP7_75t_L g1159 ( .A1(n_1088), .A2(n_118), .B(n_119), .C(n_120), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_993), .Y(n_1160) );
OAI221xp5_ASAP7_75t_SL g1161 ( .A1(n_1053), .A2(n_118), .B1(n_120), .B2(n_253), .C(n_257), .Y(n_1161) );
OA21x2_ASAP7_75t_L g1162 ( .A1(n_964), .A2(n_259), .B(n_260), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1014), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_939), .A2(n_269), .B1(n_270), .B2(n_272), .Y(n_1164) );
INVx2_ASAP7_75t_L g1165 ( .A(n_985), .Y(n_1165) );
OA21x2_ASAP7_75t_L g1166 ( .A1(n_976), .A2(n_279), .B(n_282), .Y(n_1166) );
INVx1_ASAP7_75t_SL g1167 ( .A(n_1077), .Y(n_1167) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1019), .Y(n_1168) );
AOI21xp5_ASAP7_75t_L g1169 ( .A1(n_948), .A2(n_286), .B(n_287), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1036), .B(n_288), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1000), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1063), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_992), .A2(n_291), .B1(n_292), .B2(n_293), .Y(n_1173) );
AO21x1_ASAP7_75t_L g1174 ( .A1(n_1029), .A2(n_294), .B(n_297), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_961), .B(n_298), .Y(n_1175) );
AOI21xp5_ASAP7_75t_L g1176 ( .A1(n_948), .A2(n_300), .B(n_301), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_936), .B(n_353), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_1054), .A2(n_310), .B1(n_317), .B2(n_319), .Y(n_1178) );
AND2x4_ASAP7_75t_L g1179 ( .A(n_1037), .B(n_321), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_992), .A2(n_936), .B1(n_921), .B2(n_933), .Y(n_1180) );
OAI22xp5_ASAP7_75t_SL g1181 ( .A1(n_926), .A2(n_322), .B1(n_325), .B2(n_327), .Y(n_1181) );
NAND3xp33_ASAP7_75t_L g1182 ( .A(n_923), .B(n_329), .C(n_332), .Y(n_1182) );
AOI21xp5_ASAP7_75t_L g1183 ( .A1(n_934), .A2(n_333), .B(n_334), .Y(n_1183) );
OR2x6_ASAP7_75t_L g1184 ( .A(n_973), .B(n_335), .Y(n_1184) );
OAI22xp33_ASAP7_75t_L g1185 ( .A1(n_1054), .A2(n_336), .B1(n_337), .B2(n_338), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_932), .Y(n_1186) );
OAI22xp5_ASAP7_75t_SL g1187 ( .A1(n_1047), .A2(n_339), .B1(n_999), .B2(n_1008), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_958), .B(n_1001), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_923), .A2(n_1007), .B1(n_1016), .B2(n_933), .Y(n_1189) );
OAI211xp5_ASAP7_75t_SL g1190 ( .A1(n_1067), .A2(n_1047), .B(n_921), .C(n_1087), .Y(n_1190) );
BUFx6f_ASAP7_75t_L g1191 ( .A(n_973), .Y(n_1191) );
NOR2xp33_ASAP7_75t_L g1192 ( .A(n_1081), .B(n_968), .Y(n_1192) );
BUFx8_ASAP7_75t_L g1193 ( .A(n_941), .Y(n_1193) );
NAND3xp33_ASAP7_75t_L g1194 ( .A(n_1064), .B(n_1087), .C(n_984), .Y(n_1194) );
AOI21xp5_ASAP7_75t_L g1195 ( .A1(n_934), .A2(n_994), .B(n_960), .Y(n_1195) );
OAI211xp5_ASAP7_75t_L g1196 ( .A1(n_1045), .A2(n_1016), .B(n_1007), .C(n_920), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1013), .B(n_1045), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_944), .A2(n_1032), .B1(n_1051), .B2(n_1035), .Y(n_1198) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_944), .A2(n_1032), .B1(n_1051), .B2(n_1035), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1004), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1079), .B(n_1080), .Y(n_1201) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_1011), .A2(n_999), .B1(n_1009), .B2(n_1080), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1040), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1068), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_916), .B(n_1011), .Y(n_1205) );
INVx2_ASAP7_75t_L g1206 ( .A(n_959), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_916), .B(n_1075), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_1038), .A2(n_1039), .B1(n_1078), .B2(n_938), .Y(n_1208) );
AOI21xp5_ASAP7_75t_L g1209 ( .A1(n_960), .A2(n_922), .B(n_986), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_942), .B(n_1078), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_1009), .A2(n_984), .B1(n_1090), .B2(n_1083), .Y(n_1211) );
OAI21xp5_ASAP7_75t_L g1212 ( .A1(n_930), .A2(n_937), .B(n_954), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_952), .Y(n_1213) );
AOI21xp33_ASAP7_75t_SL g1214 ( .A1(n_977), .A2(n_1090), .B(n_1083), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1215 ( .A(n_942), .B(n_938), .Y(n_1215) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_1038), .A2(n_1039), .B1(n_977), .B2(n_1086), .C(n_1064), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1048), .Y(n_1217) );
OR2x6_ASAP7_75t_L g1218 ( .A(n_938), .B(n_963), .Y(n_1218) );
AND2x4_ASAP7_75t_L g1219 ( .A(n_1027), .B(n_1069), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1040), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_952), .Y(n_1221) );
HB1xp67_ASAP7_75t_L g1222 ( .A(n_1048), .Y(n_1222) );
AOI21xp5_ASAP7_75t_L g1223 ( .A1(n_922), .A2(n_986), .B(n_930), .Y(n_1223) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_1027), .B(n_1085), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_1086), .A2(n_1034), .B1(n_953), .B2(n_937), .Y(n_1225) );
OAI22xp5_ASAP7_75t_SL g1226 ( .A1(n_1070), .A2(n_1050), .B1(n_1033), .B2(n_945), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_972), .A2(n_953), .B1(n_975), .B2(n_945), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_916), .B(n_1040), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1065), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_918), .A2(n_1065), .B1(n_975), .B2(n_1022), .Y(n_1230) );
AO21x2_ASAP7_75t_L g1231 ( .A1(n_987), .A2(n_1015), .B(n_1084), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_1030), .A2(n_987), .B1(n_918), .B2(n_1046), .Y(n_1232) );
AOI21xp5_ASAP7_75t_L g1233 ( .A1(n_918), .A2(n_1050), .B(n_996), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_1022), .A2(n_1070), .B1(n_1033), .B2(n_1060), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_967), .Y(n_1235) );
OAI222xp33_ASAP7_75t_L g1236 ( .A1(n_1026), .A2(n_1082), .B1(n_1061), .B2(n_974), .C1(n_1040), .C2(n_1089), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_916), .B(n_1089), .Y(n_1237) );
AOI221x1_ASAP7_75t_SL g1238 ( .A1(n_1089), .A2(n_1030), .B1(n_956), .B2(n_1046), .C(n_1071), .Y(n_1238) );
OAI211xp5_ASAP7_75t_L g1239 ( .A1(n_1071), .A2(n_1072), .B(n_1092), .C(n_1060), .Y(n_1239) );
BUFx12f_ASAP7_75t_L g1240 ( .A(n_1089), .Y(n_1240) );
OA21x2_ASAP7_75t_L g1241 ( .A1(n_1018), .A2(n_1055), .B(n_1066), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1242 ( .A1(n_1026), .A2(n_950), .B1(n_967), .B2(n_970), .C(n_1092), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_956), .Y(n_1243) );
OAI21xp5_ASAP7_75t_L g1244 ( .A1(n_998), .A2(n_1056), .B(n_1062), .Y(n_1244) );
AO31x2_ASAP7_75t_L g1245 ( .A1(n_956), .A2(n_1015), .A3(n_1084), .B(n_967), .Y(n_1245) );
NAND3xp33_ASAP7_75t_L g1246 ( .A(n_950), .B(n_970), .C(n_956), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_1043), .A2(n_1044), .B1(n_969), .B2(n_981), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_980), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_982), .B(n_988), .Y(n_1249) );
OAI221xp5_ASAP7_75t_L g1250 ( .A1(n_1049), .A2(n_1059), .B1(n_1057), .B2(n_1024), .C(n_1025), .Y(n_1250) );
INVx4_ASAP7_75t_L g1251 ( .A(n_995), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1076), .B(n_1073), .Y(n_1252) );
AOI21xp5_ASAP7_75t_L g1253 ( .A1(n_1012), .A2(n_1031), .B(n_1042), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_983), .A2(n_769), .B1(n_803), .B2(n_1041), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_983), .A2(n_769), .B1(n_803), .B2(n_1041), .Y(n_1255) );
OAI22xp33_ASAP7_75t_L g1256 ( .A1(n_924), .A2(n_754), .B1(n_800), .B2(n_1091), .Y(n_1256) );
INVx2_ASAP7_75t_SL g1257 ( .A(n_943), .Y(n_1257) );
AOI221xp5_ASAP7_75t_L g1258 ( .A1(n_1052), .A2(n_773), .B1(n_833), .B2(n_810), .C(n_769), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_983), .A2(n_769), .B1(n_803), .B2(n_1041), .Y(n_1259) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_1052), .A2(n_675), .B1(n_787), .B2(n_682), .C(n_746), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_955), .B(n_659), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_983), .A2(n_769), .B1(n_803), .B2(n_1041), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1172), .Y(n_1263) );
BUFx2_ASAP7_75t_SL g1264 ( .A(n_1134), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1106), .Y(n_1265) );
HB1xp67_ASAP7_75t_L g1266 ( .A(n_1235), .Y(n_1266) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1213), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1133), .B(n_1135), .Y(n_1268) );
NOR2x1_ASAP7_75t_L g1269 ( .A(n_1184), .B(n_1175), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1163), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1140), .B(n_1165), .Y(n_1271) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1221), .Y(n_1272) );
INVx3_ASAP7_75t_L g1273 ( .A(n_1124), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1261), .B(n_1147), .Y(n_1274) );
NOR3xp33_ASAP7_75t_L g1275 ( .A(n_1187), .B(n_1190), .C(n_1256), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1258), .B(n_1197), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1153), .B(n_1111), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_1167), .B(n_1204), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1167), .B(n_1254), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1255), .B(n_1259), .Y(n_1280) );
NOR2x1_ASAP7_75t_L g1281 ( .A(n_1184), .B(n_1156), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g1282 ( .A(n_1229), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1117), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1168), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1262), .B(n_1124), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1124), .B(n_1191), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1191), .B(n_1201), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1103), .Y(n_1288) );
NAND2xp33_ASAP7_75t_SL g1289 ( .A(n_1211), .B(n_1149), .Y(n_1289) );
OAI222xp33_ASAP7_75t_L g1290 ( .A1(n_1141), .A2(n_1149), .B1(n_1118), .B2(n_1199), .C1(n_1198), .C2(n_1107), .Y(n_1290) );
INVx2_ASAP7_75t_SL g1291 ( .A(n_1191), .Y(n_1291) );
AND2x4_ASAP7_75t_L g1292 ( .A(n_1148), .B(n_1151), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1105), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1237), .B(n_1171), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1200), .B(n_1113), .Y(n_1295) );
BUFx2_ASAP7_75t_L g1296 ( .A(n_1184), .Y(n_1296) );
AO21x2_ASAP7_75t_L g1297 ( .A1(n_1233), .A2(n_1195), .B(n_1209), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1139), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1113), .B(n_1206), .Y(n_1299) );
NOR2x1_ASAP7_75t_L g1300 ( .A(n_1122), .B(n_1101), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g1301 ( .A(n_1210), .Y(n_1301) );
AO31x2_ASAP7_75t_L g1302 ( .A1(n_1228), .A2(n_1234), .A3(n_1230), .B(n_1220), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1180), .B(n_1203), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1207), .B(n_1205), .Y(n_1304) );
AOI21xp5_ASAP7_75t_SL g1305 ( .A1(n_1234), .A2(n_1179), .B(n_1170), .Y(n_1305) );
NOR2x1_ASAP7_75t_L g1306 ( .A(n_1155), .B(n_1160), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1307 ( .A(n_1146), .B(n_1097), .Y(n_1307) );
OAI21xp5_ASAP7_75t_L g1308 ( .A1(n_1196), .A2(n_1194), .B(n_1189), .Y(n_1308) );
AO31x2_ASAP7_75t_L g1309 ( .A1(n_1174), .A2(n_1243), .A3(n_1251), .B(n_1248), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1170), .B(n_1179), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1142), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1154), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1102), .B(n_1144), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1107), .Y(n_1314) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_1240), .Y(n_1315) );
INVx2_ASAP7_75t_SL g1316 ( .A(n_1095), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1257), .B(n_1202), .Y(n_1317) );
INVx2_ASAP7_75t_SL g1318 ( .A(n_1095), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1128), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1152), .B(n_1260), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1192), .B(n_1126), .Y(n_1321) );
INVx2_ASAP7_75t_SL g1322 ( .A(n_1095), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1186), .B(n_1129), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1189), .B(n_1137), .Y(n_1324) );
OAI222xp33_ASAP7_75t_L g1325 ( .A1(n_1145), .A2(n_1161), .B1(n_1131), .B2(n_1100), .C1(n_1114), .C2(n_1125), .Y(n_1325) );
INVxp67_ASAP7_75t_L g1326 ( .A(n_1188), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1132), .B(n_1216), .Y(n_1327) );
BUFx2_ASAP7_75t_L g1328 ( .A(n_1217), .Y(n_1328) );
OAI22xp33_ASAP7_75t_L g1329 ( .A1(n_1194), .A2(n_1115), .B1(n_1214), .B2(n_1225), .Y(n_1329) );
NOR2xp67_ASAP7_75t_L g1330 ( .A(n_1222), .B(n_1215), .Y(n_1330) );
BUFx2_ASAP7_75t_L g1331 ( .A(n_1218), .Y(n_1331) );
INVx2_ASAP7_75t_SL g1332 ( .A(n_1224), .Y(n_1332) );
BUFx6f_ASAP7_75t_L g1333 ( .A(n_1093), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1158), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1224), .B(n_1159), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1123), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1143), .B(n_1138), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1109), .Y(n_1338) );
INVx3_ASAP7_75t_L g1339 ( .A(n_1218), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1219), .B(n_1150), .Y(n_1340) );
OAI21xp5_ASAP7_75t_L g1341 ( .A1(n_1208), .A2(n_1212), .B(n_1227), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1219), .B(n_1157), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1110), .B(n_1108), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1127), .B(n_1112), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1120), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1187), .B(n_1099), .Y(n_1346) );
BUFx12f_ASAP7_75t_L g1347 ( .A(n_1193), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1177), .B(n_1098), .Y(n_1348) );
NOR2xp33_ASAP7_75t_L g1349 ( .A(n_1236), .B(n_1218), .Y(n_1349) );
HB1xp67_ASAP7_75t_L g1350 ( .A(n_1246), .Y(n_1350) );
INVx3_ASAP7_75t_SL g1351 ( .A(n_1193), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1181), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1181), .Y(n_1353) );
BUFx3_ASAP7_75t_L g1354 ( .A(n_1104), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1099), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1119), .Y(n_1356) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_1246), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1119), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1212), .B(n_1096), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1164), .B(n_1178), .Y(n_1360) );
OR2x2_ASAP7_75t_L g1361 ( .A(n_1182), .B(n_1173), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1238), .B(n_1094), .Y(n_1362) );
AND2x4_ASAP7_75t_SL g1363 ( .A(n_1251), .B(n_1252), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1182), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1249), .Y(n_1365) );
AND2x4_ASAP7_75t_L g1366 ( .A(n_1116), .B(n_1121), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1238), .B(n_1185), .Y(n_1367) );
INVx2_ASAP7_75t_L g1368 ( .A(n_1136), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1162), .B(n_1223), .Y(n_1369) );
BUFx2_ASAP7_75t_L g1370 ( .A(n_1162), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1232), .B(n_1231), .Y(n_1371) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1245), .Y(n_1372) );
HB1xp67_ASAP7_75t_L g1373 ( .A(n_1245), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1231), .B(n_1245), .Y(n_1374) );
OAI21xp5_ASAP7_75t_L g1375 ( .A1(n_1183), .A2(n_1253), .B(n_1130), .Y(n_1375) );
HB1xp67_ASAP7_75t_L g1376 ( .A(n_1242), .Y(n_1376) );
NAND3xp33_ASAP7_75t_L g1377 ( .A(n_1169), .B(n_1176), .C(n_1247), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1378 ( .A(n_1166), .B(n_1226), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1166), .B(n_1226), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1244), .B(n_1241), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1241), .Y(n_1381) );
INVx3_ASAP7_75t_L g1382 ( .A(n_1239), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1244), .B(n_1250), .Y(n_1383) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1235), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1261), .B(n_659), .Y(n_1385) );
INVx2_ASAP7_75t_L g1386 ( .A(n_1235), .Y(n_1386) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1235), .Y(n_1387) );
BUFx6f_ASAP7_75t_L g1388 ( .A(n_1124), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1172), .Y(n_1389) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1235), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1172), .Y(n_1391) );
INVxp67_ASAP7_75t_L g1392 ( .A(n_1261), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1133), .B(n_1135), .Y(n_1393) );
INVx2_ASAP7_75t_L g1394 ( .A(n_1235), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1172), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1294), .B(n_1304), .Y(n_1396) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_1275), .A2(n_1290), .B1(n_1276), .B2(n_1308), .C(n_1346), .Y(n_1397) );
INVx3_ASAP7_75t_L g1398 ( .A(n_1363), .Y(n_1398) );
INVx2_ASAP7_75t_L g1399 ( .A(n_1384), .Y(n_1399) );
OAI21xp33_ASAP7_75t_L g1400 ( .A1(n_1281), .A2(n_1280), .B(n_1352), .Y(n_1400) );
INVx2_ASAP7_75t_SL g1401 ( .A(n_1363), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1294), .B(n_1304), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1268), .B(n_1393), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1303), .B(n_1266), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1303), .B(n_1266), .Y(n_1405) );
BUFx3_ASAP7_75t_L g1406 ( .A(n_1286), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1365), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1386), .B(n_1387), .Y(n_1408) );
INVx4_ASAP7_75t_L g1409 ( .A(n_1296), .Y(n_1409) );
NAND3xp33_ASAP7_75t_L g1410 ( .A(n_1353), .B(n_1300), .C(n_1334), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1386), .Y(n_1411) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_1282), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1387), .Y(n_1413) );
INVx4_ASAP7_75t_L g1414 ( .A(n_1310), .Y(n_1414) );
AO21x2_ASAP7_75t_L g1415 ( .A1(n_1383), .A2(n_1375), .B(n_1368), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1390), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1390), .B(n_1394), .Y(n_1417) );
AND2x4_ASAP7_75t_L g1418 ( .A(n_1339), .B(n_1315), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1394), .B(n_1282), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_1310), .A2(n_1305), .B1(n_1269), .B2(n_1355), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1268), .B(n_1393), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1267), .Y(n_1422) );
AOI33xp33_ASAP7_75t_L g1423 ( .A1(n_1279), .A2(n_1385), .A3(n_1319), .B1(n_1311), .B2(n_1312), .B3(n_1274), .Y(n_1423) );
INVx2_ASAP7_75t_SL g1424 ( .A(n_1388), .Y(n_1424) );
AOI221xp5_ASAP7_75t_SL g1425 ( .A1(n_1326), .A2(n_1392), .B1(n_1321), .B2(n_1344), .C(n_1329), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1341), .B(n_1271), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1272), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1272), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1271), .B(n_1295), .Y(n_1429) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1301), .B(n_1278), .Y(n_1430) );
NOR2xp67_ASAP7_75t_L g1431 ( .A(n_1347), .B(n_1315), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1381), .Y(n_1432) );
AOI221xp5_ASAP7_75t_L g1433 ( .A1(n_1329), .A2(n_1289), .B1(n_1336), .B2(n_1327), .C(n_1345), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1373), .Y(n_1434) );
BUFx2_ASAP7_75t_L g1435 ( .A(n_1339), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1295), .B(n_1299), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1299), .B(n_1371), .Y(n_1437) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1263), .Y(n_1438) );
OR2x2_ASAP7_75t_L g1439 ( .A(n_1301), .B(n_1317), .Y(n_1439) );
AOI22xp33_ASAP7_75t_SL g1440 ( .A1(n_1314), .A2(n_1340), .B1(n_1342), .B2(n_1331), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1371), .B(n_1284), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1373), .Y(n_1442) );
INVx2_ASAP7_75t_L g1443 ( .A(n_1372), .Y(n_1443) );
INVx2_ASAP7_75t_L g1444 ( .A(n_1380), .Y(n_1444) );
AOI221xp5_ASAP7_75t_L g1445 ( .A1(n_1289), .A2(n_1338), .B1(n_1325), .B2(n_1313), .C(n_1324), .Y(n_1445) );
BUFx3_ASAP7_75t_L g1446 ( .A(n_1388), .Y(n_1446) );
INVxp67_ASAP7_75t_L g1447 ( .A(n_1287), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1265), .B(n_1270), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1288), .B(n_1293), .Y(n_1449) );
HB1xp67_ASAP7_75t_L g1450 ( .A(n_1330), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1374), .B(n_1298), .Y(n_1451) );
BUFx2_ASAP7_75t_L g1452 ( .A(n_1339), .Y(n_1452) );
BUFx3_ASAP7_75t_L g1453 ( .A(n_1388), .Y(n_1453) );
NAND2xp5_ASAP7_75t_L g1454 ( .A(n_1389), .B(n_1395), .Y(n_1454) );
HB1xp67_ASAP7_75t_L g1455 ( .A(n_1292), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1391), .B(n_1283), .Y(n_1456) );
NOR3xp33_ASAP7_75t_SL g1457 ( .A(n_1351), .B(n_1347), .C(n_1343), .Y(n_1457) );
INVx1_ASAP7_75t_SL g1458 ( .A(n_1264), .Y(n_1458) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1362), .B(n_1320), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1374), .B(n_1305), .Y(n_1460) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1350), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_1277), .B(n_1313), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1350), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1302), .B(n_1357), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1285), .B(n_1292), .Y(n_1465) );
HB1xp67_ASAP7_75t_L g1466 ( .A(n_1292), .Y(n_1466) );
INVx3_ASAP7_75t_L g1467 ( .A(n_1382), .Y(n_1467) );
OR2x6_ASAP7_75t_SL g1468 ( .A(n_1367), .B(n_1379), .Y(n_1468) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_1332), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1302), .B(n_1357), .Y(n_1470) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1302), .Y(n_1471) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1302), .Y(n_1472) );
AOI22xp5_ASAP7_75t_L g1473 ( .A1(n_1340), .A2(n_1342), .B1(n_1337), .B2(n_1335), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1376), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1475 ( .A1(n_1337), .A2(n_1335), .B1(n_1360), .B2(n_1328), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1376), .B(n_1349), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1323), .B(n_1307), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1309), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1309), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1309), .Y(n_1480) );
HB1xp67_ASAP7_75t_L g1481 ( .A(n_1332), .Y(n_1481) );
INVx2_ASAP7_75t_L g1482 ( .A(n_1297), .Y(n_1482) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1309), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1306), .Y(n_1484) );
INVxp67_ASAP7_75t_L g1485 ( .A(n_1291), .Y(n_1485) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1448), .Y(n_1486) );
OR2x2_ASAP7_75t_L g1487 ( .A(n_1396), .B(n_1316), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1396), .B(n_1316), .Y(n_1488) );
OR2x2_ASAP7_75t_L g1489 ( .A(n_1402), .B(n_1318), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1448), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1491 ( .A(n_1402), .B(n_1318), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1447), .B(n_1291), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1406), .B(n_1322), .Y(n_1493) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1432), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_1397), .A2(n_1359), .B1(n_1349), .B2(n_1348), .Y(n_1495) );
AND2x4_ASAP7_75t_L g1496 ( .A(n_1460), .B(n_1382), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1430), .B(n_1322), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1449), .B(n_1273), .Y(n_1498) );
NAND5xp2_ASAP7_75t_SL g1499 ( .A(n_1445), .B(n_1351), .C(n_1273), .D(n_1388), .E(n_1382), .Y(n_1499) );
INVx2_ASAP7_75t_L g1500 ( .A(n_1432), .Y(n_1500) );
NAND2x1_ASAP7_75t_L g1501 ( .A(n_1398), .B(n_1273), .Y(n_1501) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_1430), .B(n_1378), .Y(n_1502) );
AND2x4_ASAP7_75t_L g1503 ( .A(n_1460), .B(n_1333), .Y(n_1503) );
AND2x4_ASAP7_75t_L g1504 ( .A(n_1444), .B(n_1404), .Y(n_1504) );
NOR3xp33_ASAP7_75t_SL g1505 ( .A(n_1400), .B(n_1377), .C(n_1358), .Y(n_1505) );
NOR3xp33_ASAP7_75t_SL g1506 ( .A(n_1410), .B(n_1356), .C(n_1364), .Y(n_1506) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1449), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1451), .B(n_1361), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1437), .B(n_1297), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1437), .B(n_1370), .Y(n_1510) );
INVxp67_ASAP7_75t_L g1511 ( .A(n_1412), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1451), .B(n_1366), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1436), .B(n_1369), .Y(n_1513) );
NAND3xp33_ASAP7_75t_L g1514 ( .A(n_1425), .B(n_1366), .C(n_1333), .Y(n_1514) );
NAND2x1_ASAP7_75t_L g1515 ( .A(n_1398), .B(n_1333), .Y(n_1515) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1438), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1403), .B(n_1366), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1406), .B(n_1354), .Y(n_1518) );
INVx1_ASAP7_75t_SL g1519 ( .A(n_1458), .Y(n_1519) );
NAND3xp33_ASAP7_75t_SL g1520 ( .A(n_1457), .B(n_1354), .C(n_1333), .Y(n_1520) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_1429), .B(n_1462), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_1429), .B(n_1476), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1523 ( .A(n_1421), .B(n_1423), .Y(n_1523) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1454), .Y(n_1524) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1456), .Y(n_1525) );
AND2x4_ASAP7_75t_L g1526 ( .A(n_1444), .B(n_1404), .Y(n_1526) );
AND2x4_ASAP7_75t_SL g1527 ( .A(n_1398), .B(n_1401), .Y(n_1527) );
OR2x2_ASAP7_75t_L g1528 ( .A(n_1419), .B(n_1439), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1476), .B(n_1414), .Y(n_1529) );
OR2x2_ASAP7_75t_L g1530 ( .A(n_1439), .B(n_1477), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1414), .B(n_1426), .Y(n_1531) );
NOR2x1p5_ASAP7_75t_L g1532 ( .A(n_1409), .B(n_1414), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1407), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_1436), .B(n_1441), .Y(n_1534) );
BUFx3_ASAP7_75t_L g1535 ( .A(n_1401), .Y(n_1535) );
NOR2xp33_ASAP7_75t_L g1536 ( .A(n_1459), .B(n_1473), .Y(n_1536) );
INVx2_ASAP7_75t_L g1537 ( .A(n_1443), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1441), .B(n_1405), .Y(n_1538) );
OR2x2_ASAP7_75t_L g1539 ( .A(n_1465), .B(n_1405), .Y(n_1539) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1407), .Y(n_1540) );
INVx2_ASAP7_75t_L g1541 ( .A(n_1443), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1542 ( .A(n_1426), .B(n_1433), .Y(n_1542) );
INVxp33_ASAP7_75t_L g1543 ( .A(n_1450), .Y(n_1543) );
INVx2_ASAP7_75t_L g1544 ( .A(n_1399), .Y(n_1544) );
NOR2xp33_ASAP7_75t_L g1545 ( .A(n_1459), .B(n_1409), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1455), .B(n_1466), .Y(n_1546) );
NOR2xp33_ASAP7_75t_L g1547 ( .A(n_1409), .B(n_1468), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1464), .B(n_1470), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1464), .B(n_1470), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1411), .B(n_1416), .Y(n_1550) );
INVx1_ASAP7_75t_SL g1551 ( .A(n_1446), .Y(n_1551) );
NAND4xp25_ASAP7_75t_L g1552 ( .A(n_1475), .B(n_1440), .C(n_1420), .D(n_1474), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1411), .B(n_1413), .Y(n_1553) );
AND2x4_ASAP7_75t_L g1554 ( .A(n_1418), .B(n_1474), .Y(n_1554) );
BUFx2_ASAP7_75t_L g1555 ( .A(n_1446), .Y(n_1555) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1537), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_1509), .B(n_1463), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1509), .B(n_1463), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1486), .B(n_1461), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1490), .B(n_1461), .Y(n_1560) );
OAI211xp5_ASAP7_75t_L g1561 ( .A1(n_1547), .A2(n_1431), .B(n_1485), .C(n_1484), .Y(n_1561) );
AND2x4_ASAP7_75t_L g1562 ( .A(n_1503), .B(n_1472), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1494), .Y(n_1563) );
OR2x2_ASAP7_75t_L g1564 ( .A(n_1528), .B(n_1434), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1507), .B(n_1434), .Y(n_1565) );
OAI31xp33_ASAP7_75t_L g1566 ( .A1(n_1532), .A2(n_1452), .A3(n_1435), .B(n_1418), .Y(n_1566) );
INVx2_ASAP7_75t_L g1567 ( .A(n_1537), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1548), .B(n_1472), .Y(n_1568) );
INVx2_ASAP7_75t_L g1569 ( .A(n_1541), .Y(n_1569) );
OR2x2_ASAP7_75t_L g1570 ( .A(n_1534), .B(n_1442), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1548), .B(n_1471), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1549), .B(n_1471), .Y(n_1572) );
AND2x4_ASAP7_75t_L g1573 ( .A(n_1503), .B(n_1482), .Y(n_1573) );
OR2x2_ASAP7_75t_L g1574 ( .A(n_1534), .B(n_1442), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1508), .B(n_1468), .Y(n_1575) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1494), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1549), .B(n_1415), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1524), .B(n_1417), .Y(n_1578) );
INVx1_ASAP7_75t_SL g1579 ( .A(n_1535), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1513), .B(n_1415), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1581 ( .A(n_1525), .B(n_1408), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1513), .B(n_1538), .Y(n_1582) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_1539), .B(n_1413), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1538), .B(n_1415), .Y(n_1584) );
OR2x2_ASAP7_75t_L g1585 ( .A(n_1502), .B(n_1416), .Y(n_1585) );
NAND2xp5_ASAP7_75t_SL g1586 ( .A(n_1547), .B(n_1418), .Y(n_1586) );
HB1xp67_ASAP7_75t_L g1587 ( .A(n_1511), .Y(n_1587) );
INVx3_ASAP7_75t_L g1588 ( .A(n_1503), .Y(n_1588) );
OAI31xp33_ASAP7_75t_L g1589 ( .A1(n_1552), .A2(n_1452), .A3(n_1435), .B(n_1467), .Y(n_1589) );
INVx2_ASAP7_75t_L g1590 ( .A(n_1544), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1504), .B(n_1482), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1504), .B(n_1478), .Y(n_1592) );
HB1xp67_ASAP7_75t_L g1593 ( .A(n_1511), .Y(n_1593) );
OR2x2_ASAP7_75t_L g1594 ( .A(n_1530), .B(n_1422), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1533), .B(n_1422), .Y(n_1595) );
NAND2xp5_ASAP7_75t_L g1596 ( .A(n_1540), .B(n_1428), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1504), .B(n_1478), .Y(n_1597) );
NOR2xp33_ASAP7_75t_L g1598 ( .A(n_1519), .B(n_1481), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1526), .B(n_1483), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1526), .B(n_1483), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1526), .B(n_1480), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1602 ( .A(n_1500), .B(n_1427), .Y(n_1602) );
OAI321xp33_ASAP7_75t_L g1603 ( .A1(n_1561), .A2(n_1542), .A3(n_1514), .B1(n_1495), .B2(n_1512), .C(n_1523), .Y(n_1603) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1570), .Y(n_1604) );
NAND4xp25_ASAP7_75t_L g1605 ( .A(n_1589), .B(n_1495), .C(n_1536), .D(n_1545), .Y(n_1605) );
OAI221xp5_ASAP7_75t_L g1606 ( .A1(n_1589), .A2(n_1536), .B1(n_1545), .B2(n_1506), .C(n_1505), .Y(n_1606) );
INVx2_ASAP7_75t_L g1607 ( .A(n_1556), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1582), .B(n_1522), .Y(n_1608) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1570), .Y(n_1609) );
OAI22xp5_ASAP7_75t_L g1610 ( .A1(n_1561), .A2(n_1535), .B1(n_1543), .B2(n_1527), .Y(n_1610) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1574), .Y(n_1611) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1574), .Y(n_1612) );
A2O1A1Ixp33_ASAP7_75t_L g1613 ( .A1(n_1566), .A2(n_1527), .B(n_1543), .C(n_1506), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1582), .B(n_1496), .Y(n_1614) );
AO32x1_ASAP7_75t_L g1615 ( .A1(n_1580), .A2(n_1493), .A3(n_1518), .B1(n_1529), .B2(n_1516), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1616 ( .A(n_1582), .B(n_1521), .Y(n_1616) );
AND2x4_ASAP7_75t_L g1617 ( .A(n_1588), .B(n_1496), .Y(n_1617) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1587), .Y(n_1618) );
AOI22xp5_ASAP7_75t_L g1619 ( .A1(n_1575), .A2(n_1496), .B1(n_1531), .B2(n_1554), .Y(n_1619) );
A2O1A1Ixp33_ASAP7_75t_L g1620 ( .A1(n_1566), .A2(n_1586), .B(n_1579), .C(n_1575), .Y(n_1620) );
AOI21xp5_ASAP7_75t_L g1621 ( .A1(n_1579), .A2(n_1499), .B(n_1520), .Y(n_1621) );
NAND4xp25_ASAP7_75t_SL g1622 ( .A(n_1571), .B(n_1488), .C(n_1487), .D(n_1489), .Y(n_1622) );
OAI21xp33_ASAP7_75t_SL g1623 ( .A1(n_1598), .A2(n_1491), .B(n_1546), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1571), .B(n_1554), .Y(n_1624) );
OAI21xp5_ASAP7_75t_SL g1625 ( .A1(n_1593), .A2(n_1554), .B(n_1492), .Y(n_1625) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1594), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1571), .B(n_1517), .Y(n_1627) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1594), .Y(n_1628) );
OAI22xp5_ASAP7_75t_L g1629 ( .A1(n_1583), .A2(n_1497), .B1(n_1498), .B2(n_1501), .Y(n_1629) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1583), .Y(n_1630) );
NOR2x1_ASAP7_75t_L g1631 ( .A(n_1564), .B(n_1515), .Y(n_1631) );
INVx1_ASAP7_75t_SL g1632 ( .A(n_1591), .Y(n_1632) );
INVxp67_ASAP7_75t_L g1633 ( .A(n_1559), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1572), .B(n_1510), .Y(n_1634) );
A2O1A1Ixp33_ASAP7_75t_L g1635 ( .A1(n_1577), .A2(n_1505), .B(n_1467), .C(n_1555), .Y(n_1635) );
OAI21xp5_ASAP7_75t_L g1636 ( .A1(n_1578), .A2(n_1469), .B(n_1551), .Y(n_1636) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1564), .Y(n_1637) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1578), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1572), .B(n_1510), .Y(n_1639) );
INVx2_ASAP7_75t_L g1640 ( .A(n_1607), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1623), .B(n_1584), .Y(n_1641) );
OAI21xp5_ASAP7_75t_L g1642 ( .A1(n_1620), .A2(n_1584), .B(n_1581), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1618), .Y(n_1643) );
AOI31xp33_ASAP7_75t_SL g1644 ( .A1(n_1621), .A2(n_1557), .A3(n_1558), .B(n_1585), .Y(n_1644) );
HB1xp67_ASAP7_75t_L g1645 ( .A(n_1632), .Y(n_1645) );
OAI21xp33_ASAP7_75t_L g1646 ( .A1(n_1625), .A2(n_1584), .B(n_1558), .Y(n_1646) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1638), .Y(n_1647) );
INVxp67_ASAP7_75t_L g1648 ( .A(n_1626), .Y(n_1648) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1630), .Y(n_1649) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1628), .Y(n_1650) );
OAI221xp5_ASAP7_75t_SL g1651 ( .A1(n_1625), .A2(n_1577), .B1(n_1580), .B2(n_1585), .C(n_1557), .Y(n_1651) );
INVx2_ASAP7_75t_L g1652 ( .A(n_1632), .Y(n_1652) );
OAI21xp5_ASAP7_75t_L g1653 ( .A1(n_1603), .A2(n_1581), .B(n_1467), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1633), .B(n_1580), .Y(n_1654) );
INVx2_ASAP7_75t_L g1655 ( .A(n_1631), .Y(n_1655) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1637), .Y(n_1656) );
OR2x2_ASAP7_75t_L g1657 ( .A(n_1604), .B(n_1577), .Y(n_1657) );
NOR2x1_ASAP7_75t_L g1658 ( .A(n_1613), .B(n_1553), .Y(n_1658) );
AO22x2_ASAP7_75t_L g1659 ( .A1(n_1610), .A2(n_1559), .B1(n_1560), .B2(n_1565), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1608), .B(n_1572), .Y(n_1660) );
INVxp67_ASAP7_75t_SL g1661 ( .A(n_1636), .Y(n_1661) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1609), .Y(n_1662) );
AND2x4_ASAP7_75t_L g1663 ( .A(n_1617), .B(n_1588), .Y(n_1663) );
NOR2xp33_ASAP7_75t_L g1664 ( .A(n_1605), .B(n_1560), .Y(n_1664) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1611), .Y(n_1665) );
CKINVDCx5p33_ASAP7_75t_R g1666 ( .A(n_1661), .Y(n_1666) );
O2A1O1Ixp33_ASAP7_75t_L g1667 ( .A1(n_1644), .A2(n_1606), .B(n_1605), .C(n_1635), .Y(n_1667) );
AOI221xp5_ASAP7_75t_L g1668 ( .A1(n_1664), .A2(n_1622), .B1(n_1629), .B2(n_1612), .C(n_1627), .Y(n_1668) );
AOI21xp33_ASAP7_75t_L g1669 ( .A1(n_1664), .A2(n_1565), .B(n_1619), .Y(n_1669) );
AOI21xp33_ASAP7_75t_L g1670 ( .A1(n_1653), .A2(n_1595), .B(n_1596), .Y(n_1670) );
AOI22xp5_ASAP7_75t_L g1671 ( .A1(n_1658), .A2(n_1617), .B1(n_1614), .B2(n_1592), .Y(n_1671) );
INVx1_ASAP7_75t_SL g1672 ( .A(n_1645), .Y(n_1672) );
OAI22xp5_ASAP7_75t_L g1673 ( .A1(n_1641), .A2(n_1616), .B1(n_1639), .B2(n_1634), .Y(n_1673) );
OAI21x1_ASAP7_75t_SL g1674 ( .A1(n_1642), .A2(n_1615), .B(n_1595), .Y(n_1674) );
AOI21xp5_ASAP7_75t_SL g1675 ( .A1(n_1646), .A2(n_1615), .B(n_1596), .Y(n_1675) );
AOI22x1_ASAP7_75t_L g1676 ( .A1(n_1659), .A2(n_1624), .B1(n_1615), .B2(n_1588), .Y(n_1676) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1647), .Y(n_1677) );
AOI211x1_ASAP7_75t_SL g1678 ( .A1(n_1655), .A2(n_1602), .B(n_1556), .C(n_1567), .Y(n_1678) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1647), .Y(n_1679) );
OAI221xp5_ASAP7_75t_L g1680 ( .A1(n_1651), .A2(n_1588), .B1(n_1601), .B2(n_1600), .C(n_1599), .Y(n_1680) );
AOI21xp5_ASAP7_75t_L g1681 ( .A1(n_1659), .A2(n_1602), .B(n_1601), .Y(n_1681) );
OAI21xp33_ASAP7_75t_L g1682 ( .A1(n_1659), .A2(n_1601), .B(n_1600), .Y(n_1682) );
AOI221x1_ASAP7_75t_L g1683 ( .A1(n_1659), .A2(n_1480), .B1(n_1479), .B2(n_1563), .C(n_1576), .Y(n_1683) );
NOR3xp33_ASAP7_75t_L g1684 ( .A(n_1667), .B(n_1655), .C(n_1643), .Y(n_1684) );
AOI211xp5_ASAP7_75t_L g1685 ( .A1(n_1675), .A2(n_1648), .B(n_1663), .C(n_1652), .Y(n_1685) );
OAI211xp5_ASAP7_75t_L g1686 ( .A1(n_1666), .A2(n_1654), .B(n_1652), .C(n_1650), .Y(n_1686) );
AOI32xp33_ASAP7_75t_L g1687 ( .A1(n_1668), .A2(n_1663), .A3(n_1656), .B1(n_1649), .B2(n_1665), .Y(n_1687) );
O2A1O1Ixp33_ASAP7_75t_L g1688 ( .A1(n_1674), .A2(n_1662), .B(n_1657), .C(n_1660), .Y(n_1688) );
AOI221xp5_ASAP7_75t_L g1689 ( .A1(n_1682), .A2(n_1663), .B1(n_1657), .B2(n_1640), .C(n_1600), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1673), .B(n_1640), .Y(n_1690) );
OAI21xp5_ASAP7_75t_L g1691 ( .A1(n_1666), .A2(n_1599), .B(n_1597), .Y(n_1691) );
OAI211xp5_ASAP7_75t_L g1692 ( .A1(n_1675), .A2(n_1599), .B(n_1592), .C(n_1597), .Y(n_1692) );
BUFx2_ASAP7_75t_L g1693 ( .A(n_1672), .Y(n_1693) );
AOI221xp5_ASAP7_75t_L g1694 ( .A1(n_1670), .A2(n_1597), .B1(n_1592), .B2(n_1568), .C(n_1591), .Y(n_1694) );
OAI21xp33_ASAP7_75t_L g1695 ( .A1(n_1671), .A2(n_1591), .B(n_1568), .Y(n_1695) );
NAND3xp33_ASAP7_75t_SL g1696 ( .A(n_1678), .B(n_1568), .C(n_1550), .Y(n_1696) );
HB1xp67_ASAP7_75t_L g1697 ( .A(n_1693), .Y(n_1697) );
NOR4xp75_ASAP7_75t_SL g1698 ( .A(n_1690), .B(n_1676), .C(n_1669), .D(n_1683), .Y(n_1698) );
NAND2xp5_ASAP7_75t_L g1699 ( .A(n_1684), .B(n_1679), .Y(n_1699) );
NOR2x1_ASAP7_75t_L g1700 ( .A(n_1692), .B(n_1681), .Y(n_1700) );
INVx1_ASAP7_75t_SL g1701 ( .A(n_1691), .Y(n_1701) );
NAND2x1p5_ASAP7_75t_L g1702 ( .A(n_1685), .B(n_1453), .Y(n_1702) );
XNOR2x1_ASAP7_75t_L g1703 ( .A(n_1687), .B(n_1677), .Y(n_1703) );
INVx2_ASAP7_75t_L g1704 ( .A(n_1696), .Y(n_1704) );
OR3x1_ASAP7_75t_L g1705 ( .A(n_1688), .B(n_1680), .C(n_1576), .Y(n_1705) );
INVx2_ASAP7_75t_SL g1706 ( .A(n_1697), .Y(n_1706) );
OAI222xp33_ASAP7_75t_L g1707 ( .A1(n_1701), .A2(n_1686), .B1(n_1689), .B2(n_1695), .C1(n_1694), .C2(n_1562), .Y(n_1707) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1699), .Y(n_1708) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1699), .Y(n_1709) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1704), .Y(n_1710) );
INVx3_ASAP7_75t_L g1711 ( .A(n_1702), .Y(n_1711) );
OAI22xp5_ASAP7_75t_L g1712 ( .A1(n_1711), .A2(n_1705), .B1(n_1701), .B2(n_1703), .Y(n_1712) );
OR2x2_ASAP7_75t_L g1713 ( .A(n_1706), .B(n_1698), .Y(n_1713) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1706), .B(n_1700), .Y(n_1714) );
INVx1_ASAP7_75t_SL g1715 ( .A(n_1710), .Y(n_1715) );
HB1xp67_ASAP7_75t_L g1716 ( .A(n_1715), .Y(n_1716) );
OAI22xp5_ASAP7_75t_L g1717 ( .A1(n_1712), .A2(n_1711), .B1(n_1709), .B2(n_1708), .Y(n_1717) );
XNOR2xp5_ASAP7_75t_L g1718 ( .A(n_1713), .B(n_1711), .Y(n_1718) );
AOI22x1_ASAP7_75t_L g1719 ( .A1(n_1718), .A2(n_1714), .B1(n_1707), .B2(n_1424), .Y(n_1719) );
AOI22xp33_ASAP7_75t_SL g1720 ( .A1(n_1717), .A2(n_1453), .B1(n_1573), .B2(n_1562), .Y(n_1720) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1716), .Y(n_1721) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1721), .Y(n_1722) );
AOI22x1_ASAP7_75t_L g1723 ( .A1(n_1722), .A2(n_1719), .B1(n_1720), .B2(n_1573), .Y(n_1723) );
AOI21xp5_ASAP7_75t_L g1724 ( .A1(n_1723), .A2(n_1590), .B(n_1569), .Y(n_1724) );
endmodule