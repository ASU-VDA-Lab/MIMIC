module fake_jpeg_29372_n_544 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_544);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_544;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g137 ( 
.A(n_55),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_59),
.Y(n_153)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_7),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_66),
.Y(n_113)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_7),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_7),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_91),
.Y(n_121)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_26),
.Y(n_70)
);

NAND2x1_ASAP7_75t_SL g133 ( 
.A(n_70),
.B(n_51),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_35),
.B(n_6),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_95),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_105),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_51),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_104),
.B(n_106),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_28),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_108),
.Y(n_142)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_110),
.Y(n_154)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_112),
.B(n_96),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_52),
.B1(n_44),
.B2(n_37),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_115),
.A2(n_128),
.B1(n_136),
.B2(n_45),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_48),
.B1(n_53),
.B2(n_52),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g217 ( 
.A1(n_117),
.A2(n_156),
.B1(n_97),
.B2(n_36),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_48),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_120),
.B(n_145),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_87),
.B(n_52),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_103),
.C(n_71),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_101),
.B1(n_56),
.B2(n_82),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_78),
.A2(n_44),
.B1(n_37),
.B2(n_45),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_64),
.B(n_22),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_141),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_60),
.B(n_22),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_64),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_150),
.B(n_163),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_67),
.B(n_54),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_151),
.B(n_155),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_54),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_41),
.B1(n_47),
.B2(n_43),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_41),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_58),
.B(n_20),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_164),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_108),
.B(n_47),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_63),
.B(n_29),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_173),
.Y(n_183)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_178),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_29),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_192),
.Y(n_243)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_113),
.A2(n_57),
.B1(n_88),
.B2(n_75),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_182),
.B(n_186),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_184),
.A2(n_177),
.B1(n_138),
.B2(n_135),
.Y(n_235)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_185),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_121),
.B(n_100),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_187),
.B(n_191),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_134),
.A2(n_61),
.B1(n_83),
.B2(n_76),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_188),
.A2(n_195),
.B1(n_200),
.B2(n_202),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_113),
.B(n_23),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_132),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_197),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_147),
.B1(n_152),
.B2(n_153),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_132),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_142),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_211),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_152),
.A2(n_72),
.B1(n_65),
.B2(n_45),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_126),
.B(n_43),
.C(n_34),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_201),
.B(n_222),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_37),
.B1(n_45),
.B2(n_23),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_37),
.B1(n_34),
.B2(n_51),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_231),
.B1(n_114),
.B2(n_174),
.Y(n_241)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_205),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_126),
.B(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_220),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_125),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_213),
.Y(n_259)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_216),
.Y(n_249)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_116),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_217),
.A2(n_157),
.B1(n_166),
.B2(n_130),
.Y(n_258)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_133),
.B(n_110),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_219),
.A2(n_227),
.B(n_14),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_118),
.B(n_9),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_36),
.B1(n_9),
.B2(n_15),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_115),
.B1(n_168),
.B2(n_166),
.Y(n_240)
);

AO22x2_ASAP7_75t_L g222 ( 
.A1(n_158),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_226),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_12),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_117),
.B(n_12),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_158),
.A2(n_6),
.B(n_15),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_230),
.Y(n_268)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_183),
.B(n_154),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_137),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_235),
.B(n_179),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_198),
.A2(n_128),
.B1(n_165),
.B2(n_136),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_239),
.B(n_203),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_245),
.B1(n_266),
.B2(n_261),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_241),
.A2(n_242),
.B1(n_256),
.B2(n_228),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_182),
.A2(n_198),
.B1(n_135),
.B2(n_114),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_161),
.B1(n_168),
.B2(n_130),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_210),
.B(n_219),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_218),
.A2(n_165),
.B1(n_111),
.B2(n_143),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_180),
.B(n_160),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_271),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_267),
.B1(n_191),
.B2(n_224),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_217),
.A2(n_127),
.B1(n_129),
.B2(n_143),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_187),
.A2(n_129),
.B1(n_111),
.B2(n_167),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_137),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_272),
.A2(n_273),
.B(n_279),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_237),
.A2(n_189),
.B1(n_213),
.B2(n_178),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_278),
.B1(n_280),
.B2(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_217),
.B1(n_222),
.B2(n_227),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_276),
.A2(n_282),
.B1(n_283),
.B2(n_300),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_277),
.B(n_271),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_258),
.B1(n_263),
.B2(n_248),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_239),
.A2(n_193),
.B1(n_223),
.B2(n_209),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_187),
.B1(n_192),
.B2(n_214),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_219),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_292),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_222),
.B1(n_212),
.B2(n_190),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_249),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_247),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_207),
.C(n_201),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_288),
.C(n_290),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_186),
.B(n_208),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_293),
.B(n_297),
.Y(n_324)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_229),
.C(n_215),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_222),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_291),
.B(n_233),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_216),
.C(n_205),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_263),
.B(n_185),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_296),
.Y(n_316)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_230),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_167),
.B(n_226),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_234),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_254),
.B(n_181),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_267),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_235),
.A2(n_179),
.B1(n_137),
.B2(n_55),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_257),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_301)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_304),
.A2(n_268),
.B(n_261),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_310),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_290),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_314),
.B(n_333),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_317),
.B(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_233),
.B(n_268),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_320),
.A2(n_261),
.B(n_265),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_274),
.A2(n_240),
.B1(n_243),
.B2(n_232),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_321),
.A2(n_330),
.B1(n_283),
.B2(n_276),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_247),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_323),
.Y(n_362)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_243),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_291),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_328),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_329),
.A2(n_297),
.B(n_303),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_282),
.A2(n_259),
.B1(n_238),
.B2(n_246),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_253),
.Y(n_332)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_332),
.Y(n_345)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_281),
.B(n_259),
.CI(n_253),
.CON(n_333),
.SN(n_333)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_331),
.A2(n_304),
.B1(n_293),
.B2(n_278),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_335),
.A2(n_342),
.B1(n_352),
.B2(n_320),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_336),
.B(n_332),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_338),
.A2(n_346),
.B1(n_350),
.B2(n_351),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_328),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_339),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_341),
.B(n_358),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_331),
.A2(n_293),
.B1(n_304),
.B2(n_294),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_296),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_327),
.C(n_334),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_321),
.A2(n_293),
.B1(n_272),
.B2(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_288),
.B1(n_292),
.B2(n_286),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_312),
.A2(n_285),
.B1(n_277),
.B2(n_280),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_301),
.B1(n_281),
.B2(n_302),
.Y(n_352)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_265),
.Y(n_356)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_312),
.A2(n_302),
.B1(n_238),
.B2(n_246),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_364),
.B1(n_313),
.B2(n_310),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_360),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_361),
.A2(n_309),
.B(n_269),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_330),
.A2(n_238),
.B1(n_244),
.B2(n_236),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_370),
.C(n_371),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_355),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_369),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_327),
.C(n_334),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_334),
.C(n_307),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_362),
.B(n_323),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_372),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_307),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_379),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_333),
.C(n_316),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_377),
.C(n_347),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_333),
.C(n_316),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_362),
.B(n_326),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_378),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_333),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_381),
.A2(n_389),
.B1(n_342),
.B2(n_358),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_340),
.B(n_325),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_382),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_335),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_393),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_384),
.B(n_319),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_318),
.Y(n_386)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_387),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_324),
.B1(n_309),
.B2(n_329),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_337),
.Y(n_391)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_391),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_392),
.A2(n_364),
.B1(n_343),
.B2(n_355),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_320),
.Y(n_393)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

XOR2x2_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_346),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_398),
.B(n_405),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_410),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_403),
.A2(n_365),
.B1(n_395),
.B2(n_389),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_345),
.B1(n_360),
.B2(n_359),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_407),
.Y(n_426)
);

XOR2x2_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_387),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_345),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_357),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_418),
.C(n_420),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_386),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_413),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_343),
.Y(n_414)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_414),
.Y(n_430)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_375),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_337),
.C(n_348),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_419),
.A2(n_425),
.B1(n_381),
.B2(n_415),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_319),
.C(n_306),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_394),
.Y(n_422)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_422),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_251),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_384),
.C(n_394),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_365),
.A2(n_313),
.B1(n_305),
.B2(n_353),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_428),
.A2(n_443),
.B1(n_447),
.B2(n_407),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_432),
.B(n_402),
.Y(n_454)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_397),
.Y(n_433)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_433),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_448),
.Y(n_456)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_414),
.Y(n_436)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_436),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_376),
.C(n_385),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_439),
.C(n_442),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_399),
.B(n_412),
.C(n_424),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_413),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_440),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_366),
.Y(n_441)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_379),
.C(n_366),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_423),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_428),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_420),
.A2(n_390),
.B(n_367),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_446),
.A2(n_419),
.B(n_401),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_425),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_396),
.B(n_380),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_468),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_SL g451 ( 
.A(n_446),
.B(n_417),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_451),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_442),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_457),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_438),
.B(n_406),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_461),
.Y(n_470)
);

FAx1_ASAP7_75t_SL g459 ( 
.A(n_438),
.B(n_406),
.CI(n_405),
.CON(n_459),
.SN(n_459)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_465),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_400),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_463),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_429),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_398),
.C(n_410),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_467),
.B(n_469),
.C(n_452),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_427),
.A2(n_411),
.B(n_400),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_408),
.C(n_305),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_471),
.B(n_452),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_472),
.B(n_478),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g476 ( 
.A(n_463),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_479),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_437),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_453),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_448),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_481),
.B(n_484),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_464),
.A2(n_427),
.B1(n_440),
.B2(n_444),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_482),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g483 ( 
.A(n_450),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_483),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_436),
.B1(n_430),
.B2(n_433),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_431),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_468),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_461),
.A2(n_430),
.B1(n_431),
.B2(n_449),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_459),
.C(n_408),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_460),
.A2(n_426),
.B1(n_434),
.B2(n_467),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_487),
.A2(n_456),
.B1(n_468),
.B2(n_462),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_488),
.B(n_501),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_494),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_454),
.C(n_458),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_475),
.C(n_482),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_426),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_497),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_470),
.B(n_459),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_500),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_449),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_416),
.B1(n_353),
.B2(n_308),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_480),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_502),
.B(n_236),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_251),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_270),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_496),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_516),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_509),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_475),
.C(n_483),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_507),
.C(n_503),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_490),
.C(n_495),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_492),
.A2(n_308),
.B(n_234),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_508),
.A2(n_513),
.B(n_6),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g512 ( 
.A(n_497),
.B(n_236),
.CI(n_295),
.CON(n_512),
.SN(n_512)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_512),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_492),
.A2(n_234),
.B(n_269),
.Y(n_513)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_498),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_515),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_523),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_SL g520 ( 
.A1(n_504),
.A2(n_493),
.B1(n_270),
.B2(n_262),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_520),
.B(n_521),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_507),
.A2(n_262),
.B(n_260),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_505),
.A2(n_179),
.B(n_13),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_522),
.A2(n_508),
.B(n_506),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_527),
.C(n_512),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_511),
.A2(n_14),
.B(n_15),
.Y(n_527)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_528),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_524),
.A2(n_514),
.B(n_510),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_532),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_518),
.A2(n_510),
.B(n_516),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_533),
.A2(n_526),
.B(n_3),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_529),
.A2(n_520),
.B(n_519),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_537),
.Y(n_539)
);

OAI311xp33_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_530),
.A3(n_3),
.B1(n_5),
.C1(n_0),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_535),
.C(n_3),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_540),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_539),
.C(n_3),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_5),
.B(n_386),
.Y(n_543)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_543),
.Y(n_544)
);


endmodule