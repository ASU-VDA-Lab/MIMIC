module fake_jpeg_7027_n_214 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g21 ( 
.A(n_9),
.B(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_31),
.B(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_8),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_47),
.B(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_54),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_29),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_29),
.B(n_27),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_75),
.Y(n_96)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_59),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_14),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_67),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_15),
.B1(n_25),
.B2(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_65),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_107)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_26),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_73),
.Y(n_101)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_20),
.C(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_24),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_18),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_53),
.B1(n_56),
.B2(n_48),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_65),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_22),
.B1(n_20),
.B2(n_25),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_98),
.B1(n_107),
.B2(n_109),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_25),
.B1(n_15),
.B2(n_4),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_77),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_106),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_75),
.C(n_68),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_114),
.C(n_119),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_63),
.C(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_51),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_57),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_72),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_6),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_58),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_134),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_84),
.B(n_60),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_104),
.B(n_90),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_58),
.Y(n_132)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_153),
.B(n_154),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_134),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_89),
.C(n_106),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_126),
.C(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_155),
.B(n_133),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_89),
.B(n_100),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_101),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_87),
.B(n_60),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_150),
.B1(n_152),
.B2(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_145),
.B1(n_138),
.B2(n_141),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_127),
.B1(n_119),
.B2(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_165),
.B1(n_154),
.B2(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_169),
.Y(n_183)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_123),
.B1(n_112),
.B2(n_124),
.C(n_113),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_137),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_114),
.B1(n_121),
.B2(n_130),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_124),
.C(n_92),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.C(n_153),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_69),
.C(n_101),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_140),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_138),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_158),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_168),
.B1(n_166),
.B2(n_170),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_160),
.B(n_140),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_175),
.C(n_176),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_169),
.B(n_154),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_165),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_145),
.C(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_173),
.C(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_187),
.B(n_190),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_189),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_159),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_168),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_157),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_149),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_194),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_162),
.B1(n_159),
.B2(n_178),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_177),
.B(n_136),
.C(n_188),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_199),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_192),
.B(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_204),
.A3(n_193),
.B1(n_186),
.B2(n_136),
.C1(n_147),
.C2(n_143),
.Y(n_205)
);

OAI31xp33_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_195),
.A3(n_198),
.B(n_199),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_186),
.B(n_163),
.C(n_69),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_149),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_143),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_211),
.B(n_87),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_105),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);


endmodule