module fake_aes_4518_n_589 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_589);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_589;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_476;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_163;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_65), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_7), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_6), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_52), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_33), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_78), .Y(n_88) );
BUFx2_ASAP7_75t_SL g89 ( .A(n_53), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_36), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_56), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_59), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_9), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_66), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_3), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_32), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_5), .Y(n_99) );
NOR2xp33_ASAP7_75t_L g100 ( .A(n_15), .B(n_18), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_80), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_69), .Y(n_102) );
BUFx5_ASAP7_75t_L g103 ( .A(n_72), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_73), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_16), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_14), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_24), .B(n_4), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_9), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_4), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_22), .Y(n_112) );
INVxp33_ASAP7_75t_L g113 ( .A(n_25), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_64), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_46), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_70), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_1), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_91), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_112), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_84), .Y(n_122) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_97), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_93), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_93), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_87), .B(n_0), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_113), .B(n_1), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_105), .Y(n_130) );
INVx5_ASAP7_75t_L g131 ( .A(n_105), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_88), .B(n_2), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_106), .B(n_107), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_83), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_103), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_124), .B(n_98), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_141), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_126), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_124), .B(n_101), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_132), .A2(n_86), .B1(n_94), .B2(n_117), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_126), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_126), .B(n_109), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_125), .B(n_102), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_132), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_131), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_137), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_138), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_127), .B(n_108), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_125), .A2(n_108), .B(n_104), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_137), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_152), .B(n_121), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_173), .B(n_127), .Y(n_176) );
NOR3xp33_ASAP7_75t_SL g177 ( .A(n_150), .B(n_106), .C(n_107), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_152), .B(n_134), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_173), .B(n_120), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_157), .B(n_128), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_169), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
AOI22xp33_ASAP7_75t_SL g184 ( .A1(n_150), .A2(n_117), .B1(n_94), .B2(n_123), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_152), .B(n_92), .Y(n_185) );
OAI22x1_ASAP7_75t_SL g186 ( .A1(n_154), .A2(n_123), .B1(n_111), .B2(n_115), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_164), .Y(n_187) );
OAI221xp5_ASAP7_75t_L g188 ( .A1(n_145), .A2(n_128), .B1(n_140), .B2(n_144), .C(n_136), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_164), .B(n_140), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g191 ( .A1(n_152), .A2(n_133), .B1(n_122), .B2(n_118), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_151), .B(n_92), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_151), .B(n_96), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_164), .B(n_135), .Y(n_194) );
NOR3xp33_ASAP7_75t_SL g195 ( .A(n_145), .B(n_96), .C(n_100), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_164), .B(n_131), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_148), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_116), .B1(n_110), .B2(n_114), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
AND3x1_ASAP7_75t_SL g201 ( .A(n_169), .B(n_119), .C(n_3), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_164), .B(n_130), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_149), .B(n_130), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
NOR3xp33_ASAP7_75t_SL g206 ( .A(n_149), .B(n_89), .C(n_5), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_153), .B(n_89), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_172), .B(n_103), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_172), .B(n_2), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_156), .A2(n_130), .B(n_129), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_208), .B(n_146), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_199), .B(n_172), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_205), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_188), .A2(n_172), .B(n_160), .C(n_147), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_199), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_175), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_180), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_205), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_180), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_205), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_176), .B(n_146), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_198), .B(n_147), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
NOR2x1_ASAP7_75t_L g226 ( .A(n_210), .B(n_155), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_187), .B(n_155), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_197), .A2(n_160), .B(n_165), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_183), .Y(n_230) );
INVx4_ASAP7_75t_L g231 ( .A(n_183), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_209), .A2(n_166), .B1(n_165), .B2(n_138), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_183), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_200), .B(n_166), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_197), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_183), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_174), .B(n_156), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_189), .A2(n_156), .B(n_171), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_183), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_203), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_181), .B(n_103), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_210), .B(n_159), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_209), .A2(n_139), .B1(n_129), .B2(n_130), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_181), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_204), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_202), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_204), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_245), .A2(n_184), .B1(n_191), .B2(n_178), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_245), .Y(n_250) );
AOI21x1_ASAP7_75t_L g251 ( .A1(n_226), .A2(n_211), .B(n_171), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_217), .B(n_196), .Y(n_252) );
OAI22xp33_ASAP7_75t_L g253 ( .A1(n_243), .A2(n_179), .B1(n_194), .B2(n_207), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_243), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_243), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_212), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_217), .B(n_177), .Y(n_257) );
INVx6_ASAP7_75t_L g258 ( .A(n_231), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_230), .Y(n_259) );
AOI22xp33_ASAP7_75t_SL g260 ( .A1(n_243), .A2(n_201), .B1(n_206), .B2(n_186), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_216), .A2(n_193), .B(n_192), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_216), .A2(n_182), .B(n_185), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_228), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_212), .Y(n_265) );
AOI21x1_ASAP7_75t_L g266 ( .A1(n_226), .A2(n_182), .B(n_158), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_230), .Y(n_267) );
OA21x2_ASAP7_75t_L g268 ( .A1(n_244), .A2(n_195), .B(n_103), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_229), .A2(n_204), .B(n_170), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_229), .A2(n_159), .B(n_167), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_219), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_217), .B(n_204), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_219), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_230), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_217), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_223), .B(n_214), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_221), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_249), .A2(n_241), .B1(n_223), .B2(n_214), .C(n_237), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_250), .B(n_214), .Y(n_280) );
BUFx10_ASAP7_75t_L g281 ( .A(n_254), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_269), .A2(n_238), .B(n_218), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_277), .A2(n_232), .B1(n_223), .B2(n_240), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_277), .B(n_241), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_269), .B(n_261), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_241), .B1(n_213), .B2(n_240), .C(n_224), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_256), .A2(n_238), .B(n_225), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g289 ( .A(n_260), .B(n_244), .C(n_232), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_254), .Y(n_290) );
AOI21x1_ASAP7_75t_L g291 ( .A1(n_266), .A2(n_248), .B(n_236), .Y(n_291) );
OAI221xp5_ASAP7_75t_L g292 ( .A1(n_260), .A2(n_235), .B1(n_218), .B2(n_225), .C(n_220), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_257), .A2(n_228), .B1(n_234), .B2(n_235), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_266), .A2(n_248), .B(n_236), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_256), .A2(n_278), .B(n_265), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_264), .A2(n_228), .B1(n_234), .B2(n_215), .Y(n_296) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_263), .B(n_231), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_264), .A2(n_228), .B1(n_234), .B2(n_215), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_253), .A2(n_234), .B1(n_247), .B2(n_227), .C(n_221), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_265), .B(n_221), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
OAI221xp5_ASAP7_75t_L g302 ( .A1(n_255), .A2(n_220), .B1(n_247), .B2(n_222), .C(n_215), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_255), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_300), .B(n_273), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_290), .B(n_273), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_300), .B(n_276), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_301), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_286), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_301), .B(n_276), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_297), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_303), .B(n_265), .Y(n_312) );
NOR2xp33_ASAP7_75t_SL g313 ( .A(n_283), .B(n_275), .Y(n_313) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_281), .B(n_271), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_303), .B(n_271), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_297), .B(n_271), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_297), .B(n_278), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_280), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_278), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_295), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_291), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_281), .B(n_275), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_294), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_283), .B(n_262), .Y(n_328) );
INVx5_ASAP7_75t_SL g329 ( .A(n_308), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_318), .A2(n_292), .B1(n_289), .B2(n_279), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g331 ( .A1(n_321), .A2(n_293), .B1(n_289), .B2(n_287), .C(n_296), .Y(n_331) );
AOI222xp33_ASAP7_75t_SL g332 ( .A1(n_307), .A2(n_6), .B1(n_8), .B2(n_10), .C1(n_11), .C2(n_12), .Y(n_332) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_311), .B(n_285), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_314), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_308), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_304), .B(n_285), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_314), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g340 ( .A1(n_313), .A2(n_298), .B1(n_299), .B2(n_268), .C(n_302), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_323), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_312), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_311), .B(n_282), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_313), .A2(n_288), .B(n_285), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_304), .B(n_285), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_306), .B(n_312), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_305), .B(n_262), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_323), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_306), .B(n_261), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g350 ( .A1(n_326), .A2(n_268), .B(n_139), .C(n_261), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_316), .B(n_259), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_324), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_305), .B(n_268), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_325), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_327), .A2(n_139), .B1(n_130), .B2(n_252), .C(n_227), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_316), .A2(n_268), .B1(n_252), .B2(n_258), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_326), .A2(n_268), .B1(n_252), .B2(n_258), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_315), .B(n_103), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_309), .B(n_274), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_336), .B(n_328), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_341), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_336), .B(n_328), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_345), .B(n_327), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_345), .B(n_324), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_337), .B(n_309), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_349), .B(n_324), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_342), .B(n_310), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_337), .B(n_322), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_348), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g372 ( .A1(n_330), .A2(n_315), .B(n_319), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_349), .B(n_317), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_348), .B(n_322), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_343), .B(n_320), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_346), .B(n_8), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_346), .B(n_317), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_347), .B(n_310), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_354), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_354), .B(n_355), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_355), .B(n_320), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_352), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_347), .B(n_319), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_331), .B(n_10), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_359), .B(n_320), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_359), .B(n_320), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
NOR3xp33_ASAP7_75t_SL g388 ( .A(n_340), .B(n_272), .C(n_270), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_343), .B(n_320), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_335), .B(n_320), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_334), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_339), .B(n_333), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_333), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_343), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_329), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_353), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_338), .B(n_314), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_353), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_329), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_350), .A2(n_274), .B(n_259), .Y(n_402) );
INVx6_ASAP7_75t_L g403 ( .A(n_338), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_329), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_338), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_360), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_329), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_380), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_376), .B(n_11), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_377), .B(n_351), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_400), .B(n_344), .Y(n_413) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_399), .B(n_351), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_377), .B(n_351), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_362), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_373), .B(n_358), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_399), .B(n_258), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_373), .B(n_357), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_366), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_383), .B(n_12), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_366), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_400), .B(n_356), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_406), .B(n_384), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_371), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_364), .B(n_103), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_399), .B(n_259), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_371), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_369), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_399), .B(n_139), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_364), .B(n_13), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_379), .B(n_139), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_379), .B(n_13), .Y(n_434) );
NOR3x1_ASAP7_75t_SL g435 ( .A(n_405), .B(n_332), .C(n_15), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_370), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_365), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_398), .B(n_14), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_370), .Y(n_439) );
OAI31xp33_ASAP7_75t_L g440 ( .A1(n_392), .A2(n_252), .A3(n_267), .B(n_274), .Y(n_440) );
XNOR2x2_ASAP7_75t_L g441 ( .A(n_372), .B(n_16), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_367), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_372), .A2(n_258), .B1(n_252), .B2(n_267), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_398), .B(n_17), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_367), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_361), .B(n_17), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_396), .B(n_267), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_398), .B(n_158), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_361), .B(n_158), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_383), .B(n_170), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_363), .B(n_258), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_363), .B(n_158), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_365), .B(n_158), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_374), .B(n_158), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_374), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_403), .B(n_19), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_368), .B(n_21), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_394), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_394), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_368), .B(n_168), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_396), .B(n_161), .C(n_162), .D(n_170), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_378), .B(n_168), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_427), .B(n_381), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_408), .Y(n_464) );
OAI322xp33_ASAP7_75t_L g465 ( .A1(n_441), .A2(n_422), .A3(n_425), .B1(n_442), .B2(n_445), .C1(n_410), .C2(n_413), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_436), .B(n_381), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_411), .A2(n_393), .B1(n_388), .B2(n_396), .C(n_395), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_415), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_414), .A2(n_403), .B1(n_378), .B2(n_397), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_421), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_439), .B(n_393), .Y(n_472) );
AOI332xp33_ASAP7_75t_L g473 ( .A1(n_446), .A2(n_387), .A3(n_382), .B1(n_389), .B2(n_385), .B3(n_386), .C1(n_395), .C2(n_394), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_423), .Y(n_474) );
AOI322xp5_ASAP7_75t_L g475 ( .A1(n_432), .A2(n_385), .A3(n_386), .B1(n_395), .B2(n_382), .C1(n_387), .C2(n_389), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
AOI21xp33_ASAP7_75t_L g477 ( .A1(n_434), .A2(n_375), .B(n_390), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_426), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_420), .A2(n_375), .B1(n_390), .B2(n_403), .Y(n_479) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_443), .A2(n_397), .B(n_404), .Y(n_480) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_419), .A2(n_403), .B1(n_397), .B2(n_404), .Y(n_481) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_419), .A2(n_403), .B1(n_397), .B2(n_404), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_440), .A2(n_401), .B(n_407), .C(n_402), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_431), .B(n_401), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_409), .B(n_391), .Y(n_486) );
AOI21xp33_ASAP7_75t_L g487 ( .A1(n_434), .A2(n_444), .B(n_438), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_455), .B(n_391), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_416), .B(n_390), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_412), .B(n_375), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_451), .B(n_390), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_433), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_418), .B(n_375), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_435), .B(n_402), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_419), .A2(n_401), .B1(n_407), .B2(n_231), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_431), .A2(n_407), .B1(n_231), .B2(n_220), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_449), .B(n_162), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_428), .A2(n_227), .B1(n_222), .B2(n_215), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_457), .A2(n_222), .B1(n_233), .B2(n_242), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_413), .B(n_239), .Y(n_502) );
NAND3xp33_ASAP7_75t_L g503 ( .A(n_449), .B(n_168), .C(n_162), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_438), .A2(n_251), .B(n_270), .Y(n_504) );
NAND2xp33_ASAP7_75t_SL g505 ( .A(n_444), .B(n_246), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_428), .A2(n_222), .B1(n_251), .B2(n_242), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_458), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_452), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_475), .A2(n_424), .B(n_453), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_468), .Y(n_512) );
OAI22xp33_ASAP7_75t_SL g513 ( .A1(n_469), .A2(n_456), .B1(n_424), .B2(n_450), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_509), .B(n_453), .Y(n_514) );
XOR2x2_ASAP7_75t_L g515 ( .A(n_496), .B(n_460), .Y(n_515) );
O2A1O1Ixp5_ASAP7_75t_L g516 ( .A1(n_465), .A2(n_469), .B(n_484), .C(n_481), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_507), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_482), .B(n_460), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_476), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_490), .B(n_447), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_495), .B(n_447), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_479), .A2(n_462), .B(n_454), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_486), .B(n_462), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_507), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_502), .Y(n_525) );
OAI322xp33_ASAP7_75t_L g526 ( .A1(n_472), .A2(n_454), .A3(n_448), .B1(n_168), .B2(n_461), .C1(n_248), .C2(n_236), .Y(n_526) );
OAI21xp33_ASAP7_75t_L g527 ( .A1(n_480), .A2(n_448), .B(n_168), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_467), .A2(n_242), .B1(n_233), .B2(n_168), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_464), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_473), .A2(n_477), .B(n_497), .C(n_505), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_510), .B(n_23), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_508), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_470), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_493), .B(n_26), .Y(n_534) );
AO22x2_ASAP7_75t_L g535 ( .A1(n_489), .A2(n_242), .B1(n_233), .B2(n_30), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_503), .B(n_246), .C(n_239), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_463), .A2(n_233), .B1(n_239), .B2(n_246), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_471), .B(n_28), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_506), .A2(n_246), .B1(n_239), .B2(n_167), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_474), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_478), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_487), .A2(n_29), .B(n_31), .C(n_34), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_512), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_533), .Y(n_544) );
AOI21xp33_ASAP7_75t_SL g545 ( .A1(n_513), .A2(n_500), .B(n_477), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_516), .A2(n_530), .B(n_527), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_519), .B(n_488), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_541), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_511), .B(n_492), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_519), .B(n_494), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_515), .A2(n_487), .B1(n_483), .B2(n_498), .C(n_506), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_518), .A2(n_466), .B1(n_485), .B2(n_491), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_540), .Y(n_553) );
OAI21xp5_ASAP7_75t_SL g554 ( .A1(n_528), .A2(n_501), .B(n_504), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_529), .A2(n_504), .B1(n_499), .B2(n_246), .C(n_239), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_517), .Y(n_556) );
NAND4xp75_ASAP7_75t_L g557 ( .A(n_534), .B(n_35), .C(n_37), .D(n_38), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_523), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_532), .Y(n_559) );
AOI221x1_ASAP7_75t_SL g560 ( .A1(n_522), .A2(n_39), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_514), .A2(n_246), .B1(n_239), .B2(n_167), .C(n_163), .Y(n_561) );
OAI211xp5_ASAP7_75t_L g562 ( .A1(n_546), .A2(n_542), .B(n_539), .C(n_525), .Y(n_562) );
NAND3xp33_ASAP7_75t_SL g563 ( .A(n_551), .B(n_536), .C(n_538), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_551), .A2(n_526), .B1(n_524), .B2(n_535), .C(n_538), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_550), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_552), .A2(n_535), .B1(n_521), .B2(n_520), .Y(n_566) );
AOI221xp5_ASAP7_75t_SL g567 ( .A1(n_545), .A2(n_526), .B1(n_531), .B2(n_537), .C(n_536), .Y(n_567) );
AOI222xp33_ASAP7_75t_L g568 ( .A1(n_549), .A2(n_43), .B1(n_44), .B2(n_45), .C1(n_47), .C2(n_48), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_558), .A2(n_163), .B1(n_159), .B2(n_167), .Y(n_569) );
OAI221xp5_ASAP7_75t_SL g570 ( .A1(n_554), .A2(n_553), .B1(n_547), .B2(n_555), .C(n_556), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_560), .A2(n_49), .B1(n_50), .B2(n_51), .C(n_55), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
OAI222xp33_ASAP7_75t_L g573 ( .A1(n_570), .A2(n_548), .B1(n_544), .B2(n_543), .C1(n_561), .C2(n_557), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_566), .B(n_58), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_562), .B(n_60), .Y(n_575) );
OAI211xp5_ASAP7_75t_SL g576 ( .A1(n_564), .A2(n_61), .B(n_62), .C(n_63), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_565), .B(n_67), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_572), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_578), .B(n_563), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_573), .B(n_571), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_575), .B(n_576), .C(n_574), .Y(n_581) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_579), .B(n_577), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_580), .B(n_568), .C(n_567), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_582), .Y(n_584) );
AO22x2_ASAP7_75t_L g585 ( .A1(n_583), .A2(n_581), .B1(n_569), .B2(n_76), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_585), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_586), .A2(n_584), .B1(n_163), .B2(n_159), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_587), .A2(n_163), .B1(n_74), .B2(n_77), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_588), .A2(n_68), .B1(n_79), .B2(n_81), .Y(n_589) );
endmodule