module real_aes_12263_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1699;
wire n_730;
wire n_1023;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1691;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AO221x1_ASAP7_75t_L g1465 ( .A1(n_0), .A2(n_122), .B1(n_1435), .B2(n_1466), .C(n_1468), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g1723 ( .A(n_1), .Y(n_1723) );
AOI22xp5_ASAP7_75t_L g1453 ( .A1(n_2), .A2(n_106), .B1(n_1435), .B2(n_1439), .Y(n_1453) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_3), .A2(n_280), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
INVx1_ASAP7_75t_L g1103 ( .A(n_3), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_4), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_5), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_6), .A2(n_85), .B1(n_1221), .B2(n_1223), .Y(n_1370) );
INVx1_ASAP7_75t_L g1409 ( .A(n_6), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_7), .A2(n_191), .B1(n_554), .B2(n_556), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_7), .A2(n_191), .B1(n_576), .B2(n_578), .Y(n_575) );
INVx1_ASAP7_75t_L g798 ( .A(n_8), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_9), .A2(n_183), .B1(n_391), .B2(n_986), .C(n_987), .Y(n_1046) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_9), .A2(n_276), .B1(n_474), .B2(n_995), .Y(n_1051) );
CKINVDCx5p33_ASAP7_75t_R g1071 ( .A(n_10), .Y(n_1071) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_11), .A2(n_27), .B1(n_708), .B2(n_901), .C(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g928 ( .A(n_11), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1657 ( .A1(n_12), .A2(n_135), .B1(n_875), .B2(n_1194), .Y(n_1657) );
INVx1_ASAP7_75t_L g1691 ( .A(n_12), .Y(n_1691) );
INVx1_ASAP7_75t_L g1469 ( .A(n_13), .Y(n_1469) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_14), .A2(n_260), .B1(n_421), .B2(n_422), .C(n_423), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_14), .A2(n_260), .B1(n_451), .B2(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g846 ( .A(n_15), .Y(n_846) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_15), .A2(n_254), .B1(n_865), .B2(n_867), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g1220 ( .A1(n_16), .A2(n_63), .B1(n_1221), .B2(n_1223), .Y(n_1220) );
OAI22xp33_ASAP7_75t_L g1229 ( .A1(n_16), .A2(n_167), .B1(n_326), .B2(n_613), .Y(n_1229) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_17), .Y(n_966) );
AO22x2_ASAP7_75t_L g509 ( .A1(n_18), .A2(n_510), .B1(n_615), .B2(n_616), .Y(n_509) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_18), .Y(n_615) );
XNOR2xp5_ASAP7_75t_L g934 ( .A(n_19), .B(n_935), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_20), .A2(n_309), .B1(n_587), .B2(n_795), .Y(n_1011) );
INVxp67_ASAP7_75t_SL g1037 ( .A(n_20), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_21), .A2(n_116), .B1(n_895), .B2(n_896), .Y(n_894) );
INVx1_ASAP7_75t_L g914 ( .A(n_21), .Y(n_914) );
INVx1_ASAP7_75t_L g1215 ( .A(n_22), .Y(n_1215) );
OAI222xp33_ASAP7_75t_L g1227 ( .A1(n_22), .A2(n_216), .B1(n_287), .B2(n_599), .C1(n_680), .C2(n_1228), .Y(n_1227) );
OAI222xp33_ASAP7_75t_L g1716 ( .A1(n_23), .A2(n_59), .B1(n_129), .B2(n_1168), .C1(n_1717), .C2(n_1718), .Y(n_1716) );
INVx1_ASAP7_75t_L g1733 ( .A(n_23), .Y(n_1733) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_24), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_25), .Y(n_1342) );
AOI22xp33_ASAP7_75t_SL g1179 ( .A1(n_26), .A2(n_114), .B1(n_861), .B2(n_1077), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_26), .A2(n_114), .B1(n_1043), .B2(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g926 ( .A(n_27), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_28), .A2(n_185), .B1(n_384), .B2(n_386), .C(n_391), .Y(n_383) );
INVx1_ASAP7_75t_L g480 ( .A(n_28), .Y(n_480) );
INVx1_ASAP7_75t_L g630 ( .A(n_29), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_29), .A2(n_143), .B1(n_690), .B2(n_692), .C(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g1165 ( .A(n_30), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_30), .A2(n_290), .B1(n_422), .B2(n_986), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1369 ( .A(n_31), .B(n_1219), .Y(n_1369) );
INVx1_ASAP7_75t_L g1407 ( .A(n_31), .Y(n_1407) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_32), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_33), .A2(n_139), .B1(n_1082), .B2(n_1196), .Y(n_1316) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_33), .A2(n_139), .B1(n_562), .B2(n_1333), .Y(n_1332) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_34), .A2(n_234), .B1(n_559), .B2(n_560), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_34), .A2(n_234), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g317 ( .A(n_35), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g1217 ( .A1(n_36), .A2(n_95), .B1(n_1218), .B2(n_1219), .Y(n_1217) );
AOI22xp33_ASAP7_75t_SL g1237 ( .A1(n_36), .A2(n_95), .B1(n_1184), .B2(n_1189), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_37), .A2(n_142), .B1(n_373), .B2(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g483 ( .A(n_37), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g1479 ( .A1(n_38), .A2(n_130), .B1(n_1435), .B2(n_1439), .Y(n_1479) );
INVx1_ASAP7_75t_L g1258 ( .A(n_39), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_39), .A2(n_205), .B1(n_986), .B2(n_1129), .Y(n_1296) );
INVx1_ASAP7_75t_L g1118 ( .A(n_40), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_40), .A2(n_256), .B1(n_564), .B2(n_567), .Y(n_1147) );
INVx1_ASAP7_75t_L g1231 ( .A(n_41), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_41), .A2(n_213), .B1(n_587), .B2(n_795), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_42), .A2(n_131), .B1(n_1094), .B2(n_1129), .Y(n_1292) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_42), .A2(n_131), .B1(n_865), .B2(n_1178), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_43), .A2(n_223), .B1(n_451), .B2(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1100 ( .A(n_43), .Y(n_1100) );
INVx1_ASAP7_75t_L g653 ( .A(n_44), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_44), .A2(n_111), .B1(n_585), .B2(n_712), .Y(n_711) );
AOI22x1_ASAP7_75t_SL g1207 ( .A1(n_45), .A2(n_1208), .B1(n_1248), .B2(n_1249), .Y(n_1207) );
INVx1_ASAP7_75t_L g1248 ( .A(n_45), .Y(n_1248) );
INVx1_ASAP7_75t_L g765 ( .A(n_46), .Y(n_765) );
INVx1_ASAP7_75t_L g886 ( .A(n_47), .Y(n_886) );
AO221x2_ASAP7_75t_L g1512 ( .A1(n_48), .A2(n_248), .B1(n_1466), .B2(n_1513), .C(n_1515), .Y(n_1512) );
INVx1_ASAP7_75t_L g1010 ( .A(n_49), .Y(n_1010) );
INVx1_ASAP7_75t_L g1173 ( .A(n_50), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_50), .A2(n_164), .B1(n_1182), .B2(n_1184), .Y(n_1181) );
INVx1_ASAP7_75t_L g984 ( .A(n_51), .Y(n_984) );
OAI22xp33_ASAP7_75t_L g994 ( .A1(n_51), .A2(n_113), .B1(n_474), .B2(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1138 ( .A(n_52), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_52), .A2(n_249), .B1(n_587), .B2(n_795), .Y(n_1158) );
INVx1_ASAP7_75t_L g1140 ( .A(n_53), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_53), .A2(n_274), .B1(n_585), .B2(n_1156), .Y(n_1157) );
INVx1_ASAP7_75t_L g1737 ( .A(n_54), .Y(n_1737) );
AOI22xp33_ASAP7_75t_SL g1752 ( .A1(n_54), .A2(n_94), .B1(n_1178), .B2(n_1303), .Y(n_1752) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_55), .A2(n_158), .B1(n_587), .B2(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g973 ( .A(n_55), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_56), .B(n_343), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g809 ( .A1(n_57), .A2(n_278), .B1(n_810), .B2(n_811), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_57), .A2(n_278), .B1(n_872), .B2(n_875), .Y(n_871) );
INVx1_ASAP7_75t_L g1125 ( .A(n_58), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_58), .A2(n_288), .B1(n_597), .B2(n_1134), .Y(n_1133) );
AOI22xp33_ASAP7_75t_SL g1740 ( .A1(n_59), .A2(n_268), .B1(n_1094), .B2(n_1191), .Y(n_1740) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_60), .A2(n_270), .B1(n_1435), .B2(n_1439), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_61), .A2(n_179), .B1(n_1182), .B2(n_1290), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_61), .A2(n_179), .B1(n_583), .B2(n_1299), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1447 ( .A1(n_62), .A2(n_292), .B1(n_1448), .B2(n_1451), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_63), .A2(n_127), .B1(n_554), .B2(n_1129), .Y(n_1238) );
INVxp33_ASAP7_75t_SL g740 ( .A(n_64), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_64), .A2(n_300), .B1(n_781), .B2(n_783), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_65), .Y(n_906) );
CKINVDCx5p33_ASAP7_75t_R g1064 ( .A(n_66), .Y(n_1064) );
AOI22xp33_ASAP7_75t_SL g1235 ( .A1(n_67), .A2(n_133), .B1(n_421), .B2(n_1129), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_67), .A2(n_133), .B1(n_585), .B2(n_1244), .Y(n_1243) );
AO22x1_ASAP7_75t_L g1474 ( .A1(n_68), .A2(n_238), .B1(n_1439), .B2(n_1475), .Y(n_1474) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_69), .A2(n_226), .B1(n_698), .B2(n_701), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g919 ( .A1(n_69), .A2(n_226), .B1(n_640), .B2(n_645), .C(n_648), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_70), .A2(n_302), .B1(n_870), .B2(n_1079), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1097 ( .A1(n_70), .A2(n_835), .B1(n_1038), .B2(n_1098), .C(n_1102), .Y(n_1097) );
INVx1_ASAP7_75t_L g1259 ( .A(n_71), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g1294 ( .A1(n_71), .A2(n_152), .B1(n_1182), .B2(n_1295), .Y(n_1294) );
AO22x1_ASAP7_75t_L g1476 ( .A1(n_72), .A2(n_237), .B1(n_1448), .B2(n_1451), .Y(n_1476) );
INVx1_ASAP7_75t_L g625 ( .A(n_73), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_73), .A2(n_210), .B1(n_582), .B2(n_696), .Y(n_695) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_74), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_75), .A2(n_230), .B1(n_583), .B2(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g604 ( .A(n_75), .Y(n_604) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_76), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g788 ( .A1(n_76), .A2(n_304), .B1(n_789), .B2(n_791), .C(n_792), .Y(n_788) );
INVx1_ASAP7_75t_L g531 ( .A(n_77), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_77), .A2(n_177), .B1(n_597), .B2(n_599), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_78), .Y(n_1005) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_79), .A2(n_99), .B1(n_640), .B2(n_645), .C(n_648), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_79), .A2(n_99), .B1(n_698), .B2(n_701), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g1668 ( .A1(n_80), .A2(n_301), .B1(n_1669), .B2(n_1671), .Y(n_1668) );
OAI221xp5_ASAP7_75t_L g1686 ( .A1(n_80), .A2(n_301), .B1(n_742), .B2(n_1687), .C(n_1688), .Y(n_1686) );
BUFx2_ASAP7_75t_L g346 ( .A(n_81), .Y(n_346) );
BUFx2_ASAP7_75t_L g361 ( .A(n_81), .Y(n_361) );
INVx1_ASAP7_75t_L g471 ( .A(n_81), .Y(n_471) );
OR2x2_ASAP7_75t_L g644 ( .A(n_81), .B(n_366), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g1236 ( .A1(n_82), .A2(n_221), .B1(n_559), .B2(n_1184), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_82), .A2(n_221), .B1(n_1241), .B2(n_1242), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_83), .A2(n_296), .B1(n_865), .B2(n_1178), .Y(n_1177) );
AOI22xp33_ASAP7_75t_SL g1190 ( .A1(n_83), .A2(n_296), .B1(n_986), .B2(n_1191), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_84), .A2(n_307), .B1(n_559), .B2(n_560), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1153 ( .A1(n_84), .A2(n_307), .B1(n_705), .B2(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1365 ( .A(n_85), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g1167 ( .A1(n_86), .A2(n_144), .B1(n_1124), .B2(n_1168), .Y(n_1167) );
OAI22xp33_ASAP7_75t_L g1200 ( .A1(n_86), .A2(n_144), .B1(n_1134), .B2(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1067 ( .A(n_87), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_87), .A2(n_259), .B1(n_391), .B2(n_1093), .C(n_1094), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_88), .A2(n_166), .B1(n_640), .B2(n_648), .C(n_742), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_88), .A2(n_166), .B1(n_698), .B2(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g1120 ( .A(n_89), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_89), .A2(n_105), .B1(n_1149), .B2(n_1151), .Y(n_1148) );
AO221x1_ASAP7_75t_L g1337 ( .A1(n_90), .A2(n_184), .B1(n_555), .B2(n_988), .C(n_1131), .Y(n_1337) );
INVx1_ASAP7_75t_L g1348 ( .A(n_90), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_91), .A2(n_245), .B1(n_585), .B2(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g929 ( .A(n_91), .Y(n_929) );
INVx1_ASAP7_75t_L g1730 ( .A(n_92), .Y(n_1730) );
AOI22xp33_ASAP7_75t_L g1753 ( .A1(n_92), .A2(n_209), .B1(n_1082), .B2(n_1299), .Y(n_1753) );
AOI221xp5_ASAP7_75t_L g1654 ( .A1(n_93), .A2(n_174), .B1(n_874), .B2(n_1178), .C(n_1655), .Y(n_1654) );
INVxp67_ASAP7_75t_SL g1696 ( .A(n_93), .Y(n_1696) );
INVx1_ASAP7_75t_L g1732 ( .A(n_94), .Y(n_1732) );
XNOR2x2_ASAP7_75t_L g1110 ( .A(n_96), .B(n_1111), .Y(n_1110) );
AO221x1_ASAP7_75t_L g1434 ( .A1(n_96), .A2(n_107), .B1(n_1435), .B2(n_1439), .C(n_1440), .Y(n_1434) );
AO221x1_ASAP7_75t_L g1458 ( .A1(n_97), .A2(n_282), .B1(n_1435), .B2(n_1439), .C(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1461 ( .A(n_98), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_100), .A2(n_253), .B1(n_865), .B2(n_1121), .Y(n_1317) );
AOI221xp5_ASAP7_75t_L g1334 ( .A1(n_100), .A2(n_253), .B1(n_421), .B2(n_423), .C(n_632), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g1747 ( .A1(n_101), .A2(n_187), .B1(n_1093), .B2(n_1094), .Y(n_1747) );
AOI22xp33_ASAP7_75t_L g1749 ( .A1(n_101), .A2(n_187), .B1(n_865), .B2(n_1178), .Y(n_1749) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_102), .A2(n_178), .B1(n_489), .B2(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g991 ( .A(n_102), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g1663 ( .A1(n_103), .A2(n_138), .B1(n_457), .B2(n_779), .C(n_1178), .Y(n_1663) );
INVx1_ASAP7_75t_L g1683 ( .A(n_103), .Y(n_1683) );
INVx1_ASAP7_75t_L g1442 ( .A(n_104), .Y(n_1442) );
INVx1_ASAP7_75t_L g1114 ( .A(n_105), .Y(n_1114) );
OA22x2_ASAP7_75t_L g1354 ( .A1(n_106), .A2(n_1355), .B1(n_1412), .B2(n_1413), .Y(n_1354) );
INVxp67_ASAP7_75t_SL g1413 ( .A(n_106), .Y(n_1413) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_108), .A2(n_134), .B1(n_1448), .B2(n_1451), .Y(n_1478) );
INVx1_ASAP7_75t_L g1041 ( .A(n_109), .Y(n_1041) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_109), .A2(n_183), .B1(n_997), .B2(n_999), .Y(n_1052) );
XNOR2xp5_ASAP7_75t_L g1058 ( .A(n_110), .B(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g669 ( .A(n_111), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_112), .A2(n_149), .B1(n_578), .B2(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g611 ( .A(n_112), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_113), .A2(n_266), .B1(n_986), .B2(n_987), .C(n_988), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_115), .Y(n_827) );
INVx1_ASAP7_75t_L g918 ( .A(n_116), .Y(n_918) );
INVx1_ASAP7_75t_L g1015 ( .A(n_117), .Y(n_1015) );
OAI221xp5_ASAP7_75t_L g1031 ( .A1(n_117), .A2(n_835), .B1(n_1032), .B2(n_1035), .C(n_1038), .Y(n_1031) );
INVx1_ASAP7_75t_L g1516 ( .A(n_118), .Y(n_1516) );
INVx1_ASAP7_75t_L g1279 ( .A(n_119), .Y(n_1279) );
AOI22xp33_ASAP7_75t_SL g1302 ( .A1(n_119), .A2(n_275), .B1(n_1178), .B2(n_1303), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_120), .A2(n_145), .B1(n_1082), .B2(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1203 ( .A(n_120), .Y(n_1203) );
INVx1_ASAP7_75t_L g1653 ( .A(n_121), .Y(n_1653) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_123), .A2(n_182), .B1(n_861), .B2(n_1082), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_123), .A2(n_182), .B1(n_810), .B2(n_811), .Y(n_1105) );
INVx1_ASAP7_75t_L g842 ( .A(n_124), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_124), .A2(n_257), .B1(n_861), .B2(n_862), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_125), .Y(n_1068) );
INVx1_ASAP7_75t_L g980 ( .A(n_126), .Y(n_980) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_126), .A2(n_266), .B1(n_997), .B2(n_999), .Y(n_996) );
INVx1_ASAP7_75t_L g1212 ( .A(n_127), .Y(n_1212) );
CKINVDCx5p33_ASAP7_75t_R g1366 ( .A(n_128), .Y(n_1366) );
INVx1_ASAP7_75t_L g1735 ( .A(n_129), .Y(n_1735) );
XOR2xp5_ASAP7_75t_L g730 ( .A(n_130), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g1423 ( .A(n_132), .Y(n_1423) );
INVx1_ASAP7_75t_L g1698 ( .A(n_135), .Y(n_1698) );
INVx1_ASAP7_75t_L g1460 ( .A(n_136), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g1643 ( .A1(n_136), .A2(n_1460), .B1(n_1644), .B2(n_1703), .Y(n_1643) );
AOI22xp33_ASAP7_75t_L g1709 ( .A1(n_136), .A2(n_1710), .B1(n_1754), .B2(n_1758), .Y(n_1709) );
INVx1_ASAP7_75t_L g1271 ( .A(n_137), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_137), .A2(n_176), .B1(n_485), .B2(n_583), .Y(n_1304) );
INVx1_ASAP7_75t_L g1680 ( .A(n_138), .Y(n_1680) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_140), .A2(n_271), .B1(n_373), .B2(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_140), .A2(n_271), .B1(n_443), .B2(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g853 ( .A(n_141), .Y(n_853) );
INVx1_ASAP7_75t_L g466 ( .A(n_142), .Y(n_466) );
INVx1_ASAP7_75t_L g634 ( .A(n_143), .Y(n_634) );
INVx1_ASAP7_75t_L g1204 ( .A(n_145), .Y(n_1204) );
INVx1_ASAP7_75t_L g1424 ( .A(n_146), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1444 ( .A(n_146), .B(n_1422), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1664 ( .A1(n_147), .A2(n_198), .B1(n_1665), .B2(n_1666), .Y(n_1664) );
INVx1_ASAP7_75t_L g1678 ( .A(n_147), .Y(n_1678) );
INVx1_ASAP7_75t_L g522 ( .A(n_148), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_148), .A2(n_170), .B1(n_564), .B2(n_567), .Y(n_563) );
INVx1_ASAP7_75t_L g592 ( .A(n_149), .Y(n_592) );
INVx2_ASAP7_75t_L g329 ( .A(n_150), .Y(n_329) );
XNOR2xp5_ASAP7_75t_L g1711 ( .A(n_151), .B(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1262 ( .A(n_152), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_153), .A2(n_190), .B1(n_1024), .B2(n_1026), .Y(n_1023) );
INVx1_ASAP7_75t_L g1048 ( .A(n_153), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1745 ( .A1(n_154), .A2(n_242), .B1(n_1189), .B2(n_1746), .Y(n_1745) );
AOI22xp33_ASAP7_75t_L g1750 ( .A1(n_154), .A2(n_242), .B1(n_1076), .B2(n_1082), .Y(n_1750) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_155), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_156), .A2(n_303), .B1(n_583), .B2(n_961), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_156), .A2(n_303), .B1(n_810), .B2(n_811), .Y(n_968) );
BUFx3_ASAP7_75t_L g355 ( .A(n_157), .Y(n_355) );
INVx1_ASAP7_75t_L g449 ( .A(n_157), .Y(n_449) );
INVx1_ASAP7_75t_L g974 ( .A(n_158), .Y(n_974) );
INVx1_ASAP7_75t_L g419 ( .A(n_159), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_159), .A2(n_239), .B1(n_457), .B2(n_459), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g1376 ( .A(n_160), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1340 ( .A(n_161), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g1367 ( .A(n_162), .Y(n_1367) );
INVxp33_ASAP7_75t_SL g737 ( .A(n_163), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_163), .A2(n_261), .B1(n_585), .B2(n_775), .C(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g1174 ( .A(n_164), .Y(n_1174) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_165), .A2(n_228), .B1(n_1168), .B2(n_1264), .C(n_1267), .Y(n_1263) );
INVx1_ASAP7_75t_L g1274 ( .A(n_165), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_167), .A2(n_216), .B1(n_794), .B2(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1017 ( .A(n_168), .Y(n_1017) );
OAI211xp5_ASAP7_75t_SL g1039 ( .A1(n_168), .A2(n_813), .B(n_1040), .C(n_1047), .Y(n_1039) );
CKINVDCx5p33_ASAP7_75t_R g1325 ( .A(n_169), .Y(n_1325) );
INVx1_ASAP7_75t_L g543 ( .A(n_170), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g1322 ( .A1(n_171), .A2(n_310), .B1(n_485), .B2(n_875), .Y(n_1322) );
INVx1_ASAP7_75t_L g1329 ( .A(n_171), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_172), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g893 ( .A1(n_173), .A2(n_186), .B1(n_690), .B2(n_693), .C(n_707), .Y(n_893) );
INVx1_ASAP7_75t_L g917 ( .A(n_173), .Y(n_917) );
INVxp67_ASAP7_75t_SL g1693 ( .A(n_174), .Y(n_1693) );
INVx1_ASAP7_75t_L g1470 ( .A(n_175), .Y(n_1470) );
INVx1_ASAP7_75t_L g1272 ( .A(n_176), .Y(n_1272) );
INVx1_ASAP7_75t_L g536 ( .A(n_177), .Y(n_536) );
INVx1_ASAP7_75t_L g990 ( .A(n_178), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_180), .Y(n_820) );
INVx1_ASAP7_75t_L g1517 ( .A(n_181), .Y(n_1517) );
INVx1_ASAP7_75t_L g1350 ( .A(n_184), .Y(n_1350) );
INVx1_ASAP7_75t_L g472 ( .A(n_185), .Y(n_472) );
INVx1_ASAP7_75t_L g915 ( .A(n_186), .Y(n_915) );
INVx1_ASAP7_75t_L g350 ( .A(n_188), .Y(n_350) );
INVx1_ASAP7_75t_L g441 ( .A(n_188), .Y(n_441) );
INVx1_ASAP7_75t_L g1649 ( .A(n_189), .Y(n_1649) );
INVx1_ASAP7_75t_L g1049 ( .A(n_190), .Y(n_1049) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_192), .Y(n_1387) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_193), .Y(n_674) );
INVx1_ASAP7_75t_L g412 ( .A(n_194), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_194), .A2(n_232), .B1(n_443), .B2(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g767 ( .A(n_195), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_196), .Y(n_829) );
XOR2x2_ASAP7_75t_L g806 ( .A(n_197), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g1684 ( .A(n_198), .Y(n_1684) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_199), .A2(n_286), .B1(n_1178), .B2(n_1319), .Y(n_1318) );
OAI221xp5_ASAP7_75t_L g1336 ( .A1(n_199), .A2(n_813), .B1(n_1337), .B2(n_1338), .C(n_1341), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_200), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g1171 ( .A(n_201), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_202), .Y(n_518) );
INVx1_ASAP7_75t_L g1441 ( .A(n_203), .Y(n_1441) );
XOR2xp5_ASAP7_75t_L g620 ( .A(n_204), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g1268 ( .A(n_205), .Y(n_1268) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_206), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_206), .A2(n_263), .B1(n_794), .B2(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g656 ( .A(n_207), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_207), .A2(n_215), .B1(n_705), .B2(n_707), .C(n_708), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g1492 ( .A1(n_208), .A2(n_311), .B1(n_1448), .B2(n_1451), .Y(n_1492) );
INVx1_ASAP7_75t_L g1729 ( .A(n_209), .Y(n_1729) );
INVx1_ASAP7_75t_L g637 ( .A(n_210), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_211), .A2(n_224), .B1(n_403), .B2(n_408), .Y(n_402) );
INVx1_ASAP7_75t_L g502 ( .A(n_211), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_212), .Y(n_507) );
INVx1_ASAP7_75t_L g1232 ( .A(n_213), .Y(n_1232) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_214), .Y(n_826) );
INVx1_ASAP7_75t_L g662 ( .A(n_215), .Y(n_662) );
INVx1_ASAP7_75t_L g1673 ( .A(n_217), .Y(n_1673) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_218), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_219), .A2(n_279), .B1(n_554), .B2(n_556), .Y(n_1145) );
AOI22xp33_ASAP7_75t_SL g1155 ( .A1(n_219), .A2(n_279), .B1(n_576), .B2(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g959 ( .A(n_220), .Y(n_959) );
OAI211xp5_ASAP7_75t_SL g977 ( .A1(n_220), .A2(n_813), .B(n_978), .C(n_989), .Y(n_977) );
INVx1_ASAP7_75t_L g955 ( .A(n_222), .Y(n_955) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_222), .A2(n_428), .B1(n_835), .B2(n_970), .C(n_975), .Y(n_969) );
INVx1_ASAP7_75t_L g1101 ( .A(n_223), .Y(n_1101) );
INVx1_ASAP7_75t_L g495 ( .A(n_224), .Y(n_495) );
INVx1_ASAP7_75t_L g539 ( .A(n_225), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_225), .A2(n_297), .B1(n_554), .B2(n_556), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_227), .A2(n_244), .B1(n_1359), .B2(n_1361), .Y(n_1358) );
INVx1_ASAP7_75t_L g1396 ( .A(n_227), .Y(n_1396) );
INVx1_ASAP7_75t_L g1275 ( .A(n_228), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_229), .Y(n_943) );
INVx1_ASAP7_75t_L g608 ( .A(n_230), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g812 ( .A1(n_231), .A2(n_813), .B1(n_814), .B2(n_822), .C(n_828), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_231), .A2(n_285), .B1(n_867), .B2(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g416 ( .A(n_232), .Y(n_416) );
INVx1_ASAP7_75t_L g910 ( .A(n_233), .Y(n_910) );
OAI211xp5_ASAP7_75t_L g1362 ( .A1(n_235), .A2(n_1099), .B(n_1285), .C(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1393 ( .A(n_235), .Y(n_1393) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_236), .Y(n_908) );
INVx1_ASAP7_75t_L g401 ( .A(n_239), .Y(n_401) );
BUFx3_ASAP7_75t_L g357 ( .A(n_240), .Y(n_357) );
INVx1_ASAP7_75t_L g445 ( .A(n_240), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g1324 ( .A(n_241), .Y(n_1324) );
AO22x2_ASAP7_75t_L g1254 ( .A1(n_243), .A2(n_1255), .B1(n_1305), .B2(n_1306), .Y(n_1254) );
INVxp67_ASAP7_75t_L g1305 ( .A(n_243), .Y(n_1305) );
INVx1_ASAP7_75t_L g1395 ( .A(n_244), .Y(n_1395) );
INVx1_ASAP7_75t_L g924 ( .A(n_245), .Y(n_924) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_246), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_246), .B(n_291), .Y(n_366) );
INVx1_ASAP7_75t_L g396 ( .A(n_246), .Y(n_396) );
AND2x2_ASAP7_75t_L g400 ( .A(n_246), .B(n_395), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g1339 ( .A(n_247), .Y(n_1339) );
INVx1_ASAP7_75t_L g1136 ( .A(n_249), .Y(n_1136) );
XNOR2xp5_ASAP7_75t_L g1161 ( .A(n_250), .B(n_1162), .Y(n_1161) );
INVx2_ASAP7_75t_L g352 ( .A(n_251), .Y(n_352) );
OR2x2_ASAP7_75t_L g470 ( .A(n_251), .B(n_350), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_252), .Y(n_909) );
INVx1_ASAP7_75t_L g849 ( .A(n_254), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_255), .Y(n_1381) );
INVx1_ASAP7_75t_L g1115 ( .A(n_256), .Y(n_1115) );
INVx1_ASAP7_75t_L g839 ( .A(n_257), .Y(n_839) );
INVx1_ASAP7_75t_L g761 ( .A(n_258), .Y(n_761) );
INVx1_ASAP7_75t_L g1065 ( .A(n_259), .Y(n_1065) );
INVxp33_ASAP7_75t_L g739 ( .A(n_261), .Y(n_739) );
INVx1_ASAP7_75t_L g1726 ( .A(n_262), .Y(n_1726) );
AOI22xp33_ASAP7_75t_L g1741 ( .A1(n_262), .A2(n_273), .B1(n_1182), .B2(n_1742), .Y(n_1741) );
INVxp33_ASAP7_75t_L g745 ( .A(n_263), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_264), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_265), .A2(n_281), .B1(n_1178), .B2(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1206 ( .A(n_265), .Y(n_1206) );
AOI22x1_ASAP7_75t_L g1309 ( .A1(n_267), .A2(n_1310), .B1(n_1311), .B2(n_1351), .Y(n_1309) );
INVxp67_ASAP7_75t_SL g1351 ( .A(n_267), .Y(n_1351) );
INVx1_ASAP7_75t_L g1722 ( .A(n_268), .Y(n_1722) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_269), .A2(n_293), .B1(n_1019), .B2(n_1021), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_269), .A2(n_293), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
INVx1_ASAP7_75t_L g1002 ( .A(n_270), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_272), .Y(n_1072) );
INVx1_ASAP7_75t_L g1725 ( .A(n_273), .Y(n_1725) );
INVx1_ASAP7_75t_L g1132 ( .A(n_274), .Y(n_1132) );
INVx1_ASAP7_75t_L g1284 ( .A(n_275), .Y(n_1284) );
INVx1_ASAP7_75t_L g1045 ( .A(n_276), .Y(n_1045) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_277), .Y(n_1117) );
INVx1_ASAP7_75t_L g1104 ( .A(n_280), .Y(n_1104) );
INVx1_ASAP7_75t_L g1199 ( .A(n_281), .Y(n_1199) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_283), .B(n_317), .Y(n_1420) );
AND3x2_ASAP7_75t_L g1438 ( .A(n_283), .B(n_317), .C(n_1423), .Y(n_1438) );
INVx2_ASAP7_75t_L g330 ( .A(n_284), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g834 ( .A1(n_285), .A2(n_428), .B1(n_835), .B2(n_836), .C(n_843), .Y(n_834) );
INVx1_ASAP7_75t_L g1335 ( .A(n_286), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g1214 ( .A(n_287), .Y(n_1214) );
INVx1_ASAP7_75t_L g1122 ( .A(n_288), .Y(n_1122) );
INVx1_ASAP7_75t_L g1084 ( .A(n_289), .Y(n_1084) );
INVx1_ASAP7_75t_L g1170 ( .A(n_290), .Y(n_1170) );
INVx1_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
INVx2_ASAP7_75t_L g395 ( .A(n_291), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_294), .Y(n_1357) );
INVx1_ASAP7_75t_L g770 ( .A(n_295), .Y(n_770) );
INVx1_ASAP7_75t_L g528 ( .A(n_297), .Y(n_528) );
OAI211xp5_ASAP7_75t_L g1371 ( .A1(n_298), .A2(n_1216), .B(n_1372), .C(n_1374), .Y(n_1371) );
INVx1_ASAP7_75t_L g1410 ( .A(n_298), .Y(n_1410) );
INVx1_ASAP7_75t_L g1662 ( .A(n_299), .Y(n_1662) );
INVxp33_ASAP7_75t_SL g735 ( .A(n_300), .Y(n_735) );
OAI211xp5_ASAP7_75t_SL g1086 ( .A1(n_302), .A2(n_813), .B(n_1087), .C(n_1096), .Y(n_1086) );
INVxp33_ASAP7_75t_SL g749 ( .A(n_304), .Y(n_749) );
INVx1_ASAP7_75t_L g1009 ( .A(n_305), .Y(n_1009) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_306), .Y(n_832) );
INVx1_ASAP7_75t_L g1648 ( .A(n_308), .Y(n_1648) );
INVxp33_ASAP7_75t_SL g1036 ( .A(n_309), .Y(n_1036) );
INVx1_ASAP7_75t_L g1330 ( .A(n_310), .Y(n_1330) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_333), .B(n_1414), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_320), .Y(n_314) );
AND2x4_ASAP7_75t_L g1708 ( .A(n_315), .B(n_321), .Y(n_1708) );
NOR2xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_SL g1757 ( .A(n_316), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_316), .B(n_318), .Y(n_1760) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_318), .B(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g614 ( .A(n_323), .B(n_346), .Y(n_614) );
OR2x6_ASAP7_75t_L g1142 ( .A(n_323), .B(n_346), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g552 ( .A(n_324), .B(n_332), .Y(n_552) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g423 ( .A(n_325), .B(n_424), .Y(n_423) );
INVx8_ASAP7_75t_L g610 ( .A(n_326), .Y(n_610) );
OR2x6_ASAP7_75t_L g326 ( .A(n_327), .B(n_331), .Y(n_326) );
OR2x6_ASAP7_75t_L g613 ( .A(n_327), .B(n_603), .Y(n_613) );
INVx1_ASAP7_75t_L g655 ( .A(n_327), .Y(n_655) );
OR2x2_ASAP7_75t_L g728 ( .A(n_327), .B(n_644), .Y(n_728) );
INVx2_ASAP7_75t_SL g748 ( .A(n_327), .Y(n_748) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_327), .Y(n_819) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g369 ( .A(n_329), .B(n_330), .Y(n_369) );
INVx2_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
AND2x4_ASAP7_75t_L g381 ( .A(n_329), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g390 ( .A(n_329), .Y(n_390) );
INVx1_ASAP7_75t_L g432 ( .A(n_329), .Y(n_432) );
INVx1_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
INVx2_ASAP7_75t_L g382 ( .A(n_330), .Y(n_382) );
INVx1_ASAP7_75t_L g406 ( .A(n_330), .Y(n_406) );
INVx1_ASAP7_75t_L g431 ( .A(n_330), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_330), .B(n_375), .Y(n_668) );
AND2x4_ASAP7_75t_L g598 ( .A(n_331), .B(n_406), .Y(n_598) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g599 ( .A(n_332), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g1134 ( .A(n_332), .B(n_600), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_1053), .B2(n_1054), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
XNOR2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_802), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_618), .B1(n_800), .B2(n_801), .Y(n_336) );
INVx1_ASAP7_75t_L g800 ( .A(n_337), .Y(n_800) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI21x1_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_508), .B(n_617), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g617 ( .A(n_340), .B(n_509), .Y(n_617) );
XOR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_507), .Y(n_340) );
NOR3xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_370), .C(n_435), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_344), .B(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_344), .B(n_966), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_344), .B(n_1005), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_344), .B(n_1084), .Y(n_1083) );
OR2x6_ASAP7_75t_L g344 ( .A(n_345), .B(n_358), .Y(n_344) );
INVx2_ASAP7_75t_L g729 ( .A(n_345), .Y(n_729) );
AOI222xp33_ASAP7_75t_L g1347 ( .A1(n_345), .A2(n_467), .B1(n_481), .B2(n_1339), .C1(n_1342), .C2(n_1348), .Y(n_1347) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AND2x4_ASAP7_75t_L g463 ( .A(n_346), .B(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g589 ( .A(n_346), .B(n_464), .Y(n_589) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_353), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_348), .B(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g699 ( .A(n_348), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g702 ( .A(n_348), .B(n_491), .Y(n_702) );
INVx1_ASAP7_75t_L g717 ( .A(n_348), .Y(n_717) );
BUFx2_ASAP7_75t_L g1659 ( .A(n_348), .Y(n_1659) );
AND2x4_ASAP7_75t_L g1670 ( .A(n_348), .B(n_700), .Y(n_1670) );
AND2x4_ASAP7_75t_L g1672 ( .A(n_348), .B(n_491), .Y(n_1672) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g464 ( .A(n_351), .B(n_441), .Y(n_464) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g440 ( .A(n_352), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g516 ( .A(n_352), .Y(n_516) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_352), .Y(n_521) );
INVx1_ASAP7_75t_L g525 ( .A(n_352), .Y(n_525) );
BUFx2_ASAP7_75t_L g451 ( .A(n_353), .Y(n_451) );
INVx2_ASAP7_75t_L g458 ( .A(n_353), .Y(n_458) );
AND2x4_ASAP7_75t_L g519 ( .A(n_353), .B(n_520), .Y(n_519) );
INVx6_ASAP7_75t_L g542 ( .A(n_353), .Y(n_542) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g492 ( .A(n_354), .Y(n_492) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g444 ( .A(n_355), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g455 ( .A(n_355), .B(n_357), .Y(n_455) );
INVx1_ASAP7_75t_L g500 ( .A(n_356), .Y(n_500) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g448 ( .A(n_357), .B(n_449), .Y(n_448) );
NOR2xp67_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
INVx2_ASAP7_75t_L g434 ( .A(n_359), .Y(n_434) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g438 ( .A(n_360), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g551 ( .A(n_360), .B(n_552), .Y(n_551) );
OR2x6_ASAP7_75t_L g573 ( .A(n_360), .B(n_574), .Y(n_573) );
OAI31xp33_ASAP7_75t_L g808 ( .A1(n_360), .A2(n_809), .A3(n_812), .B(n_834), .Y(n_808) );
BUFx2_ASAP7_75t_L g992 ( .A(n_360), .Y(n_992) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_360), .B(n_552), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_360), .B(n_574), .Y(n_1315) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g547 ( .A(n_361), .Y(n_547) );
OR2x6_ASAP7_75t_L g651 ( .A(n_361), .B(n_423), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_367), .Y(n_362) );
AND2x2_ASAP7_75t_L g830 ( .A(n_363), .B(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
OR2x6_ASAP7_75t_L g408 ( .A(n_364), .B(n_409), .Y(n_408) );
OR2x6_ASAP7_75t_L g428 ( .A(n_364), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_364), .B(n_429), .Y(n_1038) );
INVx1_ASAP7_75t_L g1345 ( .A(n_364), .Y(n_1345) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g986 ( .A(n_367), .Y(n_986) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g555 ( .A(n_368), .Y(n_555) );
INVx2_ASAP7_75t_SL g636 ( .A(n_368), .Y(n_636) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_369), .Y(n_385) );
AOI31xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_410), .A3(n_417), .B(n_433), .Y(n_370) );
AOI221xp5_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_383), .B1(n_397), .B2(n_401), .C(n_402), .Y(n_371) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g411 ( .A(n_374), .B(n_400), .Y(n_411) );
BUFx2_ASAP7_75t_L g559 ( .A(n_374), .Y(n_559) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_374), .Y(n_566) );
AND2x4_ASAP7_75t_L g602 ( .A(n_374), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g1183 ( .A(n_374), .Y(n_1183) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_374), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g1333 ( .A(n_374), .Y(n_1333) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g757 ( .A(n_379), .Y(n_757) );
INVx2_ASAP7_75t_L g1185 ( .A(n_379), .Y(n_1185) );
INVx2_ASAP7_75t_L g1291 ( .A(n_379), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_379), .B(n_629), .Y(n_1679) );
INVx2_ASAP7_75t_L g1743 ( .A(n_379), .Y(n_1743) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g628 ( .A(n_380), .Y(n_628) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_380), .Y(n_764) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_381), .Y(n_562) );
INVx1_ASAP7_75t_L g607 ( .A(n_381), .Y(n_607) );
AND2x4_ASAP7_75t_L g389 ( .A(n_382), .B(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g418 ( .A(n_385), .B(n_400), .Y(n_418) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
INVx3_ASAP7_75t_L g1095 ( .A(n_385), .Y(n_1095) );
AOI211xp5_ASAP7_75t_L g591 ( .A1(n_386), .A2(n_592), .B(n_593), .C(n_596), .Y(n_591) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g1093 ( .A(n_387), .Y(n_1093) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g397 ( .A(n_388), .B(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_389), .Y(n_422) );
AND2x4_ASAP7_75t_L g593 ( .A(n_389), .B(n_594), .Y(n_593) );
BUFx3_ASAP7_75t_L g632 ( .A(n_389), .Y(n_632) );
BUFx6f_ASAP7_75t_L g1131 ( .A(n_389), .Y(n_1131) );
BUFx2_ASAP7_75t_L g1282 ( .A(n_389), .Y(n_1282) );
INVx1_ASAP7_75t_L g821 ( .A(n_391), .Y(n_821) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g570 ( .A(n_393), .B(n_494), .Y(n_570) );
BUFx2_ASAP7_75t_L g988 ( .A(n_393), .Y(n_988) );
NAND2x1p5_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g595 ( .A(n_394), .Y(n_595) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
INVx8_ASAP7_75t_L g813 ( .A(n_397), .Y(n_813) );
AND2x4_ASAP7_75t_L g413 ( .A(n_398), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g629 ( .A(n_400), .B(n_471), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
NAND2x1_ASAP7_75t_SL g642 ( .A(n_404), .B(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g1344 ( .A1(n_404), .A2(n_1277), .B1(n_1324), .B2(n_1325), .Y(n_1344) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_406), .Y(n_831) );
CKINVDCx11_ASAP7_75t_R g833 ( .A(n_408), .Y(n_833) );
INVx1_ASAP7_75t_L g647 ( .A(n_409), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_413), .B2(n_416), .Y(n_410) );
INVx3_ASAP7_75t_L g810 ( .A(n_411), .Y(n_810) );
INVx3_ASAP7_75t_L g1029 ( .A(n_411), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_411), .A2(n_413), .B1(n_1329), .B2(n_1330), .Y(n_1328) );
INVx3_ASAP7_75t_L g811 ( .A(n_413), .Y(n_811) );
INVx3_ASAP7_75t_L g1030 ( .A(n_413), .Y(n_1030) );
INVx1_ASAP7_75t_L g1044 ( .A(n_414), .Y(n_1044) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g426 ( .A(n_415), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_425), .C(n_427), .Y(n_417) );
CKINVDCx6p67_ASAP7_75t_R g835 ( .A(n_418), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_418), .A2(n_1332), .B1(n_1334), .B2(n_1335), .Y(n_1331) );
INVx1_ASAP7_75t_L g1150 ( .A(n_421), .Y(n_1150) );
INVx2_ASAP7_75t_SL g557 ( .A(n_422), .Y(n_557) );
BUFx6f_ASAP7_75t_L g987 ( .A(n_422), .Y(n_987) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_422), .B(n_629), .Y(n_1681) );
INVx1_ASAP7_75t_L g603 ( .A(n_424), .Y(n_603) );
INVx1_ASAP7_75t_L g983 ( .A(n_426), .Y(n_983) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_429), .Y(n_750) );
INVx1_ASAP7_75t_L g845 ( .A(n_429), .Y(n_845) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g680 ( .A(n_430), .Y(n_680) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_430), .Y(n_1034) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_431), .B(n_432), .Y(n_660) );
INVx1_ASAP7_75t_L g600 ( .A(n_432), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_433), .A2(n_685), .B1(n_725), .B2(n_726), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_433), .A2(n_726), .B1(n_772), .B2(n_798), .Y(n_771) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI31xp33_ASAP7_75t_L g1027 ( .A1(n_434), .A2(n_1028), .A3(n_1031), .B(n_1039), .Y(n_1027) );
NAND4xp25_ASAP7_75t_L g435 ( .A(n_436), .B(n_465), .C(n_479), .D(n_487), .Y(n_435) );
AOI33xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_442), .A3(n_450), .B1(n_456), .B2(n_461), .B3(n_463), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g1176 ( .A(n_437), .B(n_1177), .C(n_1179), .Y(n_1176) );
NAND3xp33_ASAP7_75t_L g1297 ( .A(n_437), .B(n_1298), .C(n_1300), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1748 ( .A(n_437), .B(n_1749), .C(n_1750), .Y(n_1748) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g574 ( .A(n_440), .Y(n_574) );
INVx2_ASAP7_75t_SL g710 ( .A(n_440), .Y(n_710) );
INVx1_ASAP7_75t_L g792 ( .A(n_440), .Y(n_792) );
BUFx3_ASAP7_75t_L g1656 ( .A(n_440), .Y(n_1656) );
INVx1_ASAP7_75t_L g546 ( .A(n_441), .Y(n_546) );
BUFx3_ASAP7_75t_L g582 ( .A(n_443), .Y(n_582) );
AND2x4_ASAP7_75t_L g687 ( .A(n_443), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g782 ( .A(n_443), .Y(n_782) );
INVx2_ASAP7_75t_SL g790 ( .A(n_443), .Y(n_790) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g486 ( .A(n_444), .Y(n_486) );
AND2x6_ASAP7_75t_L g544 ( .A(n_444), .B(n_515), .Y(n_544) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_444), .Y(n_588) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_444), .Y(n_706) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_444), .Y(n_874) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_444), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1076 ( .A(n_444), .Y(n_1076) );
BUFx2_ASAP7_75t_L g1299 ( .A(n_444), .Y(n_1299) );
HB1xp67_ASAP7_75t_L g1665 ( .A(n_444), .Y(n_1665) );
INVx1_ASAP7_75t_L g478 ( .A(n_445), .Y(n_478) );
BUFx2_ASAP7_75t_L g696 ( .A(n_446), .Y(n_696) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g468 ( .A(n_447), .B(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g995 ( .A(n_447), .B(n_469), .Y(n_995) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_448), .Y(n_462) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_448), .Y(n_526) );
INVx2_ASAP7_75t_L g724 ( .A(n_448), .Y(n_724) );
INVx1_ASAP7_75t_L g796 ( .A(n_448), .Y(n_796) );
INVx1_ASAP7_75t_L g477 ( .A(n_449), .Y(n_477) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g1178 ( .A(n_453), .Y(n_1178) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g505 ( .A(n_454), .Y(n_505) );
AND2x4_ASAP7_75t_L g513 ( .A(n_454), .B(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_454), .Y(n_530) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_454), .Y(n_580) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_455), .Y(n_460) );
AND2x2_ASAP7_75t_L g481 ( .A(n_457), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g585 ( .A(n_458), .Y(n_585) );
BUFx2_ASAP7_75t_SL g791 ( .A(n_459), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_459), .B(n_506), .Y(n_880) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g714 ( .A(n_460), .B(n_688), .Y(n_714) );
INVx2_ASAP7_75t_SL g868 ( .A(n_460), .Y(n_868) );
BUFx4f_ASAP7_75t_L g1121 ( .A(n_460), .Y(n_1121) );
BUFx3_ASAP7_75t_L g1244 ( .A(n_460), .Y(n_1244) );
AND2x4_ASAP7_75t_L g1658 ( .A(n_460), .B(n_1659), .Y(n_1658) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_462), .Y(n_583) );
BUFx3_ASAP7_75t_L g905 ( .A(n_462), .Y(n_905) );
INVx1_ASAP7_75t_L g950 ( .A(n_462), .Y(n_950) );
INVx1_ASAP7_75t_L g877 ( .A(n_463), .Y(n_877) );
AOI33xp33_ASAP7_75t_L g1073 ( .A1(n_463), .A2(n_1074), .A3(n_1075), .B1(n_1078), .B2(n_1080), .B3(n_1081), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g1192 ( .A(n_463), .B(n_1193), .C(n_1195), .Y(n_1192) );
NAND3xp33_ASAP7_75t_L g1301 ( .A(n_463), .B(n_1302), .C(n_1304), .Y(n_1301) );
AOI33xp33_ASAP7_75t_L g1313 ( .A1(n_463), .A2(n_1314), .A3(n_1316), .B1(n_1317), .B2(n_1318), .B3(n_1322), .Y(n_1313) );
INVx2_ASAP7_75t_L g694 ( .A(n_464), .Y(n_694) );
INVx2_ASAP7_75t_SL g779 ( .A(n_464), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_472), .B2(n_473), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_467), .A2(n_473), .B1(n_816), .B2(n_827), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_467), .A2(n_473), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
CKINVDCx6p67_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_L g474 ( .A(n_469), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g482 ( .A(n_469), .Y(n_482) );
OR2x2_ASAP7_75t_L g997 ( .A(n_469), .B(n_998), .Y(n_997) );
OR2x2_ASAP7_75t_L g999 ( .A(n_469), .B(n_1000), .Y(n_999) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g688 ( .A(n_470), .Y(n_688) );
OR2x2_ASAP7_75t_L g720 ( .A(n_470), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g723 ( .A(n_470), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g494 ( .A(n_471), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g1349 ( .A1(n_473), .A2(n_484), .B1(n_1340), .B2(n_1350), .Y(n_1349) );
CKINVDCx6p67_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g1392 ( .A(n_475), .Y(n_1392) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx4f_ASAP7_75t_L g947 ( .A(n_476), .Y(n_947) );
INVx1_ASAP7_75t_L g958 ( .A(n_476), .Y(n_958) );
INVx1_ASAP7_75t_L g1720 ( .A(n_476), .Y(n_1720) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
OR2x2_ASAP7_75t_L g721 ( .A(n_477), .B(n_478), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_483), .B2(n_484), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_481), .A2(n_484), .B1(n_820), .B2(n_826), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_481), .A2(n_484), .B1(n_1067), .B2(n_1068), .Y(n_1066) );
AND2x2_ASAP7_75t_L g484 ( .A(n_482), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g1196 ( .A(n_486), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_486), .A2(n_1395), .B1(n_1396), .B2(n_1397), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_495), .B1(n_496), .B2(n_502), .C(n_503), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_488), .A2(n_829), .B1(n_832), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_488), .A2(n_1025), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_488), .A2(n_496), .B1(n_503), .B2(n_1324), .C(n_1325), .Y(n_1323) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .Y(n_489) );
OR2x2_ASAP7_75t_L g786 ( .A(n_490), .B(n_717), .Y(n_786) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_490), .B(n_493), .Y(n_1026) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x6_ASAP7_75t_L g537 ( .A(n_492), .B(n_516), .Y(n_537) );
INVx2_ASAP7_75t_SL g501 ( .A(n_493), .Y(n_501) );
INVx1_ASAP7_75t_L g506 ( .A(n_493), .Y(n_506) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g857 ( .A(n_497), .Y(n_857) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_497), .Y(n_964) );
INVx1_ASAP7_75t_L g1025 ( .A(n_497), .Y(n_1025) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g700 ( .A(n_499), .Y(n_700) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g535 ( .A(n_500), .Y(n_535) );
BUFx2_ASAP7_75t_L g937 ( .A(n_503), .Y(n_937) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g707 ( .A(n_505), .Y(n_707) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g616 ( .A(n_510), .Y(n_616) );
AOI211x1_ASAP7_75t_SL g510 ( .A1(n_511), .A2(n_545), .B(n_548), .C(n_590), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_512), .B(n_517), .C(n_527), .D(n_538), .Y(n_511) );
NAND4xp25_ASAP7_75t_SL g1112 ( .A(n_512), .B(n_1113), .C(n_1116), .D(n_1119), .Y(n_1112) );
INVx5_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g1164 ( .A1(n_513), .A2(n_1165), .B(n_1166), .C(n_1167), .Y(n_1164) );
CKINVDCx8_ASAP7_75t_R g1216 ( .A(n_513), .Y(n_1216) );
NOR2xp33_ASAP7_75t_L g1715 ( .A(n_513), .B(n_1716), .Y(n_1715) );
OAI21xp33_ASAP7_75t_L g1267 ( .A1(n_514), .A2(n_580), .B(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g1222 ( .A(n_515), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_515), .B(n_530), .Y(n_1373) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_522), .B2(n_523), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_518), .A2(n_610), .B1(n_611), .B2(n_612), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_519), .A2(n_523), .B1(n_1117), .B2(n_1118), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_519), .A2(n_540), .B1(n_1170), .B2(n_1171), .Y(n_1169) );
INVx4_ASAP7_75t_L g1223 ( .A(n_519), .Y(n_1223) );
AOI221xp5_ASAP7_75t_L g1260 ( .A1(n_519), .A2(n_544), .B1(n_1261), .B2(n_1262), .C(n_1263), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1721 ( .A1(n_519), .A2(n_540), .B1(n_1722), .B2(n_1723), .Y(n_1721) );
AND2x4_ASAP7_75t_L g533 ( .A(n_520), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_SL g1377 ( .A(n_520), .B(n_534), .Y(n_1377) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_523), .A2(n_544), .B1(n_1173), .B2(n_1174), .Y(n_1172) );
INVx4_ASAP7_75t_L g1219 ( .A(n_523), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_523), .A2(n_540), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1724 ( .A1(n_523), .A2(n_544), .B1(n_1725), .B2(n_1726), .Y(n_1724) );
AND2x6_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
AND2x4_ASAP7_75t_L g540 ( .A(n_524), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_525), .B(n_1266), .Y(n_1265) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_526), .Y(n_712) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_526), .Y(n_875) );
INVx2_ASAP7_75t_L g1022 ( .A(n_526), .Y(n_1022) );
INVx1_ASAP7_75t_L g1397 ( .A(n_526), .Y(n_1397) );
INVx1_ASAP7_75t_L g1667 ( .A(n_526), .Y(n_1667) );
AOI222xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B1(n_531), .B2(n_532), .C1(n_536), .C2(n_537), .Y(n_527) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_530), .Y(n_692) );
HB1xp67_ASAP7_75t_L g1166 ( .A(n_530), .Y(n_1166) );
BUFx4f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g1124 ( .A(n_533), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_533), .A2(n_537), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g1266 ( .A(n_535), .Y(n_1266) );
AOI222xp33_ASAP7_75t_L g1119 ( .A1(n_537), .A2(n_1120), .B1(n_1121), .B2(n_1122), .C1(n_1123), .C2(n_1125), .Y(n_1119) );
INVx3_ASAP7_75t_L g1168 ( .A(n_537), .Y(n_1168) );
AOI322xp5_ASAP7_75t_L g1374 ( .A1(n_537), .A2(n_874), .A3(n_1366), .B1(n_1367), .B2(n_1375), .C1(n_1376), .C2(n_1377), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_543), .B2(n_544), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_540), .A2(n_544), .B1(n_1114), .B2(n_1115), .Y(n_1113) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g577 ( .A(n_542), .Y(n_577) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_542), .Y(n_691) );
INVx2_ASAP7_75t_L g866 ( .A(n_542), .Y(n_866) );
INVx1_ASAP7_75t_L g1303 ( .A(n_542), .Y(n_1303) );
INVx2_ASAP7_75t_SL g1321 ( .A(n_542), .Y(n_1321) );
CKINVDCx6p67_ASAP7_75t_R g1218 ( .A(n_544), .Y(n_1218) );
BUFx6f_ASAP7_75t_L g1126 ( .A(n_545), .Y(n_1126) );
AO211x2_ASAP7_75t_L g1162 ( .A1(n_545), .A2(n_1163), .B(n_1175), .C(n_1197), .Y(n_1162) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_546), .B(n_547), .Y(n_1224) );
INVx2_ASAP7_75t_L g890 ( .A(n_547), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_571), .Y(n_548) );
AOI33xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_553), .A3(n_558), .B1(n_563), .B2(n_568), .B3(n_569), .Y(n_549) );
AOI33xp33_ASAP7_75t_L g1144 ( .A1(n_550), .A2(n_569), .A3(n_1145), .B1(n_1146), .B2(n_1147), .B3(n_1148), .Y(n_1144) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g1187 ( .A(n_551), .B(n_1188), .C(n_1190), .Y(n_1187) );
INVx1_ASAP7_75t_L g851 ( .A(n_552), .Y(n_851) );
BUFx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI211xp5_ASAP7_75t_L g1198 ( .A1(n_556), .A2(n_593), .B(n_1199), .C(n_1200), .Y(n_1198) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g1151 ( .A(n_557), .Y(n_1151) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_561), .A2(n_663), .B1(n_897), .B2(n_909), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_561), .A2(n_824), .B1(n_1036), .B2(n_1037), .Y(n_1035) );
INVx4_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx3_ASAP7_75t_L g567 ( .A(n_562), .Y(n_567) );
INVx2_ASAP7_75t_SL g675 ( .A(n_562), .Y(n_675) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g638 ( .A(n_566), .B(n_629), .Y(n_638) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_566), .B(n_629), .Y(n_1685) );
AOI33xp33_ASAP7_75t_L g1233 ( .A1(n_569), .A2(n_1234), .A3(n_1235), .B1(n_1236), .B2(n_1237), .B3(n_1238), .Y(n_1233) );
INVx2_ASAP7_75t_L g1411 ( .A(n_569), .Y(n_1411) );
INVx6_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx5_ASAP7_75t_L g683 ( .A(n_570), .Y(n_683) );
AOI33xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .A3(n_581), .B1(n_584), .B2(n_586), .B3(n_589), .Y(n_571) );
AOI33xp33_ASAP7_75t_L g1152 ( .A1(n_572), .A2(n_1153), .A3(n_1155), .B1(n_1157), .B2(n_1158), .B3(n_1159), .Y(n_1152) );
AOI33xp33_ASAP7_75t_L g1239 ( .A1(n_572), .A2(n_589), .A3(n_1240), .B1(n_1243), .B2(n_1245), .B3(n_1247), .Y(n_1239) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_573), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_573), .Y(n_859) );
OAI22xp5_ASAP7_75t_SL g938 ( .A1(n_573), .A2(n_939), .B1(n_951), .B2(n_952), .Y(n_938) );
OAI22xp5_ASAP7_75t_SL g1007 ( .A1(n_573), .A2(n_1008), .B1(n_1012), .B2(n_1014), .Y(n_1007) );
INVx2_ASAP7_75t_L g1074 ( .A(n_573), .Y(n_1074) );
BUFx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_577), .Y(n_794) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g715 ( .A(n_580), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g776 ( .A(n_580), .Y(n_776) );
INVx1_ASAP7_75t_L g903 ( .A(n_580), .Y(n_903) );
BUFx6f_ASAP7_75t_L g1246 ( .A(n_580), .Y(n_1246) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx4f_ASAP7_75t_L g861 ( .A(n_588), .Y(n_861) );
INVx1_ASAP7_75t_L g1000 ( .A(n_588), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_588), .B(n_688), .Y(n_1661) );
INVx4_ASAP7_75t_L g951 ( .A(n_589), .Y(n_951) );
BUFx4f_ASAP7_75t_L g1013 ( .A(n_589), .Y(n_1013) );
BUFx4f_ASAP7_75t_L g1159 ( .A(n_589), .Y(n_1159) );
AOI31xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_601), .A3(n_609), .B(n_614), .Y(n_590) );
AOI211xp5_ASAP7_75t_L g1128 ( .A1(n_593), .A2(n_1129), .B(n_1132), .C(n_1133), .Y(n_1128) );
NOR3xp33_ASAP7_75t_L g1226 ( .A(n_593), .B(n_1227), .C(n_1229), .Y(n_1226) );
CKINVDCx11_ASAP7_75t_R g1285 ( .A(n_593), .Y(n_1285) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVxp67_ASAP7_75t_L g1278 ( .A(n_595), .Y(n_1278) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g1201 ( .A(n_598), .Y(n_1201) );
INVx2_ASAP7_75t_L g1228 ( .A(n_598), .Y(n_1228) );
AOI222xp33_ASAP7_75t_L g1273 ( .A1(n_598), .A2(n_1274), .B1(n_1275), .B2(n_1276), .C1(n_1279), .C2(n_1280), .Y(n_1273) );
AOI322xp5_ASAP7_75t_L g1363 ( .A1(n_598), .A2(n_1276), .A3(n_1360), .B1(n_1364), .B2(n_1365), .C1(n_1366), .C2(n_1367), .Y(n_1363) );
INVx1_ASAP7_75t_L g1277 ( .A(n_600), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .B1(n_605), .B2(n_608), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_602), .A2(n_1136), .B1(n_1137), .B2(n_1138), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g1202 ( .A1(n_602), .A2(n_605), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_602), .A2(n_605), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_602), .A2(n_1137), .B1(n_1271), .B2(n_1272), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1728 ( .A1(n_602), .A2(n_1137), .B1(n_1729), .B2(n_1730), .Y(n_1728) );
AND2x4_ASAP7_75t_L g605 ( .A(n_603), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g1137 ( .A(n_603), .B(n_606), .Y(n_1137) );
INVx1_ASAP7_75t_L g1360 ( .A(n_603), .Y(n_1360) );
INVx5_ASAP7_75t_SL g1361 ( .A(n_605), .Y(n_1361) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_607), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_610), .A2(n_1117), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g1205 ( .A1(n_610), .A2(n_612), .B1(n_1171), .B2(n_1206), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_610), .A2(n_1141), .B1(n_1261), .B2(n_1284), .Y(n_1283) );
AOI211xp5_ASAP7_75t_L g1356 ( .A1(n_610), .A2(n_1357), .B(n_1358), .C(n_1362), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g1736 ( .A1(n_610), .A2(n_612), .B1(n_1723), .B2(n_1737), .Y(n_1736) );
INVx5_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx4_ASAP7_75t_L g1141 ( .A(n_613), .Y(n_1141) );
OAI211xp5_ASAP7_75t_L g1355 ( .A1(n_614), .A2(n_1356), .B(n_1368), .C(n_1378), .Y(n_1355) );
INVx1_ASAP7_75t_L g801 ( .A(n_618), .Y(n_801) );
AO22x2_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B1(n_730), .B2(n_799), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_684), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_639), .C(n_650), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_633), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_630), .B2(n_631), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_626), .A2(n_631), .B1(n_914), .B2(n_915), .Y(n_913) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g736 ( .A(n_627), .Y(n_736) );
AND2x4_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx2_ASAP7_75t_L g1697 ( .A(n_628), .Y(n_1697) );
AND2x6_ASAP7_75t_L g631 ( .A(n_629), .B(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_L g635 ( .A(n_629), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_631), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g649 ( .A(n_632), .B(n_643), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_637), .B2(n_638), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_635), .A2(n_638), .B1(n_739), .B2(n_740), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_635), .A2(n_638), .B1(n_917), .B2(n_918), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g1682 ( .A1(n_635), .A2(n_1683), .B1(n_1684), .B2(n_1685), .Y(n_1682) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g1687 ( .A(n_641), .Y(n_1687) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_643), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx4f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx4f_ASAP7_75t_L g742 ( .A(n_646), .Y(n_742) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx3_ASAP7_75t_L g1688 ( .A(n_649), .Y(n_1688) );
OAI33xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .A3(n_661), .B1(n_673), .B2(n_677), .B3(n_682), .Y(n_650) );
OAI33xp33_ASAP7_75t_L g743 ( .A1(n_651), .A2(n_682), .A3(n_744), .B1(n_751), .B2(n_758), .B3(n_766), .Y(n_743) );
INVx1_ASAP7_75t_L g922 ( .A(n_651), .Y(n_922) );
OAI33xp33_ASAP7_75t_L g1398 ( .A1(n_651), .A2(n_1399), .A3(n_1400), .B1(n_1403), .B2(n_1408), .B3(n_1411), .Y(n_1398) );
OAI33xp33_ASAP7_75t_L g1689 ( .A1(n_651), .A2(n_1411), .A3(n_1690), .B1(n_1694), .B2(n_1699), .B3(n_1702), .Y(n_1689) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g678 ( .A(n_655), .Y(n_678) );
BUFx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g769 ( .A(n_659), .Y(n_769) );
BUFx3_ASAP7_75t_L g932 ( .A(n_659), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_659), .B(n_1344), .Y(n_1343) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_669), .B2(n_670), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_663), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_663), .A2(n_675), .B1(n_928), .B2(n_929), .Y(n_927) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g753 ( .A(n_666), .Y(n_753) );
INVx2_ASAP7_75t_SL g1404 ( .A(n_666), .Y(n_1404) );
INVx2_ASAP7_75t_L g1695 ( .A(n_666), .Y(n_1695) );
BUFx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g838 ( .A(n_667), .Y(n_838) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g760 ( .A(n_668), .Y(n_760) );
INVx1_ASAP7_75t_L g825 ( .A(n_668), .Y(n_825) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_672), .A2(n_824), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_674), .A2(n_687), .B1(n_689), .B2(n_695), .C(n_697), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_675), .A2(n_823), .B1(n_826), .B2(n_827), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_676), .A2(n_679), .B1(n_719), .B2(n_722), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_678), .A2(n_924), .B1(n_925), .B2(n_926), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_680), .A2(n_850), .B1(n_943), .B2(n_944), .C(n_976), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_681), .A2(n_704), .B1(n_711), .B2(n_713), .C(n_715), .Y(n_703) );
OAI33xp33_ASAP7_75t_L g920 ( .A1(n_682), .A2(n_921), .A3(n_923), .B1(n_927), .B2(n_930), .B3(n_931), .Y(n_920) );
CKINVDCx8_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g1180 ( .A(n_683), .B(n_1181), .C(n_1186), .Y(n_1180) );
NAND3xp33_ASAP7_75t_L g1293 ( .A(n_683), .B(n_1294), .C(n_1296), .Y(n_1293) );
NAND3xp33_ASAP7_75t_L g1739 ( .A(n_683), .B(n_1740), .C(n_1741), .Y(n_1739) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_703), .C(n_718), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_687), .A2(n_761), .B1(n_774), .B2(n_780), .C(n_785), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_687), .A2(n_893), .B1(n_894), .B2(n_897), .C(n_898), .Y(n_892) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx4_ASAP7_75t_L g870 ( .A(n_691), .Y(n_870) );
INVx2_ASAP7_75t_L g1194 ( .A(n_691), .Y(n_1194) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
BUFx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_L g901 ( .A(n_706), .Y(n_901) );
INVx1_ASAP7_75t_L g962 ( .A(n_706), .Y(n_962) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_713), .A2(n_715), .B1(n_770), .B2(n_788), .C(n_793), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_713), .A2(n_715), .B1(n_900), .B2(n_904), .C(n_906), .Y(n_899) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g1652 ( .A(n_714), .Y(n_1652) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_719), .A2(n_722), .B1(n_765), .B2(n_767), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_719), .A2(n_722), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g1647 ( .A1(n_719), .A2(n_722), .B1(n_1648), .B2(n_1649), .Y(n_1647) );
INVx6_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g942 ( .A(n_721), .Y(n_942) );
INVx2_ASAP7_75t_L g954 ( .A(n_721), .Y(n_954) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_721), .B(n_1222), .Y(n_1221) );
INVx4_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g784 ( .A(n_724), .Y(n_784) );
INVx1_ASAP7_75t_L g1385 ( .A(n_724), .Y(n_1385) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_726), .A2(n_889), .B1(n_891), .B2(n_910), .Y(n_888) );
INVx5_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g1674 ( .A(n_727), .Y(n_1674) );
AND2x4_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g799 ( .A(n_730), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_771), .Y(n_731) );
NOR3xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_741), .C(n_743), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_738), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_749), .B2(n_750), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_746), .A2(n_767), .B1(n_768), .B2(n_770), .Y(n_766) );
OAI22xp33_ASAP7_75t_L g931 ( .A1(n_746), .A2(n_906), .B1(n_908), .B2(n_932), .Y(n_931) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp33_ASAP7_75t_L g1690 ( .A1(n_747), .A2(n_1691), .B1(n_1692), .B2(n_1693), .Y(n_1690) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_755), .A2(n_971), .B1(n_973), .B2(n_974), .Y(n_970) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_761), .B1(n_762), .B2(n_765), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_760), .B(n_1360), .Y(n_1359) );
INVx2_ASAP7_75t_L g1402 ( .A(n_760), .Y(n_1402) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g841 ( .A(n_764), .Y(n_841) );
INVx2_ASAP7_75t_L g1295 ( .A(n_764), .Y(n_1295) );
INVx2_ASAP7_75t_SL g1406 ( .A(n_764), .Y(n_1406) );
OAI22xp33_ASAP7_75t_L g1408 ( .A1(n_768), .A2(n_819), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g815 ( .A(n_769), .Y(n_815) );
INVx1_ASAP7_75t_L g925 ( .A(n_769), .Y(n_925) );
NAND3xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_787), .C(n_797), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_783), .Y(n_896) );
BUFx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g863 ( .A(n_784), .Y(n_863) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g895 ( .A(n_790), .Y(n_895) );
INVx1_ASAP7_75t_L g1241 ( .A(n_790), .Y(n_1241) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g1242 ( .A(n_796), .Y(n_1242) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
XNOR2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_933), .Y(n_803) );
AOI22x1_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_884), .B2(n_885), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_852), .C(n_854), .Y(n_807) );
OAI221xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_817), .B2(n_820), .C(n_821), .Y(n_814) );
OAI221xp5_ASAP7_75t_L g1032 ( .A1(n_817), .A2(n_850), .B1(n_1009), .B2(n_1010), .C(n_1033), .Y(n_1032) );
OAI221xp5_ASAP7_75t_L g1098 ( .A1(n_817), .A2(n_850), .B1(n_1099), .B2(n_1100), .C(n_1101), .Y(n_1098) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g848 ( .A(n_819), .Y(n_848) );
BUFx2_ASAP7_75t_L g976 ( .A(n_819), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_819), .A2(n_844), .B1(n_1387), .B2(n_1389), .Y(n_1399) );
OAI22xp33_ASAP7_75t_L g1702 ( .A1(n_819), .A2(n_932), .B1(n_1648), .B2(n_1653), .Y(n_1702) );
BUFx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_824), .A2(n_1185), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g1089 ( .A(n_825), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1701 ( .A(n_825), .Y(n_1701) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .B1(n_832), .B2(n_833), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_830), .A2(n_833), .B1(n_990), .B2(n_991), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_830), .A2(n_833), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_830), .A2(n_833), .B1(n_1071), .B2(n_1072), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_839), .B1(n_840), .B2(n_842), .Y(n_836) );
BUFx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g972 ( .A(n_838), .Y(n_972) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_846), .B1(n_847), .B2(n_849), .C(n_850), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g1692 ( .A(n_845), .Y(n_1692) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NOR2xp33_ASAP7_75t_SL g854 ( .A(n_855), .B(n_881), .Y(n_854) );
NAND3xp33_ASAP7_75t_SL g855 ( .A(n_856), .B(n_858), .C(n_878), .Y(n_855) );
AOI33xp33_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .A3(n_864), .B1(n_869), .B2(n_871), .B3(n_876), .Y(n_858) );
INVx2_ASAP7_75t_SL g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g1077 ( .A(n_863), .Y(n_1077) );
INVx1_ASAP7_75t_L g1082 ( .A(n_863), .Y(n_1082) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g1079 ( .A(n_868), .Y(n_1079) );
INVx2_ASAP7_75t_L g1156 ( .A(n_868), .Y(n_1156) );
INVx1_ASAP7_75t_L g1382 ( .A(n_872), .Y(n_1382) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NAND3xp33_ASAP7_75t_L g1751 ( .A(n_876), .B(n_1752), .C(n_1753), .Y(n_1751) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NAND3xp33_ASAP7_75t_L g1069 ( .A(n_878), .B(n_1070), .C(n_1073), .Y(n_1069) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
INVx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
XNOR2x1_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
AND2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_911), .Y(n_887) );
INVx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
BUFx8_ASAP7_75t_SL g1346 ( .A(n_890), .Y(n_1346) );
NAND3xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_899), .C(n_907), .Y(n_891) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR3xp33_ASAP7_75t_SL g911 ( .A(n_912), .B(n_919), .C(n_920), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_916), .Y(n_912) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
XOR2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_1001), .Y(n_933) );
AND4x1_ASAP7_75t_L g935 ( .A(n_936), .B(n_965), .C(n_967), .D(n_993), .Y(n_935) );
NOR3xp33_ASAP7_75t_SL g936 ( .A(n_937), .B(n_938), .C(n_963), .Y(n_936) );
NOR3xp33_ASAP7_75t_SL g1006 ( .A(n_937), .B(n_1007), .C(n_1023), .Y(n_1006) );
OAI221xp5_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_943), .B1(n_944), .B2(n_945), .C(n_948), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_940), .A2(n_945), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1008) );
BUFx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
BUFx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1016 ( .A(n_947), .Y(n_1016) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
OAI33xp33_ASAP7_75t_L g1379 ( .A1(n_951), .A2(n_1315), .A3(n_1380), .B1(n_1386), .B2(n_1391), .B3(n_1394), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_955), .B1(n_956), .B2(n_959), .C(n_960), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g1014 ( .A1(n_953), .A2(n_1015), .B1(n_1016), .B2(n_1017), .C(n_1018), .Y(n_1014) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g998 ( .A(n_954), .Y(n_998) );
INVx2_ASAP7_75t_L g1388 ( .A(n_954), .Y(n_1388) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
BUFx2_ASAP7_75t_L g1390 ( .A(n_958), .Y(n_1390) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
OAI31xp33_ASAP7_75t_SL g967 ( .A1(n_968), .A2(n_969), .A3(n_977), .B(n_992), .Y(n_967) );
INVx2_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx2_ASAP7_75t_L g979 ( .A(n_972), .Y(n_979) );
OAI221xp5_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_980), .B1(n_981), .B2(n_984), .C(n_985), .Y(n_978) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_979), .A2(n_1041), .B1(n_1042), .B2(n_1045), .C(n_1046), .Y(n_1040) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g1699 ( .A1(n_983), .A2(n_1649), .B1(n_1662), .B2(n_1700), .Y(n_1699) );
CKINVDCx8_ASAP7_75t_R g1107 ( .A(n_992), .Y(n_1107) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_994), .B(n_996), .Y(n_993) );
XNOR2xp5_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
AND4x1_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1006), .C(n_1027), .D(n_1050), .Y(n_1003) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_1013), .Y(n_1012) );
BUFx3_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1022), .Y(n_1154) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1034), .Y(n_1099) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1044), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_1044), .A2(n_1381), .B1(n_1383), .B2(n_1401), .Y(n_1400) );
NOR2xp33_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_1054), .Y(n_1053) );
XNOR2xp5_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1250), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
XOR2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1108), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
NAND3xp33_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1083), .C(n_1085), .Y(n_1060) );
NOR2xp33_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1069), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1066), .Y(n_1062) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_1064), .A2(n_1068), .B1(n_1088), .B2(n_1090), .C(n_1092), .Y(n_1087) );
OAI31xp33_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1097), .A3(n_1105), .B(n_1106), .Y(n_1085) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
A2O1A1Ixp33_ASAP7_75t_L g1341 ( .A1(n_1094), .A2(n_1342), .B(n_1343), .C(n_1345), .Y(n_1341) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1095), .Y(n_1364) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1645 ( .A1(n_1107), .A2(n_1646), .B1(n_1673), .B2(n_1674), .Y(n_1645) );
XNOR2xp5_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1160), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AOI211x1_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1126), .B(n_1127), .C(n_1143), .Y(n_1111) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
AOI221x1_ASAP7_75t_L g1255 ( .A1(n_1126), .A2(n_1256), .B1(n_1269), .B2(n_1286), .C(n_1287), .Y(n_1255) );
AOI221x1_ASAP7_75t_L g1713 ( .A1(n_1126), .A2(n_1286), .B1(n_1714), .B2(n_1727), .C(n_1738), .Y(n_1713) );
AOI31xp33_ASAP7_75t_L g1127 ( .A1(n_1128), .A2(n_1135), .A3(n_1139), .B(n_1142), .Y(n_1127) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_SL g1130 ( .A(n_1131), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_1131), .Y(n_1191) );
AOI31xp33_ASAP7_75t_L g1197 ( .A1(n_1142), .A2(n_1198), .A3(n_1202), .B(n_1205), .Y(n_1197) );
AO21x1_ASAP7_75t_SL g1225 ( .A1(n_1142), .A2(n_1226), .B(n_1230), .Y(n_1225) );
CKINVDCx16_ASAP7_75t_R g1286 ( .A(n_1142), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1152), .Y(n_1143) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
AOI222xp33_ASAP7_75t_L g1731 ( .A1(n_1151), .A2(n_1276), .B1(n_1732), .B2(n_1733), .C1(n_1734), .C2(n_1735), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1156), .B(n_1212), .Y(n_1211) );
XNOR2x1_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1207), .Y(n_1160) );
NAND3xp33_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1169), .C(n_1172), .Y(n_1163) );
NAND4xp25_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1180), .C(n_1187), .D(n_1192), .Y(n_1175) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1201), .Y(n_1734) );
AND4x1_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1225), .C(n_1233), .D(n_1239), .Y(n_1208) );
NAND4xp25_ASAP7_75t_L g1249 ( .A(n_1209), .B(n_1225), .C(n_1233), .D(n_1239), .Y(n_1249) );
OAI31xp33_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1217), .A3(n_1220), .B(n_1224), .Y(n_1209) );
NAND3xp33_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1213), .C(n_1216), .Y(n_1210) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1222), .Y(n_1375) );
OAI31xp33_ASAP7_75t_SL g1368 ( .A1(n_1224), .A2(n_1369), .A3(n_1370), .B(n_1371), .Y(n_1368) );
NAND3xp33_ASAP7_75t_L g1288 ( .A(n_1234), .B(n_1289), .C(n_1292), .Y(n_1288) );
NAND3xp33_ASAP7_75t_L g1744 ( .A(n_1234), .B(n_1745), .C(n_1747), .Y(n_1744) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1252), .B1(n_1352), .B2(n_1353), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
XOR2xp5_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1307), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1255), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1260), .Y(n_1256) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx2_ASAP7_75t_L g1717 ( .A(n_1265), .Y(n_1717) );
NAND4xp25_ASAP7_75t_SL g1269 ( .A(n_1270), .B(n_1273), .C(n_1283), .D(n_1285), .Y(n_1269) );
AND2x4_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NAND4xp25_ASAP7_75t_SL g1727 ( .A(n_1285), .B(n_1728), .C(n_1731), .D(n_1736), .Y(n_1727) );
NAND4xp25_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1293), .C(n_1297), .D(n_1301), .Y(n_1287) );
INVx2_ASAP7_75t_SL g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx2_ASAP7_75t_SL g1308 ( .A(n_1309), .Y(n_1308) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NAND4xp75_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1326), .C(n_1347), .D(n_1349), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1323), .Y(n_1312) );
INVx1_ASAP7_75t_SL g1314 ( .A(n_1315), .Y(n_1314) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
OAI21xp5_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1336), .B(n_1346), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1331), .Y(n_1327) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
HB1xp67_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1355), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g1391 ( .A1(n_1357), .A2(n_1388), .B1(n_1392), .B2(n_1393), .Y(n_1391) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g1403 ( .A1(n_1376), .A2(n_1404), .B1(n_1405), .B2(n_1407), .Y(n_1403) );
NOR2xp33_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1398), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_1381), .A2(n_1382), .B1(n_1383), .B2(n_1384), .Y(n_1380) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
OAI22xp33_ASAP7_75t_SL g1386 ( .A1(n_1387), .A2(n_1388), .B1(n_1389), .B2(n_1390), .Y(n_1386) );
INVx2_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
OAI221xp5_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1425), .B1(n_1641), .B2(n_1704), .C(n_1709), .Y(n_1414) );
CKINVDCx16_ASAP7_75t_R g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
OAI22xp33_ASAP7_75t_L g1515 ( .A1(n_1417), .A2(n_1516), .B1(n_1517), .B2(n_1518), .Y(n_1515) );
BUFx3_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
OAI22xp5_ASAP7_75t_L g1440 ( .A1(n_1418), .A2(n_1441), .B1(n_1442), .B2(n_1443), .Y(n_1440) );
OAI22xp33_ASAP7_75t_L g1459 ( .A1(n_1418), .A2(n_1443), .B1(n_1460), .B2(n_1461), .Y(n_1459) );
OAI22xp33_ASAP7_75t_L g1468 ( .A1(n_1418), .A2(n_1469), .B1(n_1470), .B2(n_1471), .Y(n_1468) );
BUFx6f_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1421), .Y(n_1419) );
OR2x2_ASAP7_75t_L g1443 ( .A(n_1420), .B(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1420), .Y(n_1450) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1421), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1424), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1424), .Y(n_1437) );
NOR3xp33_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1602), .C(n_1624), .Y(n_1425) );
AOI22xp5_ASAP7_75t_L g1426 ( .A1(n_1427), .A2(n_1498), .B1(n_1564), .B2(n_1576), .Y(n_1426) );
AOI311xp33_ASAP7_75t_L g1427 ( .A1(n_1428), .A2(n_1462), .A3(n_1477), .B(n_1480), .C(n_1493), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1454), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1430), .B(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
OAI22xp33_ASAP7_75t_L g1500 ( .A1(n_1431), .A2(n_1473), .B1(n_1501), .B2(n_1504), .Y(n_1500) );
NOR2xp33_ASAP7_75t_L g1582 ( .A(n_1431), .B(n_1532), .Y(n_1582) );
OAI21xp33_ASAP7_75t_SL g1589 ( .A1(n_1431), .A2(n_1531), .B(n_1590), .Y(n_1589) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1445), .Y(n_1431) );
INVx2_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1433), .B(n_1458), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1433), .B(n_1445), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1433), .B(n_1484), .Y(n_1526) );
NOR2xp33_ASAP7_75t_L g1558 ( .A(n_1433), .B(n_1445), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1433), .B(n_1508), .Y(n_1595) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1434), .B(n_1484), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1434), .B(n_1458), .Y(n_1541) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1435), .Y(n_1514) );
AND2x4_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1438), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1436), .B(n_1438), .Y(n_1475) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_1437), .B(n_1438), .Y(n_1439) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1439), .Y(n_1467) );
HB1xp67_ASAP7_75t_L g1471 ( .A(n_1443), .Y(n_1471) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1443), .Y(n_1519) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1444), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1445), .B(n_1456), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1445), .B(n_1477), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1445), .B(n_1507), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1445), .B(n_1587), .Y(n_1622) );
BUFx3_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1446), .B(n_1483), .Y(n_1494) );
INVx2_ASAP7_75t_L g1508 ( .A(n_1446), .Y(n_1508) );
OR2x2_ASAP7_75t_L g1528 ( .A(n_1446), .B(n_1529), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1446), .B(n_1526), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1446), .B(n_1541), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1446), .B(n_1457), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1446), .B(n_1507), .Y(n_1607) );
O2A1O1Ixp33_ASAP7_75t_L g1616 ( .A1(n_1446), .A2(n_1617), .B(n_1621), .C(n_1623), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1453), .Y(n_1446) );
AND2x4_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1450), .Y(n_1448) );
OAI21xp33_ASAP7_75t_SL g1759 ( .A1(n_1449), .A2(n_1757), .B(n_1760), .Y(n_1759) );
AND2x4_ASAP7_75t_L g1451 ( .A(n_1450), .B(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
AOI21xp5_ASAP7_75t_L g1527 ( .A1(n_1456), .A2(n_1528), .B(n_1530), .Y(n_1527) );
AOI32xp33_ASAP7_75t_L g1580 ( .A1(n_1456), .A2(n_1481), .A3(n_1534), .B1(n_1581), .B2(n_1582), .Y(n_1580) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_1457), .B(n_1532), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1457), .B(n_1485), .Y(n_1606) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1458), .Y(n_1484) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1458), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_1462), .B(n_1544), .Y(n_1543) );
AOI22xp33_ASAP7_75t_SL g1605 ( .A1(n_1462), .A2(n_1562), .B1(n_1606), .B2(n_1607), .Y(n_1605) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1472), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1464), .B(n_1473), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_1464), .B(n_1538), .Y(n_1599) );
AND2x4_ASAP7_75t_SL g1615 ( .A(n_1464), .B(n_1472), .Y(n_1615) );
INVx2_ASAP7_75t_SL g1464 ( .A(n_1465), .Y(n_1464) );
INVx2_ASAP7_75t_L g1496 ( .A(n_1465), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1537 ( .A(n_1465), .B(n_1538), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1465), .B(n_1472), .Y(n_1640) );
INVx2_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_1472), .B(n_1487), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_1472), .B(n_1490), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1472), .B(n_1534), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1472), .B(n_1573), .Y(n_1596) );
CKINVDCx6p67_ASAP7_75t_R g1472 ( .A(n_1473), .Y(n_1472) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_1473), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1473), .B(n_1490), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1473), .B(n_1524), .Y(n_1523) );
AOI221xp5_ASAP7_75t_L g1631 ( .A1(n_1473), .A2(n_1566), .B1(n_1632), .B2(n_1636), .C(n_1637), .Y(n_1631) );
OR2x6_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1476), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1477), .B(n_1490), .Y(n_1489) );
INVx4_ASAP7_75t_L g1502 ( .A(n_1477), .Y(n_1502) );
INVx3_ASAP7_75t_L g1532 ( .A(n_1477), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1477), .B(n_1526), .Y(n_1590) );
NOR2xp67_ASAP7_75t_SL g1612 ( .A(n_1477), .B(n_1488), .Y(n_1612) );
OR2x2_ASAP7_75t_L g1628 ( .A(n_1477), .B(n_1490), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1636 ( .A(n_1477), .B(n_1523), .Y(n_1636) );
AND2x4_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1479), .Y(n_1477) );
OAI21xp33_ASAP7_75t_L g1480 ( .A1(n_1481), .A2(n_1482), .B(n_1486), .Y(n_1480) );
A2O1A1Ixp33_ASAP7_75t_L g1571 ( .A1(n_1481), .A2(n_1538), .B(n_1572), .C(n_1574), .Y(n_1571) );
OAI211xp5_ASAP7_75t_SL g1577 ( .A1(n_1482), .A2(n_1522), .B(n_1578), .C(n_1580), .Y(n_1577) );
OR2x2_ASAP7_75t_L g1625 ( .A(n_1482), .B(n_1538), .Y(n_1625) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1482), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1485), .Y(n_1482) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1483), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1483), .B(n_1502), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1483), .B(n_1581), .Y(n_1604) );
INVxp67_ASAP7_75t_L g1638 ( .A(n_1487), .Y(n_1638) );
NOR2xp33_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1489), .Y(n_1487) );
INVx1_ASAP7_75t_SL g1524 ( .A(n_1490), .Y(n_1524) );
CKINVDCx5p33_ASAP7_75t_R g1534 ( .A(n_1490), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1490), .B(n_1502), .Y(n_1549) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1490), .Y(n_1563) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1490), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1603 ( .A(n_1490), .B(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1490), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1492), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1495), .Y(n_1493) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1494), .Y(n_1600) );
OAI21xp33_ASAP7_75t_L g1565 ( .A1(n_1495), .A2(n_1566), .B(n_1567), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1497), .Y(n_1495) );
INVx2_ASAP7_75t_L g1509 ( .A(n_1496), .Y(n_1509) );
INVx2_ASAP7_75t_L g1553 ( .A(n_1496), .Y(n_1553) );
OAI211xp5_ASAP7_75t_SL g1624 ( .A1(n_1496), .A2(n_1625), .B(n_1626), .C(n_1631), .Y(n_1624) );
NOR2xp33_ASAP7_75t_L g1627 ( .A(n_1496), .B(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1497), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1499), .B(n_1535), .Y(n_1498) );
AOI211xp5_ASAP7_75t_L g1499 ( .A1(n_1500), .A2(n_1509), .B(n_1510), .C(n_1527), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1502), .B(n_1503), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1502), .B(n_1506), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1502), .B(n_1540), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1502), .B(n_1523), .Y(n_1570) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1502), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1502), .B(n_1508), .Y(n_1581) );
AOI22xp5_ASAP7_75t_L g1594 ( .A1(n_1503), .A2(n_1506), .B1(n_1595), .B2(n_1596), .Y(n_1594) );
AOI31xp33_ASAP7_75t_L g1610 ( .A1(n_1504), .A2(n_1528), .A3(n_1588), .B(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
NOR2x1_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1508), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1508), .B(n_1526), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1508), .B(n_1541), .Y(n_1540) );
OR2x2_ASAP7_75t_L g1575 ( .A(n_1508), .B(n_1555), .Y(n_1575) );
NAND2xp5_ASAP7_75t_L g1550 ( .A(n_1509), .B(n_1551), .Y(n_1550) );
OAI21xp33_ASAP7_75t_L g1556 ( .A1(n_1509), .A2(n_1557), .B(n_1559), .Y(n_1556) );
AOI211xp5_ASAP7_75t_L g1576 ( .A1(n_1509), .A2(n_1577), .B(n_1583), .C(n_1593), .Y(n_1576) );
OAI221xp5_ASAP7_75t_L g1602 ( .A1(n_1509), .A2(n_1603), .B1(n_1605), .B2(n_1608), .C(n_1609), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1520), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
BUFx3_ASAP7_75t_L g1592 ( .A(n_1512), .Y(n_1592) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_1522), .B(n_1525), .Y(n_1521) );
OAI21xp33_ASAP7_75t_L g1583 ( .A1(n_1522), .A2(n_1584), .B(n_1586), .Y(n_1583) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1525), .Y(n_1566) );
OR2x2_ASAP7_75t_L g1614 ( .A(n_1525), .B(n_1532), .Y(n_1614) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1526), .Y(n_1619) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1528), .B(n_1630), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1533), .Y(n_1530) );
OR2x2_ASAP7_75t_L g1578 ( .A(n_1531), .B(n_1579), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1531), .B(n_1540), .Y(n_1585) );
INVx2_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1532), .B(n_1546), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1567 ( .A(n_1532), .B(n_1558), .Y(n_1567) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1533), .Y(n_1601) );
INVx3_ASAP7_75t_L g1538 ( .A(n_1534), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1534), .B(n_1615), .Y(n_1623) );
AOI211xp5_ASAP7_75t_SL g1535 ( .A1(n_1536), .A2(n_1539), .B(n_1542), .C(n_1547), .Y(n_1535) );
AOI221xp5_ASAP7_75t_L g1586 ( .A1(n_1536), .A2(n_1587), .B1(n_1588), .B2(n_1589), .C(n_1591), .Y(n_1586) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1541), .Y(n_1620) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1546), .Y(n_1630) );
OAI21xp5_ASAP7_75t_SL g1547 ( .A1(n_1548), .A2(n_1550), .B(n_1552), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
OAI211xp5_ASAP7_75t_L g1552 ( .A1(n_1553), .A2(n_1554), .B(n_1556), .C(n_1560), .Y(n_1552) );
OAI222xp33_ASAP7_75t_L g1593 ( .A1(n_1553), .A2(n_1594), .B1(n_1597), .B2(n_1599), .C1(n_1600), .C2(n_1601), .Y(n_1593) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVxp33_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1558), .B(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1563), .Y(n_1561) );
AND3x1_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1568), .C(n_1571), .Y(n_1564) );
OAI21xp33_ASAP7_75t_L g1626 ( .A1(n_1569), .A2(n_1627), .B(n_1629), .Y(n_1626) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1588), .Y(n_1608) );
INVx2_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
AOI21xp5_ASAP7_75t_L g1637 ( .A1(n_1597), .A2(n_1638), .B(n_1639), .Y(n_1637) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
O2A1O1Ixp33_ASAP7_75t_L g1609 ( .A1(n_1610), .A2(n_1613), .B(n_1615), .C(n_1616), .Y(n_1609) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1620), .Y(n_1618) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1633), .B(n_1635), .Y(n_1632) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
HB1xp67_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1644), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1645), .B(n_1675), .Y(n_1644) );
NAND3xp33_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1650), .C(n_1660), .Y(n_1646) );
AOI221xp5_ASAP7_75t_L g1650 ( .A1(n_1651), .A2(n_1653), .B1(n_1654), .B2(n_1657), .C(n_1658), .Y(n_1650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
INVx3_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
AOI221xp5_ASAP7_75t_L g1660 ( .A1(n_1661), .A2(n_1662), .B1(n_1663), .B2(n_1664), .C(n_1668), .Y(n_1660) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_SL g1669 ( .A(n_1670), .Y(n_1669) );
INVx2_ASAP7_75t_SL g1671 ( .A(n_1672), .Y(n_1671) );
NOR3xp33_ASAP7_75t_L g1675 ( .A(n_1676), .B(n_1686), .C(n_1689), .Y(n_1675) );
NAND2xp5_ASAP7_75t_SL g1676 ( .A(n_1677), .B(n_1682), .Y(n_1676) );
AOI22xp33_ASAP7_75t_L g1677 ( .A1(n_1678), .A2(n_1679), .B1(n_1680), .B2(n_1681), .Y(n_1677) );
OAI22xp5_ASAP7_75t_L g1694 ( .A1(n_1695), .A2(n_1696), .B1(n_1697), .B2(n_1698), .Y(n_1694) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1697), .Y(n_1746) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
CKINVDCx5p33_ASAP7_75t_R g1704 ( .A(n_1705), .Y(n_1704) );
BUFx2_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVxp33_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
HB1xp67_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
NAND3xp33_ASAP7_75t_L g1714 ( .A(n_1715), .B(n_1721), .C(n_1724), .Y(n_1714) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
NAND4xp25_ASAP7_75t_L g1738 ( .A(n_1739), .B(n_1744), .C(n_1748), .D(n_1751), .Y(n_1738) );
INVx2_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
CKINVDCx5p33_ASAP7_75t_R g1755 ( .A(n_1756), .Y(n_1755) );
HB1xp67_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
endmodule