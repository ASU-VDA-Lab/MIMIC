module fake_jpeg_20121_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_45),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_14),
.Y(n_45)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_40),
.C(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_60),
.B1(n_22),
.B2(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_53),
.Y(n_77)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_55),
.Y(n_95)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_68),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_25),
.B1(n_19),
.B2(n_44),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_65),
.B1(n_78),
.B2(n_86),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_25),
.B1(n_44),
.B2(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_69),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_74),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_45),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_81),
.C(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_31),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_21),
.B1(n_19),
.B2(n_31),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_16),
.B1(n_21),
.B2(n_43),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_43),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_95),
.B1(n_68),
.B2(n_76),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_38),
.B(n_1),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_94),
.B(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_62),
.B1(n_57),
.B2(n_52),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_56),
.B1(n_55),
.B2(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_20),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_97),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_62),
.B1(n_57),
.B2(n_52),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_116),
.B1(n_117),
.B2(n_86),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_115),
.B1(n_94),
.B2(n_95),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_21),
.B1(n_47),
.B2(n_56),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_78),
.B1(n_65),
.B2(n_70),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_63),
.A2(n_55),
.B1(n_16),
.B2(n_38),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_27),
.B1(n_24),
.B2(n_32),
.Y(n_117)
);

XNOR2x1_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_28),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_32),
.C(n_27),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_0),
.B(n_1),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_0),
.B(n_2),
.Y(n_152)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_75),
.A3(n_94),
.B1(n_89),
.B2(n_87),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_143),
.B(n_152),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_136),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_132),
.B1(n_148),
.B2(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_66),
.B1(n_73),
.B2(n_72),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_150),
.B1(n_153),
.B2(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_121),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_113),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_91),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_97),
.C(n_118),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_112),
.C(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_93),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_154),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_95),
.B1(n_92),
.B2(n_67),
.Y(n_146)
);

OAI22x1_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_112),
.B1(n_99),
.B2(n_120),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_67),
.B1(n_32),
.B2(n_27),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_30),
.B1(n_26),
.B2(n_14),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_30),
.B1(n_26),
.B2(n_88),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_88),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_112),
.A3(n_106),
.B1(n_99),
.B2(n_117),
.C1(n_122),
.C2(n_116),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_156),
.A2(n_20),
.A3(n_23),
.B1(n_33),
.B2(n_29),
.C1(n_18),
.C2(n_17),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_160),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_183),
.C(n_153),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_169),
.B(n_174),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_120),
.B1(n_125),
.B2(n_114),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_171),
.B1(n_54),
.B2(n_23),
.Y(n_204)
);

AOI22x1_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_103),
.B1(n_113),
.B2(n_23),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_173),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_120),
.B1(n_114),
.B2(n_110),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_110),
.B1(n_119),
.B2(n_88),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_140),
.B1(n_150),
.B2(n_137),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_69),
.B(n_2),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_130),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_186),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_162),
.B1(n_169),
.B2(n_168),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_185),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_139),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_54),
.C(n_29),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_136),
.B(n_28),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_29),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_28),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_28),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_135),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_205),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_195),
.B1(n_204),
.B2(n_163),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_132),
.B1(n_148),
.B2(n_151),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_160),
.B1(n_183),
.B2(n_178),
.Y(n_223)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_197),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_152),
.B1(n_139),
.B2(n_143),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_198),
.A2(n_164),
.B1(n_161),
.B2(n_159),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_200),
.B(n_213),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_207),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_175),
.C(n_187),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_28),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_29),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_33),
.B(n_20),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_155),
.B(n_180),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_219),
.B(n_3),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_172),
.B1(n_185),
.B2(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_29),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

BUFx4f_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

AOI22x1_ASAP7_75t_L g217 ( 
.A1(n_155),
.A2(n_20),
.B1(n_33),
.B2(n_29),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_0),
.B(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_237),
.B1(n_238),
.B2(n_201),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_223),
.B1(n_231),
.B2(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_225),
.C(n_235),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_165),
.C(n_18),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_13),
.B(n_4),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_18),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_202),
.C(n_205),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_18),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_243),
.Y(n_252)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_18),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_17),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_199),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_17),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_219),
.B(n_217),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_192),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_248),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_206),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_206),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_196),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_251),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_188),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_261),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_198),
.CI(n_212),
.CON(n_255),
.SN(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_262),
.B1(n_263),
.B2(n_220),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_199),
.C(n_188),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_239),
.C(n_227),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_191),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_207),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_223),
.B1(n_230),
.B2(n_193),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_281),
.B1(n_236),
.B2(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_221),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_241),
.C(n_224),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_224),
.C(n_231),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_244),
.C(n_242),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_283),
.C(n_261),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_236),
.B1(n_237),
.B2(n_217),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_197),
.C(n_228),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_249),
.C(n_250),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_292),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_297),
.Y(n_308)
);

OAI221xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_245),
.B1(n_254),
.B2(n_263),
.C(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_215),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_279),
.B1(n_275),
.B2(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_252),
.C(n_228),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_190),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_190),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_228),
.B(n_4),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_228),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_3),
.C(n_6),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_270),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_280),
.B1(n_267),
.B2(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_279),
.B1(n_292),
.B2(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_285),
.B(n_7),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_11),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_285),
.C(n_7),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_6),
.C(n_8),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_6),
.B(n_8),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_316),
.B1(n_300),
.B2(n_301),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_10),
.B1(n_11),
.B2(n_308),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_8),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_10),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_314),
.B(n_305),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_320),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_301),
.B(n_308),
.Y(n_323)
);

NAND2x1_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_324),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_328),
.B(n_326),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_313),
.B(n_325),
.C(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_316),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_10),
.B(n_11),
.Y(n_334)
);


endmodule