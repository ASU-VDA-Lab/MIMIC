module fake_jpeg_3498_n_591 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_591);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_591;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_60),
.B(n_61),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_0),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_65),
.B(n_72),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_29),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_74),
.Y(n_132)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_73),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_0),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_19),
.A2(n_20),
.B(n_58),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_76),
.A2(n_78),
.B(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g196 ( 
.A(n_77),
.B(n_79),
.Y(n_196)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_19),
.B(n_2),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_58),
.B1(n_46),
.B2(n_37),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_19),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_86),
.Y(n_141)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_85),
.B(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_20),
.B(n_3),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_R g88 ( 
.A(n_38),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_119),
.Y(n_147)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_92),
.B(n_100),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_20),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_93),
.A2(n_25),
.B1(n_42),
.B2(n_41),
.Y(n_186)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_106),
.B(n_40),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_43),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_115),
.Y(n_154)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_57),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_23),
.Y(n_118)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_43),
.B(n_3),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_5),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_32),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_63),
.A2(n_55),
.B1(n_57),
.B2(n_56),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_126),
.A2(n_143),
.B1(n_159),
.B2(n_169),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_128),
.B(n_193),
.Y(n_265)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_77),
.A2(n_55),
.B1(n_37),
.B2(n_58),
.Y(n_143)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_79),
.A2(n_55),
.B1(n_46),
.B2(n_25),
.Y(n_159)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_163),
.Y(n_252)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_93),
.A2(n_51),
.B1(n_55),
.B2(n_46),
.Y(n_166)
);

OA22x2_ASAP7_75t_SL g244 ( 
.A1(n_166),
.A2(n_54),
.B1(n_49),
.B2(n_8),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_113),
.A2(n_34),
.B1(n_52),
.B2(n_48),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_86),
.A2(n_34),
.B1(n_52),
.B2(n_48),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_172),
.A2(n_186),
.B1(n_187),
.B2(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_174),
.B(n_179),
.Y(n_224)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_175),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_32),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_176),
.B(n_182),
.Y(n_236)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_88),
.B(n_56),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_105),
.A2(n_30),
.B1(n_45),
.B2(n_44),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_181),
.A2(n_185),
.B1(n_195),
.B2(n_75),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_30),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_111),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_70),
.A2(n_27),
.B1(n_42),
.B2(n_41),
.Y(n_187)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_81),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_191),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_109),
.A2(n_40),
.B1(n_35),
.B2(n_54),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_67),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_197),
.Y(n_249)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_71),
.A2(n_98),
.B1(n_90),
.B2(n_104),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_202),
.B(n_220),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_141),
.B(n_64),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_203),
.B(n_204),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_91),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_112),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_205),
.B(n_213),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_206),
.Y(n_284)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_208),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_169),
.A2(n_121),
.B1(n_96),
.B2(n_103),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_210),
.A2(n_215),
.B1(n_217),
.B2(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_82),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_212),
.B(n_241),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_147),
.B(n_35),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_127),
.B(n_99),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_214),
.B(n_242),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_118),
.B1(n_107),
.B2(n_117),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_124),
.A2(n_83),
.B(n_73),
.C(n_110),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_217),
.A2(n_10),
.B(n_14),
.C(n_15),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_218),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_164),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_222),
.B(n_243),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g318 ( 
.A1(n_223),
.A2(n_244),
.B1(n_239),
.B2(n_226),
.Y(n_318)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_110),
.B(n_118),
.C(n_107),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_229),
.A2(n_184),
.B(n_138),
.Y(n_286)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_232),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_128),
.A2(n_38),
.B1(n_54),
.B2(n_39),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_235),
.A2(n_247),
.B(n_249),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_192),
.A2(n_54),
.B1(n_49),
.B2(n_38),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_166),
.A2(n_54),
.B1(n_38),
.B2(n_49),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_238),
.A2(n_213),
.B1(n_233),
.B2(n_208),
.Y(n_309)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_162),
.Y(n_239)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_239),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_132),
.B(n_5),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_6),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_173),
.B(n_6),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_167),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_248),
.B(n_257),
.Y(n_308)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

INVx11_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_156),
.Y(n_251)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_123),
.Y(n_253)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_255),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_183),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_256),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_150),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_150),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_264),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_155),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_266),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_125),
.B(n_6),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_271),
.C(n_157),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_7),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_261),
.B(n_262),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_134),
.B(n_7),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_133),
.B(n_8),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_158),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_135),
.B(n_9),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_269),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_184),
.Y(n_270)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_270),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_137),
.B(n_10),
.C(n_11),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_195),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_272),
.A2(n_130),
.B1(n_142),
.B2(n_10),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_265),
.A2(n_185),
.B1(n_181),
.B2(n_159),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_274),
.A2(n_282),
.B1(n_287),
.B2(n_309),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_276),
.B(n_286),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_143),
.B(n_198),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_278),
.A2(n_281),
.B(n_311),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_153),
.B(n_157),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_235),
.A2(n_170),
.B1(n_180),
.B2(n_144),
.Y(n_282)
);

NAND3xp33_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_300),
.C(n_314),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_233),
.A2(n_144),
.B1(n_129),
.B2(n_170),
.Y(n_287)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_204),
.A2(n_178),
.A3(n_158),
.B1(n_129),
.B2(n_180),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_298),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_203),
.B(n_178),
.C(n_130),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_304),
.C(n_328),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_292),
.A2(n_269),
.B(n_246),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_206),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_221),
.A2(n_14),
.B1(n_142),
.B2(n_244),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_301),
.A2(n_318),
.B1(n_305),
.B2(n_274),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_210),
.A2(n_215),
.B1(n_244),
.B2(n_205),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_302),
.A2(n_216),
.B1(n_219),
.B2(n_252),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_236),
.B(n_230),
.C(n_214),
.Y(n_304)
);

AO22x1_ASAP7_75t_SL g310 ( 
.A1(n_211),
.A2(n_209),
.B1(n_228),
.B2(n_245),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_254),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_263),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_321),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_234),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_242),
.A2(n_268),
.B(n_228),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_323),
.A2(n_331),
.B(n_320),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_231),
.B(n_273),
.C(n_260),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_209),
.Y(n_329)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_224),
.A2(n_260),
.B(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_255),
.Y(n_333)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_334),
.A2(n_336),
.B1(n_355),
.B2(n_379),
.Y(n_412)
);

AND2x2_ASAP7_75t_SL g335 ( 
.A(n_285),
.B(n_252),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_335),
.B(n_348),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_302),
.A2(n_246),
.B1(n_234),
.B2(n_219),
.Y(n_336)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_275),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_341),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_278),
.A2(n_259),
.B(n_240),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_342),
.A2(n_371),
.B(n_380),
.Y(n_408)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_249),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_344),
.B(n_360),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_285),
.B(n_216),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_346),
.B(n_351),
.C(n_352),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_347),
.A2(n_364),
.B(n_368),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_254),
.C(n_270),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_283),
.B(n_207),
.C(n_253),
.Y(n_352)
);

AND2x2_ASAP7_75t_SL g354 ( 
.A(n_322),
.B(n_250),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_276),
.A2(n_225),
.B1(n_251),
.B2(n_250),
.Y(n_355)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_358),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_322),
.B(n_227),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_372),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_295),
.B(n_232),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g362 ( 
.A(n_325),
.Y(n_362)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_275),
.Y(n_363)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_287),
.A2(n_218),
.B1(n_282),
.B2(n_323),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_365),
.A2(n_369),
.B1(n_373),
.B2(n_294),
.Y(n_389)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_279),
.Y(n_366)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_290),
.B(n_218),
.C(n_331),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_324),
.C(n_303),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_318),
.A2(n_286),
.B1(n_281),
.B2(n_305),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_277),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_311),
.A2(n_286),
.B(n_320),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_310),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_318),
.A2(n_292),
.B1(n_327),
.B2(n_277),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_293),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_376),
.Y(n_397)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_293),
.Y(n_375)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_333),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_308),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_297),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_289),
.B(n_296),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_378),
.B(n_332),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_318),
.A2(n_315),
.B1(n_299),
.B2(n_329),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_297),
.B(n_313),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_377),
.B(n_315),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_383),
.B(n_388),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_330),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_396),
.C(n_401),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_389),
.A2(n_400),
.B1(n_350),
.B2(n_336),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_393),
.B(n_402),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_330),
.Y(n_396)
);

AO22x2_ASAP7_75t_L g399 ( 
.A1(n_379),
.A2(n_299),
.B1(n_326),
.B2(n_291),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_414),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_338),
.A2(n_350),
.B1(n_369),
.B2(n_373),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_376),
.B(n_324),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_303),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_403),
.B(n_409),
.C(n_335),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_312),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_407),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_291),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_351),
.B(n_345),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_410),
.B(n_415),
.Y(n_420)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_411),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_356),
.A2(n_326),
.B(n_313),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_413),
.A2(n_365),
.B(n_354),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_374),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_359),
.B(n_312),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_380),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_418),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_346),
.B(n_307),
.Y(n_418)
);

A2O1A1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_414),
.A2(n_372),
.B(n_371),
.C(n_356),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_421),
.B(n_424),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_416),
.Y(n_422)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_422),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_397),
.A2(n_347),
.B(n_350),
.C(n_339),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_425),
.A2(n_427),
.B1(n_446),
.B2(n_450),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_419),
.A2(n_342),
.B(n_348),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_426),
.A2(n_429),
.B(n_445),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_338),
.B1(n_334),
.B2(n_355),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_352),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_431),
.C(n_437),
.Y(n_476)
);

XOR2x2_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_335),
.Y(n_430)
);

XOR2x1_ASAP7_75t_L g478 ( 
.A(n_430),
.B(n_404),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_387),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_408),
.Y(n_432)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_354),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_383),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_438),
.B(n_440),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_443),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_406),
.Y(n_441)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_409),
.B(n_375),
.C(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_419),
.A2(n_357),
.B(n_353),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_370),
.B1(n_366),
.B2(n_337),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_337),
.B(n_358),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_447),
.A2(n_453),
.B(n_395),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_397),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_418),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_385),
.A2(n_341),
.B1(n_363),
.B2(n_319),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_452),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_413),
.A2(n_307),
.B(n_319),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_442),
.Y(n_454)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_454),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_425),
.A2(n_385),
.B1(n_412),
.B2(n_416),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_456),
.A2(n_448),
.B1(n_446),
.B2(n_434),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_431),
.B(n_401),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_464),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g501 ( 
.A1(n_463),
.A2(n_450),
.B(n_451),
.Y(n_501)
);

XNOR2x1_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_416),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_420),
.B(n_381),
.C(n_395),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_467),
.B(n_420),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_468),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_428),
.B(n_417),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_474),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_426),
.A2(n_411),
.B(n_405),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_471),
.A2(n_429),
.B(n_447),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_433),
.B(n_412),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_399),
.B1(n_405),
.B2(n_404),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_475),
.A2(n_479),
.B1(n_482),
.B2(n_458),
.Y(n_504)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_477),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_480),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_421),
.A2(n_399),
.B1(n_392),
.B2(n_394),
.Y(n_479)
);

XOR2x2_ASAP7_75t_L g480 ( 
.A(n_433),
.B(n_399),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_439),
.B(n_399),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_443),
.C(n_430),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_438),
.A2(n_392),
.B1(n_394),
.B2(n_398),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_454),
.A2(n_449),
.B1(n_427),
.B2(n_432),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_483),
.A2(n_484),
.B1(n_500),
.B2(n_504),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_479),
.A2(n_459),
.B1(n_475),
.B2(n_468),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_485),
.B(n_497),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_486),
.B(n_503),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_430),
.C(n_422),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_494),
.C(n_498),
.Y(n_510)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_492),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_491),
.A2(n_501),
.B(n_462),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_481),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_468),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_499),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_448),
.C(n_424),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_495),
.A2(n_508),
.B1(n_471),
.B2(n_465),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_445),
.C(n_435),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_466),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_460),
.A2(n_453),
.B1(n_440),
.B2(n_444),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_456),
.B(n_434),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_507),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_463),
.Y(n_503)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_472),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_473),
.A2(n_423),
.B1(n_436),
.B2(n_452),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_512),
.B(n_519),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_514),
.B(n_518),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_474),
.C(n_455),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_517),
.Y(n_531)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_502),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g518 ( 
.A(n_494),
.B(n_478),
.CI(n_469),
.CON(n_518),
.SN(n_518)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_423),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_522),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_496),
.B(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_455),
.C(n_480),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_436),
.Y(n_523)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_461),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_524),
.B(n_526),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

BUFx12f_ASAP7_75t_SL g527 ( 
.A(n_491),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_527),
.A2(n_506),
.B(n_501),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_487),
.B(n_462),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_529),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_487),
.B(n_464),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_530),
.B(n_497),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_514),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_534),
.A2(n_528),
.B(n_521),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_522),
.C(n_515),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_538),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_510),
.B(n_505),
.C(n_488),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_516),
.B(n_507),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_539),
.B(n_513),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_505),
.C(n_506),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_529),
.C(n_513),
.Y(n_552)
);

OAI221xp5_ASAP7_75t_L g541 ( 
.A1(n_509),
.A2(n_499),
.B1(n_489),
.B2(n_484),
.C(n_500),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_541),
.A2(n_511),
.B1(n_523),
.B2(n_526),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_512),
.B(n_390),
.Y(n_543)
);

CKINVDCx14_ASAP7_75t_R g558 ( 
.A(n_543),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_509),
.B(n_390),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_525),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_512),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_551),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_549),
.B(n_552),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_535),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_554),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_533),
.C(n_540),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_534),
.B(n_518),
.Y(n_555)
);

NOR2x1_ASAP7_75t_L g569 ( 
.A(n_555),
.B(n_547),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_556),
.A2(n_560),
.B(n_536),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_542),
.A2(n_519),
.B1(n_524),
.B2(n_525),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_559),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_536),
.B(n_511),
.C(n_526),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_561),
.B(n_545),
.C(n_537),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_550),
.B(n_544),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_562),
.B(n_566),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_564),
.A2(n_569),
.B(n_549),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_547),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_567),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_554),
.B(n_537),
.C(n_546),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_568),
.B(n_571),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_392),
.Y(n_571)
);

NOR2x1p5_ASAP7_75t_L g573 ( 
.A(n_570),
.B(n_557),
.Y(n_573)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_573),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_565),
.B(n_559),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_577),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_563),
.B(n_561),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_579),
.B(n_555),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_574),
.B(n_568),
.C(n_567),
.Y(n_580)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_580),
.A2(n_583),
.B(n_584),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_576),
.B(n_572),
.C(n_569),
.Y(n_584)
);

O2A1O1Ixp33_ASAP7_75t_SL g585 ( 
.A1(n_581),
.A2(n_583),
.B(n_527),
.C(n_578),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_585),
.A2(n_586),
.B1(n_384),
.B2(n_284),
.Y(n_588)
);

O2A1O1Ixp33_ASAP7_75t_SL g586 ( 
.A1(n_582),
.A2(n_518),
.B(n_384),
.C(n_362),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_587),
.B(n_284),
.Y(n_589)
);

BUFx24_ASAP7_75t_SL g590 ( 
.A(n_589),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_343),
.Y(n_591)
);


endmodule