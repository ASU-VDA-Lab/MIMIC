module fake_jpeg_29598_n_394 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_394);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_394;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_42),
.Y(n_128)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_49),
.B(n_52),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_26),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_68),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_25),
.B(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_61),
.Y(n_119)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_18),
.B(n_0),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_38),
.C(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_13),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_63),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_67),
.Y(n_106)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_15),
.B(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_13),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_18),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_33),
.B(n_12),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_0),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_39),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_23),
.B1(n_30),
.B2(n_27),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_82),
.B(n_96),
.C(n_115),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_23),
.B1(n_30),
.B2(n_27),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_37),
.B1(n_34),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_83),
.A2(n_127),
.B1(n_56),
.B2(n_51),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_87),
.B(n_8),
.C(n_9),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_38),
.B(n_32),
.C(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_91),
.B(n_2),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_98),
.B(n_104),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_12),
.B(n_28),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_99),
.B(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_34),
.B1(n_37),
.B2(n_22),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_103),
.A2(n_126),
.B1(n_131),
.B2(n_79),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_22),
.Y(n_104)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_114),
.Y(n_159)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_47),
.B(n_19),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_21),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_17),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_73),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_21),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_57),
.A2(n_37),
.B1(n_17),
.B2(n_33),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_70),
.A2(n_33),
.B1(n_17),
.B2(n_5),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_43),
.A2(n_53),
.B1(n_66),
.B2(n_65),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_77),
.B1(n_75),
.B2(n_62),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_134),
.A2(n_138),
.B1(n_113),
.B2(n_133),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_146),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_63),
.B1(n_52),
.B2(n_48),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_145),
.Y(n_196)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_91),
.B1(n_121),
.B2(n_82),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_90),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_167),
.Y(n_189)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_81),
.A2(n_17),
.B1(n_79),
.B2(n_42),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_106),
.Y(n_153)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_49),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_165),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_79),
.B1(n_49),
.B2(n_42),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_161),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_169),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_96),
.A2(n_49),
.B1(n_42),
.B2(n_6),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_163),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_85),
.B(n_4),
.Y(n_164)
);

INVx6_ASAP7_75t_SL g166 ( 
.A(n_95),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_7),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_97),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_89),
.B(n_7),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_150),
.C(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_89),
.B(n_8),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_11),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_107),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_175),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_97),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_180),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_11),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_102),
.B(n_9),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_183),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_109),
.B(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_9),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_92),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_197),
.B1(n_214),
.B2(n_220),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_172),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_188),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_145),
.B(n_115),
.CI(n_128),
.CON(n_194),
.SN(n_194)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_194),
.B(n_215),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_92),
.B(n_130),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_152),
.B(n_181),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_113),
.B1(n_133),
.B2(n_122),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_101),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_101),
.Y(n_207)
);

AO22x1_ASAP7_75t_SL g208 ( 
.A1(n_148),
.A2(n_127),
.B1(n_83),
.B2(n_93),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_224),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_160),
.A2(n_95),
.B1(n_122),
.B2(n_130),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_93),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_139),
.A2(n_10),
.B1(n_168),
.B2(n_137),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_10),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_225),
.A2(n_251),
.B(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_154),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_228),
.B(n_229),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_232),
.B(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_159),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_235),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_167),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_239),
.Y(n_275)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_153),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_142),
.B1(n_139),
.B2(n_144),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_240),
.A2(n_246),
.B1(n_247),
.B2(n_218),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_139),
.B1(n_165),
.B2(n_155),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_205),
.B1(n_221),
.B2(n_214),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_165),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_243),
.B(n_245),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_140),
.C(n_158),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_248),
.C(n_255),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_165),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_196),
.A2(n_139),
.B1(n_166),
.B2(n_136),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_196),
.A2(n_139),
.B1(n_151),
.B2(n_143),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_170),
.C(n_183),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_195),
.B(n_212),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_193),
.B(n_147),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_254),
.Y(n_279)
);

AO22x1_ASAP7_75t_L g253 ( 
.A1(n_205),
.A2(n_147),
.B1(n_180),
.B2(n_176),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_200),
.B(n_141),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_141),
.C(n_135),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_178),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_135),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_205),
.A2(n_10),
.B(n_178),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_208),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_262),
.A2(n_278),
.B1(n_288),
.B2(n_210),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_269),
.B1(n_268),
.B2(n_241),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_204),
.C(n_207),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_271),
.C(n_282),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_184),
.A3(n_200),
.B1(n_215),
.B2(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_268),
.B(n_284),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_240),
.A2(n_247),
.B1(n_233),
.B2(n_246),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_191),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_277),
.B(n_188),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_208),
.B1(n_211),
.B2(n_209),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_224),
.C(n_216),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_231),
.B(n_199),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_227),
.C(n_250),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_199),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_225),
.A2(n_253),
.B1(n_241),
.B2(n_238),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_253),
.A2(n_217),
.B1(n_210),
.B2(n_198),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_229),
.B(n_242),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_234),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_295),
.A2(n_296),
.B1(n_310),
.B2(n_312),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_241),
.B1(n_227),
.B2(n_255),
.Y(n_296)
);

NOR3xp33_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_245),
.C(n_243),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_297),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

BUFx12f_ASAP7_75t_SL g299 ( 
.A(n_289),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_299),
.A2(n_288),
.B1(n_264),
.B2(n_278),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_300),
.A2(n_311),
.B1(n_313),
.B2(n_283),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_235),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_302),
.C(n_305),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_236),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_230),
.Y(n_304)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_259),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_307),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_198),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_287),
.B1(n_262),
.B2(n_276),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_188),
.B(n_256),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_188),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_316),
.A2(n_327),
.B1(n_329),
.B2(n_313),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_321),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_285),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_307),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_265),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_326),
.C(n_291),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_282),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_272),
.B1(n_273),
.B2(n_280),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_272),
.B1(n_267),
.B2(n_249),
.Y(n_329)
);

AOI211xp5_ASAP7_75t_L g334 ( 
.A1(n_299),
.A2(n_237),
.B(n_223),
.C(n_222),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_309),
.B(n_249),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_296),
.A2(n_203),
.A3(n_190),
.B1(n_222),
.B2(n_223),
.C1(n_213),
.C2(n_10),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_322),
.Y(n_342)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_328),
.Y(n_338)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_346),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_342),
.A2(n_320),
.B1(n_317),
.B2(n_319),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_343),
.A2(n_345),
.B1(n_351),
.B2(n_339),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_333),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_344),
.A2(n_312),
.B1(n_318),
.B2(n_190),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_323),
.A2(n_295),
.B1(n_300),
.B2(n_314),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_329),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_347),
.A2(n_348),
.B(n_353),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_330),
.A2(n_306),
.B(n_315),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_324),
.A2(n_301),
.B1(n_302),
.B2(n_308),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_349),
.A2(n_332),
.B1(n_350),
.B2(n_341),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_305),
.C(n_304),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_352),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_351),
.A2(n_352),
.B(n_353),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_292),
.B(n_294),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_327),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_357),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_356),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_346),
.B(n_321),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_347),
.A2(n_326),
.B1(n_317),
.B2(n_325),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_358),
.A2(n_343),
.B1(n_344),
.B2(n_338),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_362),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_351),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_348),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_339),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_367),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_360),
.A2(n_351),
.B(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_369),
.B(n_376),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_361),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_371),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_373),
.A2(n_340),
.B(n_364),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_373),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_377),
.B(n_378),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_375),
.A2(n_362),
.B1(n_366),
.B2(n_367),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_379),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_381),
.B(n_376),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_378),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_380),
.A2(n_368),
.B(n_374),
.Y(n_385)
);

AOI322xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_382),
.A3(n_340),
.B1(n_363),
.B2(n_337),
.C1(n_381),
.C2(n_365),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_388),
.C(n_372),
.Y(n_391)
);

AOI322xp5_ASAP7_75t_L g389 ( 
.A1(n_386),
.A2(n_342),
.A3(n_358),
.B1(n_354),
.B2(n_372),
.C1(n_357),
.C2(n_359),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_383),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_390),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_392),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_391),
.Y(n_394)
);


endmodule