module real_aes_7896_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_729;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_0), .A2(n_128), .B1(n_134), .B2(n_722), .C1(n_723), .C2(n_726), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_1), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g125 ( .A(n_1), .Y(n_125) );
INVx1_ASAP7_75t_L g463 ( .A(n_2), .Y(n_463) );
INVx1_ASAP7_75t_L g267 ( .A(n_3), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_4), .A2(n_37), .B1(n_217), .B2(n_502), .Y(n_538) );
AOI21xp33_ASAP7_75t_L g228 ( .A1(n_5), .A2(n_150), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_6), .B(n_172), .Y(n_488) );
AND2x6_ASAP7_75t_L g155 ( .A(n_7), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_8), .A2(n_149), .B(n_157), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_9), .B(n_38), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_10), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g234 ( .A(n_11), .Y(n_234) );
INVx1_ASAP7_75t_L g147 ( .A(n_12), .Y(n_147) );
INVx1_ASAP7_75t_L g457 ( .A(n_13), .Y(n_457) );
INVx1_ASAP7_75t_L g167 ( .A(n_14), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_15), .B(n_241), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_16), .B(n_173), .Y(n_490) );
AO32x2_ASAP7_75t_L g536 ( .A1(n_17), .A2(n_172), .A3(n_188), .B1(n_476), .B2(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_18), .B(n_217), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_19), .B(n_184), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_20), .B(n_173), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_21), .A2(n_49), .B1(n_217), .B2(n_502), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_22), .B(n_150), .Y(n_177) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_23), .A2(n_77), .B1(n_217), .B2(n_241), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_24), .B(n_217), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_25), .B(n_227), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_26), .A2(n_164), .B(n_166), .C(n_168), .Y(n_163) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_27), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_28), .B(n_143), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_29), .B(n_199), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_30), .A2(n_101), .B1(n_130), .B2(n_131), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_30), .Y(n_131) );
INVx1_ASAP7_75t_L g246 ( .A(n_31), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_32), .B(n_143), .Y(n_514) );
INVx2_ASAP7_75t_L g153 ( .A(n_33), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_34), .B(n_217), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_35), .B(n_143), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_36), .A2(n_155), .B(n_160), .C(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g244 ( .A(n_39), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_40), .B(n_199), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_41), .A2(n_104), .B1(n_115), .B2(n_742), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_42), .B(n_217), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_43), .A2(n_87), .B1(n_169), .B2(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_44), .B(n_217), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_45), .B(n_217), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_46), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_47), .B(n_462), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_48), .B(n_150), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_50), .A2(n_60), .B1(n_217), .B2(n_241), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_51), .A2(n_735), .B1(n_738), .B2(n_739), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_51), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_52), .A2(n_160), .B1(n_241), .B2(n_243), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_53), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_54), .B(n_217), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_55), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_56), .B(n_217), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_57), .A2(n_232), .B(n_233), .C(n_235), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_58), .Y(n_203) );
INVx1_ASAP7_75t_L g230 ( .A(n_59), .Y(n_230) );
INVx1_ASAP7_75t_L g156 ( .A(n_61), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_62), .A2(n_129), .B1(n_132), .B2(n_133), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_62), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_63), .B(n_217), .Y(n_464) );
INVx1_ASAP7_75t_L g146 ( .A(n_64), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_65), .A2(n_76), .B1(n_736), .B2(n_737), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_65), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
AO32x2_ASAP7_75t_L g499 ( .A1(n_67), .A2(n_172), .A3(n_209), .B1(n_476), .B2(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g474 ( .A(n_68), .Y(n_474) );
INVx1_ASAP7_75t_L g509 ( .A(n_69), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_SL g254 ( .A1(n_70), .A2(n_184), .B(n_235), .C(n_255), .Y(n_254) );
INVxp67_ASAP7_75t_L g256 ( .A(n_71), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_72), .B(n_241), .Y(n_510) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_74), .Y(n_249) );
INVx1_ASAP7_75t_L g194 ( .A(n_75), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_76), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_78), .A2(n_155), .B(n_160), .C(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_79), .B(n_502), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_80), .B(n_241), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_81), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_83), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_84), .B(n_241), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_85), .A2(n_155), .B(n_160), .C(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g109 ( .A(n_86), .Y(n_109) );
OR2x2_ASAP7_75t_L g122 ( .A(n_86), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g135 ( .A(n_86), .B(n_124), .Y(n_135) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_88), .A2(n_102), .B1(n_241), .B2(n_242), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_89), .B(n_143), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_90), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_91), .A2(n_155), .B(n_160), .C(n_212), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_92), .Y(n_220) );
INVx1_ASAP7_75t_L g253 ( .A(n_93), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g158 ( .A(n_94), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_95), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_96), .B(n_181), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_97), .B(n_241), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_98), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_100), .A2(n_150), .B(n_252), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_101), .Y(n_130) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g742 ( .A(n_106), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
OR2x2_ASAP7_75t_L g446 ( .A(n_109), .B(n_124), .Y(n_446) );
NOR2x2_ASAP7_75t_L g728 ( .A(n_109), .B(n_123), .Y(n_728) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g124 ( .A(n_114), .B(n_125), .Y(n_124) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_127), .B1(n_729), .B2(n_731), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g730 ( .A(n_119), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_120), .A2(n_732), .B(n_740), .Y(n_731) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_126), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g741 ( .A(n_122), .Y(n_741) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g722 ( .A(n_128), .Y(n_722) );
INVx1_ASAP7_75t_L g132 ( .A(n_129), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B1(n_444), .B2(n_447), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_135), .A2(n_446), .B1(n_724), .B2(n_725), .Y(n_723) );
INVx2_ASAP7_75t_SL g724 ( .A(n_136), .Y(n_724) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_136), .A2(n_724), .B1(n_733), .B2(n_734), .Y(n_732) );
OR4x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_340), .C(n_399), .D(n_426), .Y(n_136) );
NAND3xp33_ASAP7_75t_SL g137 ( .A(n_138), .B(n_282), .C(n_307), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_205), .B(n_225), .C(n_258), .Y(n_138) );
AOI211xp5_ASAP7_75t_SL g430 ( .A1(n_139), .A2(n_431), .B(n_433), .C(n_436), .Y(n_430) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_174), .Y(n_139) );
INVx1_ASAP7_75t_L g305 ( .A(n_140), .Y(n_305) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g280 ( .A(n_141), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g312 ( .A(n_141), .Y(n_312) );
AND2x2_ASAP7_75t_L g367 ( .A(n_141), .B(n_336), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_141), .B(n_223), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_141), .B(n_224), .Y(n_425) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g286 ( .A(n_142), .Y(n_286) );
AND2x2_ASAP7_75t_L g329 ( .A(n_142), .B(n_192), .Y(n_329) );
AND2x2_ASAP7_75t_L g347 ( .A(n_142), .B(n_224), .Y(n_347) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_148), .B(n_171), .Y(n_142) );
INVx1_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
INVx2_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_143), .A2(n_507), .B(n_514), .Y(n_506) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_143), .A2(n_516), .B(n_524), .Y(n_515) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_L g173 ( .A(n_144), .B(n_145), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_151), .B(n_155), .Y(n_195) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
INVx1_ASAP7_75t_L g462 ( .A(n_152), .Y(n_462) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
INVx1_ASAP7_75t_L g242 ( .A(n_153), .Y(n_242) );
INVx1_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
INVx3_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
INVx4_ASAP7_75t_SL g170 ( .A(n_155), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_155), .A2(n_456), .B(n_460), .Y(n_455) );
BUFx3_ASAP7_75t_L g476 ( .A(n_155), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_155), .A2(n_482), .B(n_485), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_155), .A2(n_508), .B(n_511), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_155), .A2(n_517), .B(n_521), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_163), .C(n_170), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_159), .A2(n_170), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_159), .A2(n_170), .B(n_253), .C(n_254), .Y(n_252) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
BUFx3_ASAP7_75t_L g169 ( .A(n_161), .Y(n_169) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
INVx1_ASAP7_75t_L g502 ( .A(n_161), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_164), .B(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g459 ( .A(n_164), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_164), .A2(n_512), .B(n_513), .Y(n_511) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g243 ( .A1(n_165), .A2(n_244), .B1(n_245), .B2(n_246), .Y(n_243) );
INVx2_ASAP7_75t_L g245 ( .A(n_165), .Y(n_245) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g186 ( .A(n_169), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g239 ( .A1(n_170), .A2(n_195), .B1(n_240), .B2(n_247), .Y(n_239) );
INVx4_ASAP7_75t_L g191 ( .A(n_172), .Y(n_191) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_172), .A2(n_251), .B(n_257), .Y(n_250) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_172), .A2(n_481), .B(n_488), .Y(n_480) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
INVx4_ASAP7_75t_L g279 ( .A(n_174), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_174), .A2(n_335), .B(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g415 ( .A(n_174), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_192), .Y(n_174) );
INVx1_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
AND2x2_ASAP7_75t_L g284 ( .A(n_175), .B(n_224), .Y(n_284) );
OR2x2_ASAP7_75t_L g313 ( .A(n_175), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g327 ( .A(n_175), .Y(n_327) );
INVx3_ASAP7_75t_L g336 ( .A(n_175), .Y(n_336) );
AND2x2_ASAP7_75t_L g346 ( .A(n_175), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g379 ( .A(n_175), .B(n_285), .Y(n_379) );
AND2x2_ASAP7_75t_L g403 ( .A(n_175), .B(n_359), .Y(n_403) );
OR2x6_ASAP7_75t_L g175 ( .A(n_176), .B(n_189), .Y(n_175) );
AOI21xp5_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_178), .B(n_187), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_183), .B(n_185), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_181), .A2(n_267), .B(n_268), .C(n_269), .Y(n_266) );
INVx2_ASAP7_75t_L g465 ( .A(n_181), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_181), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_181), .A2(n_483), .B(n_484), .Y(n_482) );
O2A1O1Ixp5_ASAP7_75t_SL g508 ( .A1(n_181), .A2(n_235), .B(n_509), .C(n_510), .Y(n_508) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_182), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_182), .B(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_SL g500 ( .A1(n_182), .A2(n_199), .B1(n_501), .B2(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g520 ( .A(n_184), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_185), .A2(n_198), .B(n_200), .Y(n_197) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g201 ( .A(n_187), .Y(n_201) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_187), .A2(n_455), .B(n_466), .Y(n_454) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_187), .A2(n_469), .B(n_477), .Y(n_468) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_188), .A2(n_239), .B(n_248), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_188), .B(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_188), .A2(n_263), .B(n_270), .Y(n_262) );
NOR2xp33_ASAP7_75t_SL g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx3_ASAP7_75t_L g227 ( .A(n_191), .Y(n_227) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_191), .B(n_476), .C(n_492), .Y(n_491) );
AO21x1_ASAP7_75t_L g570 ( .A1(n_191), .A2(n_492), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g224 ( .A(n_192), .Y(n_224) );
AND2x2_ASAP7_75t_L g439 ( .A(n_192), .B(n_281), .Y(n_439) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_201), .B(n_202), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_195), .A2(n_264), .B(n_265), .Y(n_263) );
INVx4_ASAP7_75t_L g215 ( .A(n_199), .Y(n_215) );
INVx2_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_199), .A2(n_465), .B1(n_493), .B2(n_494), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_199), .A2(n_465), .B1(n_538), .B2(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_204), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_204), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_221), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_207), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g359 ( .A(n_207), .B(n_347), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_207), .B(n_336), .Y(n_421) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g281 ( .A(n_208), .Y(n_281) );
AND2x2_ASAP7_75t_L g285 ( .A(n_208), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g326 ( .A(n_208), .B(n_327), .Y(n_326) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_219), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_218), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_216), .Y(n_212) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_221), .B(n_322), .Y(n_344) );
INVx1_ASAP7_75t_L g383 ( .A(n_221), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_221), .B(n_310), .Y(n_427) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
AND2x2_ASAP7_75t_L g290 ( .A(n_222), .B(n_285), .Y(n_290) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_224), .B(n_281), .Y(n_314) );
INVx1_ASAP7_75t_L g393 ( .A(n_224), .Y(n_393) );
AOI322xp5_ASAP7_75t_L g417 ( .A1(n_225), .A2(n_332), .A3(n_392), .B1(n_418), .B2(n_420), .C1(n_422), .C2(n_424), .Y(n_417) );
AND2x2_ASAP7_75t_SL g225 ( .A(n_226), .B(n_237), .Y(n_225) );
AND2x2_ASAP7_75t_L g272 ( .A(n_226), .B(n_250), .Y(n_272) );
INVx1_ASAP7_75t_SL g275 ( .A(n_226), .Y(n_275) );
AND2x2_ASAP7_75t_L g277 ( .A(n_226), .B(n_238), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_226), .B(n_294), .Y(n_300) );
INVx2_ASAP7_75t_L g319 ( .A(n_226), .Y(n_319) );
AND2x2_ASAP7_75t_L g332 ( .A(n_226), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g370 ( .A(n_226), .B(n_294), .Y(n_370) );
BUFx2_ASAP7_75t_L g387 ( .A(n_226), .Y(n_387) );
AND2x2_ASAP7_75t_L g401 ( .A(n_226), .B(n_261), .Y(n_401) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_236), .Y(n_226) );
O2A1O1Ixp5_ASAP7_75t_L g473 ( .A1(n_232), .A2(n_461), .B(n_474), .C(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_232), .A2(n_522), .B(n_523), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_237), .B(n_289), .Y(n_316) );
AND2x2_ASAP7_75t_L g443 ( .A(n_237), .B(n_319), .Y(n_443) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_250), .Y(n_237) );
OR2x2_ASAP7_75t_L g288 ( .A(n_238), .B(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g294 ( .A(n_238), .Y(n_294) );
AND2x2_ASAP7_75t_L g339 ( .A(n_238), .B(n_262), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_238), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_238), .Y(n_423) );
INVx2_ASAP7_75t_L g269 ( .A(n_241), .Y(n_269) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g274 ( .A(n_250), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g296 ( .A(n_250), .Y(n_296) );
BUFx2_ASAP7_75t_L g302 ( .A(n_250), .Y(n_302) );
AND2x2_ASAP7_75t_L g321 ( .A(n_250), .B(n_294), .Y(n_321) );
INVx3_ASAP7_75t_L g333 ( .A(n_250), .Y(n_333) );
OR2x2_ASAP7_75t_L g343 ( .A(n_250), .B(n_294), .Y(n_343) );
AOI31xp33_ASAP7_75t_SL g258 ( .A1(n_259), .A2(n_273), .A3(n_276), .B(n_278), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_272), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_260), .B(n_295), .Y(n_306) );
OR2x2_ASAP7_75t_L g330 ( .A(n_260), .B(n_300), .Y(n_330) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_261), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g351 ( .A(n_261), .B(n_343), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_261), .B(n_333), .Y(n_361) );
AND2x2_ASAP7_75t_L g368 ( .A(n_261), .B(n_369), .Y(n_368) );
NAND2x1_ASAP7_75t_L g396 ( .A(n_261), .B(n_332), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_261), .B(n_387), .Y(n_397) );
AND2x2_ASAP7_75t_L g409 ( .A(n_261), .B(n_294), .Y(n_409) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g289 ( .A(n_262), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_269), .A2(n_457), .B(n_458), .C(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g355 ( .A(n_272), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_272), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_274), .B(n_350), .Y(n_384) );
AND2x4_ASAP7_75t_L g295 ( .A(n_275), .B(n_296), .Y(n_295) );
CKINVDCx16_ASAP7_75t_R g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g374 ( .A(n_280), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_280), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g322 ( .A(n_281), .B(n_312), .Y(n_322) );
AND2x2_ASAP7_75t_L g416 ( .A(n_281), .B(n_286), .Y(n_416) );
INVx1_ASAP7_75t_L g441 ( .A(n_281), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B1(n_290), .B2(n_291), .C(n_297), .Y(n_282) );
CKINVDCx14_ASAP7_75t_R g303 ( .A(n_283), .Y(n_303) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_284), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_287), .B(n_338), .Y(n_357) );
INVx3_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g406 ( .A(n_288), .B(n_302), .Y(n_406) );
AND2x2_ASAP7_75t_L g320 ( .A(n_289), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g350 ( .A(n_289), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_289), .B(n_333), .Y(n_378) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_289), .B(n_390), .C(n_421), .Y(n_420) );
AOI211xp5_ASAP7_75t_SL g353 ( .A1(n_290), .A2(n_354), .B(n_356), .C(n_364), .Y(n_353) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_292), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_293), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_293), .B(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g435 ( .A(n_295), .B(n_409), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_303), .B1(n_304), .B2(n_306), .Y(n_297) );
NOR2xp33_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_301), .B(n_350), .Y(n_381) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_304), .A2(n_396), .B1(n_427), .B2(n_434), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_315), .B1(n_317), .B2(n_322), .C(n_323), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_313), .A2(n_324), .B1(n_330), .B2(n_331), .C(n_334), .Y(n_323) );
INVx1_ASAP7_75t_L g366 ( .A(n_314), .Y(n_366) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_SL g338 ( .A(n_319), .Y(n_338) );
OR2x2_ASAP7_75t_L g411 ( .A(n_319), .B(n_343), .Y(n_411) );
AND2x2_ASAP7_75t_L g413 ( .A(n_319), .B(n_321), .Y(n_413) );
INVx1_ASAP7_75t_L g352 ( .A(n_322), .Y(n_352) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
AOI21xp33_ASAP7_75t_SL g382 ( .A1(n_325), .A2(n_383), .B(n_384), .Y(n_382) );
OR2x2_ASAP7_75t_L g389 ( .A(n_325), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g363 ( .A(n_326), .B(n_347), .Y(n_363) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_331), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_332), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_333), .B(n_369), .Y(n_432) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_336), .A2(n_349), .B(n_351), .C(n_352), .Y(n_348) );
NAND2x1_ASAP7_75t_SL g373 ( .A(n_336), .B(n_374), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_337), .A2(n_386), .B1(n_388), .B2(n_391), .Y(n_385) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_339), .B(n_429), .Y(n_428) );
NAND5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_353), .C(n_371), .D(n_385), .E(n_394), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_348), .Y(n_341) );
INVx1_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_346), .A2(n_365), .B1(n_405), .B2(n_407), .C(n_410), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_347), .B(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_350), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_350), .B(n_416), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_360), .B2(n_362), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_368), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g438 ( .A(n_367), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B1(n_379), .B2(n_380), .C(n_382), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g422 ( .A(n_377), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g429 ( .A(n_387), .Y(n_429) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_397), .B(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_402), .B(n_404), .C(n_417), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_402), .A2(n_427), .B(n_428), .C(n_430), .Y(n_426) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_406), .B(n_408), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_440), .B(n_442), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g725 ( .A(n_447), .Y(n_725) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR5x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_613), .C(n_671), .D(n_707), .E(n_714), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_559), .C(n_583), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_495), .B1(n_525), .B2(n_530), .C(n_540), .Y(n_451) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_452), .A2(n_694), .B(n_696), .Y(n_693) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_478), .Y(n_452) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_453), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_467), .Y(n_453) );
INVx2_ASAP7_75t_L g529 ( .A(n_454), .Y(n_529) );
AND2x2_ASAP7_75t_L g542 ( .A(n_454), .B(n_480), .Y(n_542) );
AND2x2_ASAP7_75t_L g596 ( .A(n_454), .B(n_479), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_454), .B(n_468), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B(n_464), .C(n_465), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_465), .A2(n_486), .B(n_487), .Y(n_485) );
AND2x2_ASAP7_75t_L g629 ( .A(n_467), .B(n_570), .Y(n_629) );
AND2x2_ASAP7_75t_L g662 ( .A(n_467), .B(n_480), .Y(n_662) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g569 ( .A(n_468), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g582 ( .A(n_468), .B(n_480), .Y(n_582) );
AND2x2_ASAP7_75t_L g589 ( .A(n_468), .B(n_570), .Y(n_589) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_468), .Y(n_598) );
AND2x2_ASAP7_75t_L g605 ( .A(n_468), .B(n_479), .Y(n_605) );
INVx1_ASAP7_75t_L g636 ( .A(n_468), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_473), .B(n_476), .Y(n_469) );
INVx1_ASAP7_75t_L g612 ( .A(n_478), .Y(n_612) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
INVx2_ASAP7_75t_L g568 ( .A(n_479), .Y(n_568) );
AND2x2_ASAP7_75t_L g590 ( .A(n_479), .B(n_529), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_479), .B(n_636), .Y(n_641) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_480), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g713 ( .A(n_480), .B(n_677), .Y(n_713) );
INVx2_ASAP7_75t_L g527 ( .A(n_489), .Y(n_527) );
INVx3_ASAP7_75t_L g628 ( .A(n_489), .Y(n_628) );
OR2x2_ASAP7_75t_L g658 ( .A(n_489), .B(n_659), .Y(n_658) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_489), .B(n_568), .Y(n_684) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g571 ( .A(n_490), .Y(n_571) );
AOI33xp33_ASAP7_75t_L g704 ( .A1(n_495), .A2(n_542), .A3(n_556), .B1(n_628), .B2(n_705), .B3(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_504), .Y(n_496) );
OR2x2_ASAP7_75t_L g557 ( .A(n_497), .B(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_497), .B(n_554), .Y(n_616) );
OR2x2_ASAP7_75t_L g669 ( .A(n_497), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g595 ( .A(n_498), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g620 ( .A(n_498), .B(n_504), .Y(n_620) );
AND2x2_ASAP7_75t_L g687 ( .A(n_498), .B(n_532), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_498), .A2(n_587), .B(n_713), .Y(n_712) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g534 ( .A(n_499), .Y(n_534) );
INVx1_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
AND2x2_ASAP7_75t_L g566 ( .A(n_499), .B(n_536), .Y(n_566) );
AND2x2_ASAP7_75t_L g615 ( .A(n_499), .B(n_535), .Y(n_615) );
INVx2_ASAP7_75t_SL g657 ( .A(n_504), .Y(n_657) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_515), .Y(n_504) );
INVx2_ASAP7_75t_L g577 ( .A(n_505), .Y(n_577) );
INVx1_ASAP7_75t_L g708 ( .A(n_505), .Y(n_708) );
AND2x2_ASAP7_75t_L g721 ( .A(n_505), .B(n_602), .Y(n_721) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g548 ( .A(n_506), .Y(n_548) );
OR2x2_ASAP7_75t_L g554 ( .A(n_506), .B(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_506), .Y(n_565) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_515), .Y(n_532) );
AND2x2_ASAP7_75t_L g549 ( .A(n_515), .B(n_535), .Y(n_549) );
INVx1_ASAP7_75t_L g555 ( .A(n_515), .Y(n_555) );
INVx1_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
AND2x2_ASAP7_75t_L g587 ( .A(n_515), .B(n_536), .Y(n_587) );
INVx2_ASAP7_75t_L g603 ( .A(n_515), .Y(n_603) );
AND2x2_ASAP7_75t_L g696 ( .A(n_515), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_515), .B(n_577), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
INVx1_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g551 ( .A(n_527), .Y(n_551) );
INVx1_ASAP7_75t_L g580 ( .A(n_527), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_527), .B(n_611), .Y(n_677) );
INVx1_ASAP7_75t_SL g637 ( .A(n_528), .Y(n_637) );
INVx2_ASAP7_75t_L g558 ( .A(n_529), .Y(n_558) );
AND2x2_ASAP7_75t_L g627 ( .A(n_529), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g643 ( .A(n_529), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_L g705 ( .A(n_531), .Y(n_705) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g560 ( .A(n_533), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g663 ( .A(n_533), .B(n_653), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_533), .A2(n_674), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g576 ( .A(n_534), .B(n_577), .Y(n_576) );
BUFx2_ASAP7_75t_L g601 ( .A(n_534), .Y(n_601) );
INVx1_ASAP7_75t_L g625 ( .A(n_534), .Y(n_625) );
OR2x2_ASAP7_75t_L g689 ( .A(n_535), .B(n_548), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g697 ( .A(n_535), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g602 ( .A(n_536), .B(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_L g609 ( .A(n_536), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_543), .B1(n_550), .B2(n_552), .Y(n_540) );
OR2x2_ASAP7_75t_L g619 ( .A(n_541), .B(n_569), .Y(n_619) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g660 ( .A1(n_542), .A2(n_661), .B1(n_663), .B2(n_664), .C1(n_665), .C2(n_668), .Y(n_660) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g607 ( .A(n_546), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_548), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_548), .Y(n_632) );
AND2x2_ASAP7_75t_L g680 ( .A(n_548), .B(n_549), .Y(n_680) );
INVx1_ASAP7_75t_L g698 ( .A(n_548), .Y(n_698) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g664 ( .A(n_551), .B(n_590), .Y(n_664) );
AND2x2_ASAP7_75t_L g706 ( .A(n_551), .B(n_582), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_553), .B(n_601), .Y(n_688) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_554), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g581 ( .A(n_558), .B(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g649 ( .A(n_558), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B(n_567), .C(n_572), .Y(n_559) );
INVxp67_ASAP7_75t_L g573 ( .A(n_560), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_561), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_561), .B(n_608), .Y(n_703) );
BUFx3_ASAP7_75t_L g667 ( .A(n_562), .Y(n_667) );
INVx1_ASAP7_75t_L g574 ( .A(n_563), .Y(n_574) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g593 ( .A(n_565), .B(n_587), .Y(n_593) );
INVx1_ASAP7_75t_SL g633 ( .A(n_566), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g623 ( .A(n_568), .Y(n_623) );
AND2x2_ASAP7_75t_L g646 ( .A(n_568), .B(n_629), .Y(n_646) );
INVx1_ASAP7_75t_SL g617 ( .A(n_569), .Y(n_617) );
INVx1_ASAP7_75t_L g644 ( .A(n_570), .Y(n_644) );
AOI31xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .A3(n_575), .B(n_578), .Y(n_572) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g665 ( .A(n_576), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g639 ( .A(n_577), .Y(n_639) );
BUFx2_ASAP7_75t_L g653 ( .A(n_577), .Y(n_653) );
AND2x2_ASAP7_75t_L g681 ( .A(n_577), .B(n_602), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g654 ( .A(n_581), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_582), .B(n_649), .Y(n_695) );
AND2x2_ASAP7_75t_L g702 ( .A(n_582), .B(n_628), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_588), .B(n_591), .C(n_606), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_588), .A2(n_615), .B1(n_616), .B2(n_617), .C(n_618), .Y(n_614) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g622 ( .A(n_589), .B(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g659 ( .A(n_590), .Y(n_659) );
OAI32xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .A3(n_597), .B1(n_599), .B2(n_604), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_593), .A2(n_646), .B(n_647), .C(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_601), .A2(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g670 ( .A(n_602), .Y(n_670) );
INVxp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_608), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g656 ( .A(n_608), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g673 ( .A(n_610), .Y(n_673) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND4xp25_ASAP7_75t_SL g613 ( .A(n_614), .B(n_626), .C(n_645), .D(n_660), .Y(n_613) );
AND2x2_ASAP7_75t_L g652 ( .A(n_615), .B(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g674 ( .A(n_615), .B(n_667), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_617), .B(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B1(n_621), .B2(n_624), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_619), .A2(n_670), .B1(n_701), .B2(n_703), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_619), .A2(n_708), .B(n_709), .C(n_712), .Y(n_707) );
INVx2_ASAP7_75t_L g678 ( .A(n_620), .Y(n_678) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_622), .A2(n_656), .B1(n_673), .B2(n_674), .C1(n_675), .C2(n_678), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_630), .C(n_634), .Y(n_626) );
INVx1_ASAP7_75t_L g692 ( .A(n_627), .Y(n_692) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_631), .A2(n_635), .B1(n_638), .B2(n_640), .Y(n_634) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g661 ( .A(n_643), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g719 ( .A(n_646), .Y(n_719) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_655), .B2(n_658), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_653), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g710 ( .A(n_658), .Y(n_710) );
INVx1_ASAP7_75t_L g691 ( .A(n_662), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g718 ( .A(n_664), .Y(n_718) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND5xp2_ASAP7_75t_L g671 ( .A(n_672), .B(n_679), .C(n_693), .D(n_699), .E(n_704), .Y(n_671) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B(n_682), .C(n_685), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI31xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .A3(n_689), .B(n_690), .Y(n_685) );
INVx1_ASAP7_75t_L g711 ( .A(n_687), .Y(n_711) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI222xp33_ASAP7_75t_L g714 ( .A1(n_701), .A2(n_703), .B1(n_715), .B2(n_718), .C1(n_719), .C2(n_720), .Y(n_714) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
CKINVDCx14_ASAP7_75t_R g739 ( .A(n_735), .Y(n_739) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
endmodule