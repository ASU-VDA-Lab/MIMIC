module fake_aes_1818_n_1118 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1118);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1118;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_345;
wire n_360;
wire n_1090;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1078;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1024;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_1046;
wire n_460;
wire n_910;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_192), .Y(n_254) );
INVxp67_ASAP7_75t_L g255 ( .A(n_11), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_247), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_81), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_207), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_190), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_242), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_91), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_181), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_52), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_66), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_132), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_128), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_29), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_1), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_143), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_161), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_9), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_184), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_123), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_243), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_11), .Y(n_279) );
CKINVDCx16_ASAP7_75t_R g280 ( .A(n_135), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_82), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_116), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_234), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_164), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_33), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_75), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_178), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_140), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_92), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_15), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_4), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_213), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_89), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_125), .Y(n_294) );
INVxp33_ASAP7_75t_L g295 ( .A(n_93), .Y(n_295) );
BUFx2_ASAP7_75t_SL g296 ( .A(n_146), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_71), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_94), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_26), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_48), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_230), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_97), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_245), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_105), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_6), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_107), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_211), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_170), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_17), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_10), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_197), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_159), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_47), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_100), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_62), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_122), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_57), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_232), .Y(n_318) );
BUFx10_ASAP7_75t_L g319 ( .A(n_163), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_195), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_10), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_141), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_0), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_57), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_60), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_114), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_217), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_171), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_238), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_35), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_19), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_244), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_228), .Y(n_333) );
CKINVDCx14_ASAP7_75t_R g334 ( .A(n_223), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_19), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_108), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_45), .Y(n_337) );
CKINVDCx14_ASAP7_75t_R g338 ( .A(n_172), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_151), .Y(n_339) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_41), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_64), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_224), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_4), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_183), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_204), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_69), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_39), .Y(n_347) );
INVxp33_ASAP7_75t_SL g348 ( .A(n_60), .Y(n_348) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_56), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_30), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_33), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_150), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_67), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_226), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_121), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_136), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_252), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_38), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_168), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_90), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_246), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_144), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_64), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_20), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_119), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_53), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_165), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_86), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_225), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_50), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_53), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_120), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_194), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_79), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_22), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_157), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_42), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_32), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_118), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_130), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_221), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_26), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_49), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_99), .B(n_149), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_137), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_250), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_31), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_203), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_175), .Y(n_389) );
CKINVDCx16_ASAP7_75t_R g390 ( .A(n_29), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_311), .B(n_305), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_311), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_288), .Y(n_393) );
INVx5_ASAP7_75t_L g394 ( .A(n_311), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_288), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_305), .B(n_0), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_348), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_261), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
OAI22x1_ASAP7_75t_L g400 ( .A1(n_358), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_382), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_319), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_261), .Y(n_403) );
OAI22xp5_ASAP7_75t_SL g404 ( .A1(n_343), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_261), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_261), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_289), .Y(n_407) );
CKINVDCx6p67_ASAP7_75t_R g408 ( .A(n_280), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_261), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_382), .B(n_7), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_323), .B(n_8), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_289), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_265), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_268), .B(n_8), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_265), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_323), .B(n_9), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_271), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_333), .Y(n_418) );
OAI22xp5_ASAP7_75t_SL g419 ( .A1(n_343), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_333), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_271), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_324), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_324), .Y(n_423) );
INVx4_ASAP7_75t_L g424 ( .A(n_319), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_391), .B(n_302), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_391), .B(n_320), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_393), .B(n_256), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_392), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_403), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_392), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_391), .B(n_385), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_393), .A2(n_279), .B1(n_285), .B2(n_274), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_399), .B(n_319), .Y(n_434) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_396), .B(n_384), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_399), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_395), .B(n_256), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_424), .B(n_301), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_395), .A2(n_297), .B1(n_299), .B2(n_291), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_424), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_391), .B(n_282), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_407), .B(n_282), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_403), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
OR2x6_ASAP7_75t_L g446 ( .A(n_400), .B(n_296), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_407), .B(n_257), .C(n_253), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_394), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_424), .B(n_352), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_412), .A2(n_300), .B1(n_321), .B2(n_309), .Y(n_450) );
BUFx10_ASAP7_75t_L g451 ( .A(n_396), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_412), .B(n_292), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_394), .B(n_292), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_396), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_396), .A2(n_325), .B1(n_335), .B2(n_331), .Y(n_455) );
NAND2xp33_ASAP7_75t_L g456 ( .A(n_402), .B(n_262), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_401), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_394), .B(n_304), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_394), .B(n_304), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_404), .B(n_419), .C(n_390), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_424), .B(n_334), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_403), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_411), .B(n_312), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_402), .B(n_338), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_403), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_402), .B(n_312), .Y(n_470) );
INVx2_ASAP7_75t_SL g471 ( .A(n_439), .Y(n_471) );
INVxp33_ASAP7_75t_L g472 ( .A(n_434), .Y(n_472) );
NAND3xp33_ASAP7_75t_SL g473 ( .A(n_455), .B(n_397), .C(n_290), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_441), .B(n_410), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_425), .B(n_414), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_441), .B(n_262), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_425), .B(n_408), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_436), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_426), .B(n_432), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_461), .B(n_263), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_435), .A2(n_408), .B1(n_348), .B2(n_342), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_454), .A2(n_416), .B(n_415), .C(n_413), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_436), .B(n_340), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_428), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_461), .B(n_263), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_461), .B(n_273), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_455), .B(n_397), .C(n_290), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_457), .B(n_270), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_426), .B(n_273), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_463), .A2(n_415), .B(n_417), .C(n_413), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_439), .B(n_416), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_432), .B(n_295), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_468), .B(n_277), .Y(n_494) );
OR2x6_ASAP7_75t_L g495 ( .A(n_439), .B(n_404), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_468), .B(n_277), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_467), .A2(n_355), .B(n_314), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_449), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_449), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_435), .A2(n_342), .B1(n_345), .B2(n_260), .Y(n_501) );
INVx8_ASAP7_75t_L g502 ( .A(n_449), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_463), .B(n_417), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_434), .B(n_283), .Y(n_504) );
AND2x6_ASAP7_75t_SL g505 ( .A(n_446), .B(n_419), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_430), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_434), .B(n_287), .Y(n_507) );
INVx5_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_430), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_457), .A2(n_345), .B1(n_373), .B2(n_260), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_442), .B(n_464), .Y(n_511) );
BUFx3_ASAP7_75t_L g512 ( .A(n_431), .Y(n_512) );
BUFx8_ASAP7_75t_L g513 ( .A(n_460), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_431), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_465), .B(n_287), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_465), .A2(n_400), .B1(n_422), .B2(n_421), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_465), .B(n_294), .Y(n_517) );
NOR2xp33_ASAP7_75t_R g518 ( .A(n_451), .B(n_373), .Y(n_518) );
AND2x2_ASAP7_75t_SL g519 ( .A(n_460), .B(n_384), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_456), .B(n_421), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_454), .A2(n_423), .B(n_422), .C(n_366), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_445), .Y(n_522) );
BUFx8_ASAP7_75t_L g523 ( .A(n_446), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_454), .B(n_307), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_445), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_466), .B(n_307), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_466), .B(n_329), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_466), .B(n_329), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_433), .B(n_270), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_467), .B(n_423), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_466), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_443), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_443), .Y(n_533) );
BUFx2_ASAP7_75t_L g534 ( .A(n_446), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_470), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_437), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_452), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_470), .B(n_275), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_446), .A2(n_337), .B1(n_346), .B2(n_341), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_433), .B(n_360), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_427), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_440), .B(n_360), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_427), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_440), .A2(n_315), .B1(n_317), .B2(n_313), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_450), .B(n_372), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_472), .B(n_477), .Y(n_546) );
AOI21xp5_ASAP7_75t_SL g547 ( .A1(n_532), .A2(n_459), .B(n_458), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_478), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_533), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_475), .B(n_450), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_537), .Y(n_551) );
NOR3xp33_ASAP7_75t_SL g552 ( .A(n_473), .B(n_315), .C(n_313), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_475), .B(n_438), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_479), .A2(n_446), .B1(n_447), .B2(n_363), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_512), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_471), .A2(n_498), .B1(n_499), .B2(n_473), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_502), .B(n_492), .Y(n_557) );
BUFx12f_ASAP7_75t_L g558 ( .A(n_505), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_493), .B(n_438), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_493), .B(n_446), .Y(n_560) );
NOR2xp33_ASAP7_75t_SL g561 ( .A(n_508), .B(n_446), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_508), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_511), .A2(n_453), .B(n_458), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_474), .B(n_317), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_483), .A2(n_459), .B(n_453), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_502), .B(n_330), .Y(n_566) );
NOR2xp33_ASAP7_75t_R g567 ( .A(n_523), .B(n_502), .Y(n_567) );
OAI22xp5_ASAP7_75t_SL g568 ( .A1(n_495), .A2(n_363), .B1(n_387), .B2(n_330), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_531), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_492), .B(n_387), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_490), .B(n_255), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_508), .B(n_376), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_484), .B(n_266), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_508), .B(n_349), .Y(n_574) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_497), .A2(n_448), .B(n_444), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_480), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_500), .B(n_376), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_489), .B(n_371), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_526), .A2(n_445), .B(n_365), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_528), .A2(n_445), .B(n_386), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_518), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_485), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_504), .B(n_310), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_507), .B(n_388), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_523), .Y(n_585) );
BUFx4f_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_491), .A2(n_366), .B(n_370), .C(n_351), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_534), .B(n_375), .Y(n_588) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_491), .A2(n_364), .B(n_378), .C(n_377), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_510), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_506), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_482), .B(n_383), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_503), .B(n_364), .Y(n_593) );
NAND3xp33_ASAP7_75t_SL g594 ( .A(n_516), .B(n_259), .C(n_258), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_494), .B(n_264), .Y(n_595) );
BUFx4f_ASAP7_75t_L g596 ( .A(n_495), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_503), .B(n_347), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_544), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_496), .B(n_267), .Y(n_599) );
AO32x2_ASAP7_75t_L g600 ( .A1(n_535), .A2(n_296), .A3(n_403), .B1(n_405), .B2(n_333), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_522), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_521), .A2(n_353), .B(n_347), .C(n_269), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_529), .B(n_353), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_540), .A2(n_272), .B(n_278), .C(n_276), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_515), .B(n_281), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_542), .B(n_350), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_501), .A2(n_350), .B1(n_284), .B2(n_293), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
NAND3xp33_ASAP7_75t_SL g610 ( .A(n_516), .B(n_298), .C(n_286), .Y(n_610) );
BUFx8_ASAP7_75t_L g611 ( .A(n_541), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_539), .B(n_303), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_509), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_522), .Y(n_614) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_514), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_522), .Y(n_616) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_525), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_543), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_530), .A2(n_306), .B(n_316), .C(n_308), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_530), .A2(n_322), .B(n_326), .C(n_318), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_481), .A2(n_444), .B(n_429), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_525), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_525), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_488), .B(n_254), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_539), .A2(n_328), .B(n_327), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_545), .B(n_350), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_486), .A2(n_462), .B(n_336), .Y(n_627) );
AOI33xp33_ASAP7_75t_L g628 ( .A1(n_519), .A2(n_367), .A3(n_332), .B1(n_339), .B2(n_344), .B3(n_389), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_520), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_487), .A2(n_356), .B(n_357), .C(n_354), .Y(n_630) );
AO21x1_ASAP7_75t_L g631 ( .A1(n_497), .A2(n_361), .B(n_359), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_525), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_520), .A2(n_368), .B(n_369), .C(n_362), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_524), .A2(n_462), .B(n_379), .Y(n_634) );
INVx4_ASAP7_75t_L g635 ( .A(n_536), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_476), .B(n_350), .Y(n_636) );
INVx5_ASAP7_75t_L g637 ( .A(n_519), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_527), .B(n_374), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_538), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_513), .B(n_380), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_478), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_475), .B(n_254), .Y(n_642) );
INVx4_ASAP7_75t_L g643 ( .A(n_508), .Y(n_643) );
NOR2xp33_ASAP7_75t_R g644 ( .A(n_478), .B(n_12), .Y(n_644) );
OAI22x1_ASAP7_75t_L g645 ( .A1(n_510), .A2(n_314), .B1(n_355), .B2(n_15), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_491), .A2(n_381), .B(n_398), .C(n_406), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_491), .A2(n_398), .B(n_406), .C(n_409), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_478), .B(n_13), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_532), .A2(n_398), .B1(n_409), .B2(n_418), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_478), .B(n_14), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_478), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_532), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_478), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_532), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_511), .A2(n_418), .B(n_409), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_511), .A2(n_420), .B(n_469), .Y(n_656) );
BUFx4f_ASAP7_75t_L g657 ( .A(n_502), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_475), .B(n_16), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_549), .B(n_16), .Y(n_659) );
AO31x2_ASAP7_75t_L g660 ( .A1(n_631), .A2(n_420), .A3(n_403), .B(n_405), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_590), .B(n_17), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_554), .A2(n_333), .B1(n_405), .B2(n_21), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_551), .B(n_18), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_651), .B(n_18), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_563), .A2(n_405), .B(n_72), .Y(n_665) );
OAI21x1_ASAP7_75t_SL g666 ( .A1(n_643), .A2(n_20), .B(n_21), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_651), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_667) );
BUFx12f_ASAP7_75t_L g668 ( .A(n_641), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_592), .A2(n_405), .B1(n_24), .B2(n_25), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_629), .A2(n_405), .B(n_469), .C(n_27), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_652), .B(n_23), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_557), .B(n_25), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_553), .A2(n_469), .B(n_74), .Y(n_673) );
OAI21x1_ASAP7_75t_L g674 ( .A1(n_575), .A2(n_469), .B(n_76), .Y(n_674) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_552), .A2(n_27), .B(n_28), .C(n_30), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_550), .A2(n_469), .B(n_77), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_568), .A2(n_469), .B1(n_31), .B2(n_32), .Y(n_677) );
BUFx2_ASAP7_75t_L g678 ( .A(n_548), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_559), .A2(n_469), .B(n_78), .Y(n_679) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_643), .Y(n_680) );
O2A1O1Ixp33_ASAP7_75t_L g681 ( .A1(n_589), .A2(n_28), .B(n_34), .C(n_35), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_654), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_547), .A2(n_80), .B(n_73), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_576), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_582), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_546), .B(n_34), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_639), .B(n_36), .Y(n_687) );
INVx1_ASAP7_75t_SL g688 ( .A(n_653), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_568), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_591), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_617), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_586), .A2(n_37), .B1(n_39), .B2(n_40), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g693 ( .A(n_567), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_565), .A2(n_84), .B(n_83), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_628), .B(n_40), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_556), .B(n_41), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_560), .A2(n_87), .B(n_85), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_573), .A2(n_42), .B1(n_43), .B2(n_44), .C(n_45), .Y(n_698) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_656), .A2(n_155), .B(n_249), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_613), .Y(n_700) );
AOI221xp5_ASAP7_75t_SL g701 ( .A1(n_587), .A2(n_43), .B1(n_44), .B2(n_46), .C(n_47), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_618), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_566), .B(n_46), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_658), .Y(n_704) );
INVxp67_ASAP7_75t_L g705 ( .A(n_648), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_615), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_637), .B(n_48), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_603), .B(n_49), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_606), .A2(n_158), .B(n_248), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_617), .Y(n_710) );
NOR2xp33_ASAP7_75t_SL g711 ( .A(n_657), .B(n_88), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_586), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_712) );
AOI221x1_ASAP7_75t_L g713 ( .A1(n_645), .A2(n_51), .B1(n_54), .B2(n_55), .C(n_56), .Y(n_713) );
INVx1_ASAP7_75t_SL g714 ( .A(n_574), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_657), .Y(n_715) );
AOI221xp5_ASAP7_75t_SL g716 ( .A1(n_646), .A2(n_54), .B1(n_55), .B2(n_58), .C(n_59), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_602), .A2(n_58), .B(n_59), .C(n_61), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_578), .B(n_61), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_579), .A2(n_166), .B(n_241), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_598), .A2(n_62), .B1(n_63), .B2(n_65), .Y(n_720) );
OAI21x1_ASAP7_75t_L g721 ( .A1(n_621), .A2(n_162), .B(n_240), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_561), .B(n_63), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_596), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_723) );
OAI21x1_ASAP7_75t_L g724 ( .A1(n_655), .A2(n_169), .B(n_239), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_609), .B(n_564), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_580), .A2(n_167), .B(n_237), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_585), .B(n_68), .Y(n_727) );
OAI21x1_ASAP7_75t_SL g728 ( .A1(n_635), .A2(n_68), .B(n_69), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_604), .A2(n_70), .B(n_71), .C(n_95), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_642), .A2(n_174), .B(n_96), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_637), .B(n_70), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_637), .B(n_98), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_583), .B(n_101), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_570), .B(n_102), .Y(n_734) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_601), .A2(n_103), .B(n_104), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_650), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_647), .A2(n_106), .B(n_109), .C(n_110), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g738 ( .A(n_644), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_574), .Y(n_739) );
AO31x2_ASAP7_75t_L g740 ( .A1(n_619), .A2(n_111), .A3(n_112), .B(n_113), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_596), .B(n_115), .Y(n_741) );
AOI222xp33_ASAP7_75t_SL g742 ( .A1(n_608), .A2(n_117), .B1(n_124), .B2(n_126), .C1(n_127), .C2(n_129), .Y(n_742) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_617), .Y(n_743) );
INVx6_ASAP7_75t_L g744 ( .A(n_611), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_L g745 ( .A1(n_633), .A2(n_131), .B(n_133), .C(n_134), .Y(n_745) );
AO32x2_ASAP7_75t_L g746 ( .A1(n_649), .A2(n_138), .A3(n_139), .B1(n_142), .B2(n_145), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_588), .A2(n_147), .B1(n_148), .B2(n_152), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_624), .B(n_153), .C(n_154), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_625), .A2(n_156), .B(n_160), .C(n_173), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_588), .B(n_176), .Y(n_750) );
BUFx4f_ASAP7_75t_L g751 ( .A(n_558), .Y(n_751) );
AO31x2_ASAP7_75t_L g752 ( .A1(n_620), .A2(n_177), .A3(n_180), .B(n_182), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_562), .B(n_251), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_593), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_595), .A2(n_185), .B(n_186), .C(n_187), .Y(n_755) );
BUFx2_ASAP7_75t_R g756 ( .A(n_581), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g757 ( .A1(n_630), .A2(n_188), .B(n_189), .C(n_191), .Y(n_757) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_632), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_569), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_555), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_597), .Y(n_761) );
NOR2xp67_ASAP7_75t_SL g762 ( .A(n_562), .B(n_193), .Y(n_762) );
INVx4_ASAP7_75t_L g763 ( .A(n_632), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_594), .A2(n_198), .B1(n_199), .B2(n_200), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_601), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_571), .A2(n_201), .B1(n_202), .B2(n_205), .C(n_206), .Y(n_766) );
BUFx2_ASAP7_75t_L g767 ( .A(n_611), .Y(n_767) );
AO31x2_ASAP7_75t_L g768 ( .A1(n_626), .A2(n_208), .A3(n_209), .B(n_210), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_635), .A2(n_212), .B1(n_214), .B2(n_215), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_584), .B(n_219), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_599), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_610), .A2(n_612), .B1(n_640), .B2(n_638), .Y(n_772) );
NOR2xp33_ASAP7_75t_SL g773 ( .A(n_561), .B(n_220), .Y(n_773) );
BUFx3_ASAP7_75t_L g774 ( .A(n_640), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_605), .B(n_222), .Y(n_775) );
CKINVDCx6p67_ASAP7_75t_R g776 ( .A(n_572), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_623), .Y(n_777) );
A2O1A1Ixp33_ASAP7_75t_L g778 ( .A1(n_627), .A2(n_229), .B(n_231), .C(n_233), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_624), .B(n_235), .Y(n_779) );
OAI21x1_ASAP7_75t_L g780 ( .A1(n_634), .A2(n_236), .B(n_636), .Y(n_780) );
OA21x2_ASAP7_75t_L g781 ( .A1(n_607), .A2(n_616), .B(n_622), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_614), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_688), .Y(n_783) );
A2O1A1Ixp33_ASAP7_75t_L g784 ( .A1(n_704), .A2(n_577), .B(n_600), .C(n_686), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_682), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_684), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_690), .Y(n_787) );
OR2x6_ASAP7_75t_L g788 ( .A(n_744), .B(n_600), .Y(n_788) );
AOI211xp5_ASAP7_75t_L g789 ( .A1(n_661), .A2(n_720), .B(n_727), .C(n_675), .Y(n_789) );
OAI21x1_ASAP7_75t_L g790 ( .A1(n_676), .A2(n_673), .B(n_679), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_688), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_725), .A2(n_761), .B1(n_736), .B2(n_705), .C(n_700), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_703), .A2(n_754), .B1(n_672), .B2(n_772), .Y(n_793) );
AOI21xp33_ASAP7_75t_L g794 ( .A1(n_734), .A2(n_708), .B(n_687), .Y(n_794) );
AND2x4_ASAP7_75t_L g795 ( .A(n_715), .B(n_685), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_668), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_681), .A2(n_662), .B(n_669), .C(n_729), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_678), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_693), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_774), .B(n_738), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_706), .B(n_702), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_669), .A2(n_711), .B1(n_744), .B2(n_662), .Y(n_802) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_696), .A2(n_677), .B1(n_689), .B2(n_718), .C(n_695), .Y(n_803) );
OAI22xp5_ASAP7_75t_SL g804 ( .A1(n_727), .A2(n_767), .B1(n_712), .B2(n_723), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_664), .B(n_760), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_659), .A2(n_663), .B(n_671), .Y(n_806) );
AO31x2_ASAP7_75t_L g807 ( .A1(n_670), .A2(n_737), .A3(n_713), .B(n_749), .Y(n_807) );
NAND2x1p5_ASAP7_75t_L g808 ( .A(n_680), .B(n_763), .Y(n_808) );
AOI21x1_ASAP7_75t_L g809 ( .A1(n_762), .A2(n_722), .B(n_683), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_759), .B(n_739), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_714), .B(n_771), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_741), .B(n_701), .Y(n_812) );
OR2x6_ASAP7_75t_L g813 ( .A(n_680), .B(n_753), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_728), .Y(n_814) );
A2O1A1Ixp33_ASAP7_75t_L g815 ( .A1(n_733), .A2(n_717), .B(n_707), .C(n_731), .Y(n_815) );
BUFx2_ASAP7_75t_L g816 ( .A(n_680), .Y(n_816) );
AOI222xp33_ASAP7_75t_SL g817 ( .A1(n_666), .A2(n_751), .B1(n_756), .B2(n_769), .C1(n_701), .C2(n_698), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_776), .B(n_716), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_775), .B(n_753), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_716), .B(n_692), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_773), .A2(n_726), .B(n_719), .Y(n_821) );
OAI21xp33_ASAP7_75t_L g822 ( .A1(n_711), .A2(n_773), .B(n_757), .Y(n_822) );
OAI21xp33_ASAP7_75t_L g823 ( .A1(n_764), .A2(n_747), .B(n_766), .Y(n_823) );
A2O1A1Ixp33_ASAP7_75t_L g824 ( .A1(n_745), .A2(n_732), .B(n_750), .C(n_755), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_730), .A2(n_709), .B(n_697), .Y(n_825) );
NAND2x1p5_ASAP7_75t_L g826 ( .A(n_763), .B(n_758), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_667), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_782), .B(n_777), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_765), .B(n_781), .Y(n_829) );
AND2x2_ASAP7_75t_SL g830 ( .A(n_751), .B(n_742), .Y(n_830) );
OA21x2_ASAP7_75t_L g831 ( .A1(n_699), .A2(n_721), .B(n_724), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_660), .Y(n_832) );
AOI221xp5_ASAP7_75t_SL g833 ( .A1(n_778), .A2(n_779), .B1(n_691), .B2(n_710), .C(n_743), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_781), .B(n_660), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_740), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_691), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_710), .A2(n_758), .B1(n_743), .B2(n_748), .Y(n_837) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_780), .A2(n_758), .B(n_743), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_735), .A2(n_740), .B(n_752), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_752), .A2(n_746), .B(n_768), .Y(n_840) );
OAI22xp5_ASAP7_75t_SL g841 ( .A1(n_746), .A2(n_568), .B1(n_495), .B2(n_419), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_768), .A2(n_770), .B(n_704), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_685), .Y(n_843) );
OR2x2_ASAP7_75t_L g844 ( .A(n_688), .B(n_478), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_682), .B(n_549), .Y(n_845) );
CKINVDCx16_ASAP7_75t_R g846 ( .A(n_738), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_674), .A2(n_575), .B(n_665), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_661), .A2(n_473), .B1(n_592), .B2(n_488), .C(n_460), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_688), .B(n_478), .Y(n_849) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_661), .A2(n_473), .B1(n_592), .B2(n_488), .C(n_460), .Y(n_850) );
AO31x2_ASAP7_75t_L g851 ( .A1(n_670), .A2(n_631), .A3(n_676), .B(n_737), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_661), .A2(n_495), .B1(n_473), .B2(n_568), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_682), .B(n_549), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_685), .Y(n_854) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_688), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_682), .B(n_549), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_688), .B(n_499), .Y(n_857) );
A2O1A1Ixp33_ASAP7_75t_L g858 ( .A1(n_704), .A2(n_686), .B(n_754), .C(n_560), .Y(n_858) );
A2O1A1Ixp33_ASAP7_75t_L g859 ( .A1(n_704), .A2(n_686), .B(n_754), .C(n_560), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_682), .B(n_549), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_682), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_770), .A2(n_704), .B(n_547), .Y(n_862) );
A2O1A1Ixp33_ASAP7_75t_L g863 ( .A1(n_704), .A2(n_686), .B(n_754), .C(n_560), .Y(n_863) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_704), .A2(n_550), .B(n_560), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_688), .B(n_478), .Y(n_865) );
OR2x2_ASAP7_75t_L g866 ( .A(n_688), .B(n_478), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_682), .B(n_549), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_682), .B(n_549), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_688), .B(n_499), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_682), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_669), .A2(n_501), .B1(n_510), .B2(n_435), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_661), .A2(n_495), .B1(n_473), .B2(n_568), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_682), .B(n_549), .Y(n_873) );
OR2x6_ASAP7_75t_L g874 ( .A(n_744), .B(n_668), .Y(n_874) );
AO21x2_ASAP7_75t_L g875 ( .A1(n_665), .A2(n_674), .B(n_694), .Y(n_875) );
AO21x2_ASAP7_75t_L g876 ( .A1(n_665), .A2(n_674), .B(n_694), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_688), .B(n_499), .Y(n_877) );
BUFx3_ASAP7_75t_L g878 ( .A(n_668), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_682), .B(n_549), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_661), .A2(n_495), .B1(n_473), .B2(n_568), .Y(n_880) );
CKINVDCx8_ASAP7_75t_R g881 ( .A(n_693), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_682), .B(n_549), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_669), .A2(n_501), .B1(n_510), .B2(n_435), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g884 ( .A1(n_704), .A2(n_560), .B(n_589), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_682), .B(n_549), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_688), .B(n_478), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_688), .B(n_478), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_669), .A2(n_501), .B1(n_510), .B2(n_435), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_682), .B(n_549), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_830), .B(n_857), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_843), .B(n_854), .Y(n_891) );
AND2x4_ASAP7_75t_L g892 ( .A(n_813), .B(n_812), .Y(n_892) );
OA21x2_ASAP7_75t_L g893 ( .A1(n_833), .A2(n_835), .B(n_842), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_829), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_785), .Y(n_895) );
NAND2x1_ASAP7_75t_L g896 ( .A(n_813), .B(n_788), .Y(n_896) );
BUFx5_ASAP7_75t_L g897 ( .A(n_832), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_786), .B(n_787), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_861), .B(n_870), .Y(n_899) );
AO21x2_ASAP7_75t_L g900 ( .A1(n_875), .A2(n_876), .B(n_784), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g901 ( .A1(n_852), .A2(n_872), .B1(n_880), .B2(n_850), .C(n_848), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_801), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_849), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_814), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_828), .Y(n_905) );
AO21x2_ASAP7_75t_L g906 ( .A1(n_797), .A2(n_822), .B(n_821), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_810), .B(n_864), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_884), .B(n_858), .Y(n_908) );
AOI21xp5_ASAP7_75t_SL g909 ( .A1(n_822), .A2(n_802), .B(n_859), .Y(n_909) );
AOI21xp5_ASAP7_75t_SL g910 ( .A1(n_863), .A2(n_788), .B(n_862), .Y(n_910) );
INVx3_ASAP7_75t_L g911 ( .A(n_826), .Y(n_911) );
AO21x1_ASAP7_75t_SL g912 ( .A1(n_818), .A2(n_819), .B(n_820), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_844), .B(n_866), .Y(n_913) );
AO21x2_ASAP7_75t_L g914 ( .A1(n_806), .A2(n_815), .B(n_837), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_865), .B(n_886), .Y(n_915) );
BUFx4f_ASAP7_75t_L g916 ( .A(n_874), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_845), .Y(n_917) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_887), .Y(n_918) );
AND2x4_ASAP7_75t_SL g919 ( .A(n_795), .B(n_783), .Y(n_919) );
AND2x4_ASAP7_75t_L g920 ( .A(n_836), .B(n_816), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_792), .B(n_889), .Y(n_921) );
OR2x2_ASAP7_75t_L g922 ( .A(n_791), .B(n_855), .Y(n_922) );
BUFx2_ASAP7_75t_L g923 ( .A(n_798), .Y(n_923) );
OA21x2_ASAP7_75t_L g924 ( .A1(n_825), .A2(n_824), .B(n_884), .Y(n_924) );
AND2x4_ASAP7_75t_L g925 ( .A(n_827), .B(n_809), .Y(n_925) );
AO21x2_ASAP7_75t_L g926 ( .A1(n_794), .A2(n_823), .B(n_803), .Y(n_926) );
AO21x1_ASAP7_75t_SL g927 ( .A1(n_817), .A2(n_853), .B(n_860), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_805), .B(n_873), .Y(n_928) );
OAI21xp5_ASAP7_75t_SL g929 ( .A1(n_888), .A2(n_793), .B(n_869), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_856), .B(n_885), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_867), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_868), .B(n_882), .Y(n_932) );
AOI322xp5_ASAP7_75t_L g933 ( .A1(n_877), .A2(n_846), .A3(n_879), .B1(n_795), .B2(n_841), .C1(n_811), .C2(n_878), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_831), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_808), .B(n_789), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_804), .B(n_800), .Y(n_936) );
INVx1_ASAP7_75t_SL g937 ( .A(n_796), .Y(n_937) );
AND2x4_ASAP7_75t_L g938 ( .A(n_807), .B(n_851), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_807), .B(n_851), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_851), .Y(n_940) );
INVxp67_ASAP7_75t_L g941 ( .A(n_874), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_817), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_874), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_881), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_799), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_829), .Y(n_946) );
OAI21x1_ASAP7_75t_L g947 ( .A1(n_847), .A2(n_838), .B(n_790), .Y(n_947) );
NOR2x1_ASAP7_75t_L g948 ( .A(n_788), .B(n_802), .Y(n_948) );
INVx3_ASAP7_75t_L g949 ( .A(n_826), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_849), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_834), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_844), .B(n_866), .Y(n_952) );
AND2x4_ASAP7_75t_L g953 ( .A(n_813), .B(n_812), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_829), .Y(n_954) );
AO21x2_ASAP7_75t_L g955 ( .A1(n_840), .A2(n_839), .B(n_835), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_829), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_871), .A2(n_501), .B1(n_510), .B2(n_883), .Y(n_957) );
AO21x2_ASAP7_75t_L g958 ( .A1(n_840), .A2(n_839), .B(n_835), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_904), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_934), .Y(n_960) );
OR2x2_ASAP7_75t_L g961 ( .A(n_894), .B(n_946), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_904), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_954), .B(n_956), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_942), .A2(n_901), .B1(n_957), .B2(n_927), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_942), .A2(n_927), .B1(n_936), .B2(n_948), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_908), .B(n_928), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_908), .B(n_907), .Y(n_967) );
OAI322xp33_ASAP7_75t_L g968 ( .A1(n_936), .A2(n_921), .A3(n_890), .B1(n_902), .B2(n_931), .C1(n_917), .C2(n_913), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_903), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_898), .B(n_899), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_898), .B(n_899), .Y(n_971) );
HB1xp67_ASAP7_75t_L g972 ( .A(n_951), .Y(n_972) );
BUFx2_ASAP7_75t_L g973 ( .A(n_897), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_917), .B(n_931), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g975 ( .A(n_937), .Y(n_975) );
BUFx2_ASAP7_75t_L g976 ( .A(n_897), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_939), .B(n_895), .Y(n_977) );
INVx2_ASAP7_75t_SL g978 ( .A(n_897), .Y(n_978) );
OR2x2_ASAP7_75t_L g979 ( .A(n_913), .B(n_952), .Y(n_979) );
INVxp67_ASAP7_75t_L g980 ( .A(n_912), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_891), .B(n_932), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_902), .B(n_926), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_948), .A2(n_935), .B1(n_953), .B2(n_892), .Y(n_983) );
OR2x2_ASAP7_75t_L g984 ( .A(n_922), .B(n_950), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_918), .B(n_915), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_932), .B(n_938), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_938), .B(n_892), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_938), .B(n_892), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_925), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_925), .Y(n_990) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_923), .Y(n_991) );
INVx2_ASAP7_75t_SL g992 ( .A(n_896), .Y(n_992) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_919), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_938), .B(n_892), .Y(n_994) );
NOR2x1_ASAP7_75t_L g995 ( .A(n_896), .B(n_926), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_953), .B(n_940), .Y(n_996) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_919), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_953), .B(n_925), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_926), .B(n_905), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_963), .B(n_933), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_963), .B(n_929), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_960), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_980), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1004 ( .A(n_968), .B(n_943), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_986), .B(n_958), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_977), .B(n_958), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_977), .B(n_958), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_959), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_968), .B(n_943), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_987), .B(n_955), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_996), .B(n_955), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_959), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_998), .B(n_906), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_964), .A2(n_916), .B1(n_912), .B2(n_914), .Y(n_1014) );
INVx4_ASAP7_75t_L g1015 ( .A(n_973), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_988), .B(n_906), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g1017 ( .A(n_972), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_994), .B(n_906), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_962), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_994), .B(n_900), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_984), .B(n_924), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_998), .B(n_947), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_970), .B(n_893), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_967), .B(n_941), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_965), .A2(n_930), .B1(n_905), .B2(n_944), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_967), .B(n_924), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_961), .B(n_909), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_974), .B(n_944), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_978), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1001), .B(n_970), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_1001), .B(n_971), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1002), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1008), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1028), .B(n_966), .Y(n_1034) );
NOR2xp33_ASAP7_75t_SL g1035 ( .A(n_1003), .B(n_975), .Y(n_1035) );
AND3x2_ASAP7_75t_L g1036 ( .A(n_1003), .B(n_997), .C(n_993), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1008), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1012), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1012), .Y(n_1039) );
OR2x6_ASAP7_75t_L g1040 ( .A(n_1015), .B(n_976), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1019), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_1021), .B(n_982), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_1021), .B(n_982), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_1023), .B(n_1005), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1028), .B(n_1000), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_1026), .B(n_979), .Y(n_1046) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_1026), .B(n_979), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1000), .B(n_981), .Y(n_1048) );
NOR2xp67_ASAP7_75t_L g1049 ( .A(n_1015), .B(n_978), .Y(n_1049) );
OR2x6_ASAP7_75t_L g1050 ( .A(n_1015), .B(n_978), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1023), .B(n_989), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_1006), .B(n_999), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_1005), .B(n_989), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1010), .B(n_990), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1010), .B(n_990), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_1017), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_1006), .B(n_999), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1044), .B(n_1016), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1033), .Y(n_1059) );
INVx3_ASAP7_75t_L g1060 ( .A(n_1050), .Y(n_1060) );
INVxp33_ASAP7_75t_L g1061 ( .A(n_1035), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_1052), .B(n_1007), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1045), .B(n_1007), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_1032), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1037), .Y(n_1065) );
NOR2xp67_ASAP7_75t_L g1066 ( .A(n_1049), .B(n_1029), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1038), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1032), .Y(n_1068) );
INVx1_ASAP7_75t_SL g1069 ( .A(n_1046), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1044), .B(n_1016), .Y(n_1070) );
AND2x4_ASAP7_75t_L g1071 ( .A(n_1050), .B(n_1022), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1030), .B(n_1004), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1031), .B(n_1009), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_1057), .B(n_1027), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1051), .B(n_1018), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1039), .Y(n_1076) );
AOI21xp33_ASAP7_75t_L g1077 ( .A1(n_1042), .A2(n_991), .B(n_1014), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1048), .B(n_944), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1041), .Y(n_1079) );
AND4x1_ASAP7_75t_L g1080 ( .A(n_1036), .B(n_945), .C(n_1025), .D(n_983), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1058), .B(n_1051), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1064), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1069), .B(n_1053), .Y(n_1083) );
NAND3xp33_ASAP7_75t_L g1084 ( .A(n_1080), .B(n_1056), .C(n_995), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1072), .B(n_1054), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1073), .B(n_1054), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1074), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_1061), .A2(n_1050), .B1(n_1040), .B2(n_1047), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1058), .B(n_1055), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1063), .B(n_1034), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1064), .Y(n_1091) );
AOI21xp33_ASAP7_75t_L g1092 ( .A1(n_1078), .A2(n_969), .B(n_985), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1068), .Y(n_1093) );
A2O1A1Ixp33_ASAP7_75t_L g1094 ( .A1(n_1088), .A2(n_1066), .B(n_1060), .C(n_1071), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1089), .B(n_1070), .Y(n_1095) );
NAND2xp5_ASAP7_75t_SL g1096 ( .A(n_1084), .B(n_1066), .Y(n_1096) );
O2A1O1Ixp5_ASAP7_75t_L g1097 ( .A1(n_1092), .A2(n_1060), .B(n_1077), .C(n_1071), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1087), .Y(n_1098) );
AOI221x1_ASAP7_75t_L g1099 ( .A1(n_1091), .A2(n_945), .B1(n_1067), .B2(n_1065), .C(n_1059), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_1097), .A2(n_1090), .B1(n_1085), .B2(n_1086), .C(n_1083), .Y(n_1100) );
AOI211xp5_ASAP7_75t_L g1101 ( .A1(n_1094), .A2(n_1024), .B(n_910), .C(n_1047), .Y(n_1101) );
OAI21xp33_ASAP7_75t_L g1102 ( .A1(n_1094), .A2(n_1062), .B(n_1089), .Y(n_1102) );
NOR2xp67_ASAP7_75t_L g1103 ( .A(n_1096), .B(n_1081), .Y(n_1103) );
AOI322xp5_ASAP7_75t_L g1104 ( .A1(n_1102), .A2(n_1095), .A3(n_1098), .B1(n_1075), .B2(n_1093), .C1(n_1020), .C2(n_1011), .Y(n_1104) );
NAND4xp25_ASAP7_75t_L g1105 ( .A(n_1101), .B(n_1099), .C(n_910), .D(n_974), .Y(n_1105) );
NAND2xp5_ASAP7_75t_SL g1106 ( .A(n_1103), .B(n_1100), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1106), .Y(n_1107) );
NOR3xp33_ASAP7_75t_L g1108 ( .A(n_1105), .B(n_911), .C(n_949), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1107), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1108), .B(n_1104), .Y(n_1110) );
INVx3_ASAP7_75t_SL g1111 ( .A(n_1109), .Y(n_1111) );
AND2x2_ASAP7_75t_SL g1112 ( .A(n_1109), .B(n_1110), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1111), .Y(n_1113) );
AOI22x1_ASAP7_75t_L g1114 ( .A1(n_1112), .A2(n_1110), .B1(n_1082), .B2(n_992), .Y(n_1114) );
AO21x1_ASAP7_75t_L g1115 ( .A1(n_1113), .A2(n_1079), .B(n_1065), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_1115), .A2(n_1114), .B1(n_1067), .B2(n_1076), .Y(n_1116) );
XOR2xp5_ASAP7_75t_L g1117 ( .A(n_1116), .B(n_920), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_1117), .A2(n_1022), .B1(n_1013), .B2(n_1043), .Y(n_1118) );
endmodule