module fake_jpeg_20083_n_140 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_1),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_14),
.C(n_16),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_37),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_25),
.B1(n_13),
.B2(n_29),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_38),
.B1(n_34),
.B2(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_29),
.B1(n_27),
.B2(n_13),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_51),
.B1(n_22),
.B2(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_38),
.B1(n_34),
.B2(n_35),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_24),
.C(n_23),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_60),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_24),
.C(n_23),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_14),
.B1(n_17),
.B2(n_12),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_10),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_73),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_12),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_67),
.C(n_61),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_86),
.C(n_82),
.Y(n_105)
);

NOR4xp25_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_67),
.C(n_18),
.D(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_81),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_67),
.B(n_51),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.C(n_57),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_61),
.B(n_19),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_57),
.B(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_103),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_106),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_83),
.B1(n_76),
.B2(n_74),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_94),
.B1(n_92),
.B2(n_16),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_91),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_107),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_107),
.B(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_101),
.C(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_21),
.B1(n_16),
.B2(n_5),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_122),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_109),
.B(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_2),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_21),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_107),
.B(n_7),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_113),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_120),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_21),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_3),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_9),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_127),
.B(n_125),
.C(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_133),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.C(n_135),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_5),
.B(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);


endmodule