module real_aes_11202_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_892;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_1584;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g1544 ( .A(n_0), .Y(n_1544) );
OAI22xp5_ASAP7_75t_L g1574 ( .A1(n_0), .A2(n_186), .B1(n_296), .B2(n_349), .Y(n_1574) );
INVx1_ASAP7_75t_L g815 ( .A(n_1), .Y(n_815) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_2), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_2), .A2(n_51), .B1(n_635), .B2(n_638), .Y(n_634) );
INVxp33_ASAP7_75t_L g808 ( .A(n_3), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_3), .A2(n_785), .B(n_847), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_4), .A2(n_190), .B1(n_574), .B2(n_578), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_4), .A2(n_190), .B1(n_694), .B2(n_695), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_5), .A2(n_124), .B1(n_535), .B2(n_685), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_5), .A2(n_124), .B1(n_694), .B2(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g336 ( .A(n_6), .Y(n_336) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_7), .Y(n_295) );
INVx1_ASAP7_75t_L g469 ( .A(n_7), .Y(n_469) );
AND2x2_ASAP7_75t_L g822 ( .A(n_7), .B(n_314), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_7), .B(n_210), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_8), .A2(n_74), .B1(n_1182), .B2(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1452 ( .A(n_9), .Y(n_1452) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_9), .A2(n_91), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
INVx1_ASAP7_75t_L g812 ( .A(n_10), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_11), .A2(n_101), .B1(n_425), .B2(n_1073), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_11), .A2(n_101), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
OAI21xp33_ASAP7_75t_SL g479 ( .A1(n_12), .A2(n_480), .B(n_486), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_12), .A2(n_139), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_13), .A2(n_43), .B1(n_688), .B2(n_1127), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_13), .A2(n_43), .B1(n_385), .B2(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g817 ( .A(n_14), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_14), .A2(n_280), .B1(n_830), .B2(n_837), .C(n_839), .Y(n_829) );
INVx1_ASAP7_75t_L g1099 ( .A(n_15), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g1439 ( .A1(n_16), .A2(n_238), .B1(n_1440), .B2(n_1445), .C(n_1448), .Y(n_1439) );
OAI22xp33_ASAP7_75t_L g1486 ( .A1(n_16), .A2(n_238), .B1(n_1487), .B2(n_1490), .Y(n_1486) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_17), .A2(n_216), .B1(n_613), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_17), .A2(n_216), .B1(n_631), .B2(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_18), .A2(n_273), .B1(n_696), .B2(n_934), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_18), .A2(n_273), .B1(n_574), .B2(n_578), .Y(n_981) );
INVx1_ASAP7_75t_L g490 ( .A(n_19), .Y(n_490) );
OAI222xp33_ASAP7_75t_L g502 ( .A1(n_19), .A2(n_24), .B1(n_271), .B2(n_503), .C1(n_504), .C2(n_507), .Y(n_502) );
XNOR2xp5_ASAP7_75t_L g1526 ( .A(n_20), .B(n_1527), .Y(n_1526) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_21), .A2(n_81), .B1(n_1182), .B2(n_1207), .Y(n_1211) );
INVx1_ASAP7_75t_L g1453 ( .A(n_22), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1503 ( .A1(n_22), .A2(n_252), .B1(n_1504), .B2(n_1506), .C(n_1508), .Y(n_1503) );
INVx1_ASAP7_75t_L g568 ( .A(n_23), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_24), .A2(n_188), .B1(n_544), .B2(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g363 ( .A(n_25), .Y(n_363) );
OR2x2_ASAP7_75t_L g1485 ( .A(n_25), .B(n_1479), .Y(n_1485) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_26), .A2(n_90), .B1(n_532), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_26), .A2(n_90), .B1(n_549), .B2(n_554), .Y(n_793) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_27), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_27), .A2(n_268), .B1(n_866), .B2(n_876), .Y(n_875) );
INVxp33_ASAP7_75t_L g893 ( .A(n_28), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_28), .A2(n_244), .B1(n_922), .B2(n_937), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g1210 ( .A1(n_29), .A2(n_144), .B1(n_1197), .B2(n_1203), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_30), .A2(n_243), .B1(n_710), .B2(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_30), .Y(n_745) );
INVx1_ASAP7_75t_L g1059 ( .A(n_31), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_31), .A2(n_128), .B1(n_866), .B2(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_32), .A2(n_206), .B1(n_726), .B2(n_727), .Y(n_725) );
OAI211xp5_ASAP7_75t_SL g731 ( .A1(n_32), .A2(n_350), .B(n_732), .C(n_735), .Y(n_731) );
BUFx2_ASAP7_75t_L g355 ( .A(n_33), .Y(n_355) );
BUFx2_ASAP7_75t_L g408 ( .A(n_33), .Y(n_408) );
INVx1_ASAP7_75t_L g467 ( .A(n_33), .Y(n_467) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_33), .B(n_836), .Y(n_1444) );
INVx1_ASAP7_75t_L g1000 ( .A(n_34), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_34), .A2(n_231), .B1(n_687), .B2(n_978), .Y(n_1017) );
INVx1_ASAP7_75t_L g1052 ( .A(n_35), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_35), .A2(n_106), .B1(n_953), .B2(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1243 ( .A(n_36), .Y(n_1243) );
CKINVDCx5p33_ASAP7_75t_R g1536 ( .A(n_37), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_38), .A2(n_58), .B1(n_1025), .B2(n_1548), .Y(n_1547) );
OAI211xp5_ASAP7_75t_L g1575 ( .A1(n_38), .A2(n_350), .B(n_1576), .C(n_1579), .Y(n_1575) );
INVx1_ASAP7_75t_L g1065 ( .A(n_39), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_39), .A2(n_54), .B1(n_425), .B2(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g492 ( .A(n_40), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_40), .A2(n_188), .B1(n_296), .B2(n_349), .Y(n_501) );
INVx1_ASAP7_75t_L g1102 ( .A(n_41), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_41), .A2(n_104), .B1(n_613), .B2(n_1122), .Y(n_1121) );
INVxp33_ASAP7_75t_L g810 ( .A(n_42), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_42), .A2(n_102), .B1(n_535), .B2(n_677), .C(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g1104 ( .A(n_44), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_44), .A2(n_166), .B1(n_1110), .B2(n_1111), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_45), .A2(n_194), .B1(n_611), .B2(n_613), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_45), .A2(n_194), .B1(n_432), .B2(n_718), .Y(n_717) );
INVxp33_ASAP7_75t_L g1154 ( .A(n_46), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_46), .A2(n_171), .B1(n_677), .B2(n_827), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_47), .A2(n_59), .B1(n_685), .B2(n_1125), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_47), .A2(n_59), .B1(n_626), .B2(n_724), .Y(n_1132) );
INVxp33_ASAP7_75t_SL g754 ( .A(n_48), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_48), .A2(n_57), .B1(n_799), .B2(n_800), .Y(n_798) );
AO22x2_ASAP7_75t_L g1040 ( .A1(n_49), .A2(n_1041), .B1(n_1042), .B2(n_1086), .Y(n_1040) );
INVx1_ASAP7_75t_L g1086 ( .A(n_49), .Y(n_1086) );
INVx1_ASAP7_75t_L g771 ( .A(n_50), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_50), .A2(n_189), .B1(n_778), .B2(n_784), .Y(n_783) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_51), .Y(n_609) );
INVx1_ASAP7_75t_L g902 ( .A(n_52), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_52), .A2(n_161), .B1(n_911), .B2(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_53), .A2(n_264), .B1(n_611), .B2(n_613), .Y(n_610) );
AOI221xp5_ASAP7_75t_SL g629 ( .A1(n_53), .A2(n_412), .B1(n_630), .B2(n_632), .C(n_640), .Y(n_629) );
INVx1_ASAP7_75t_L g1061 ( .A(n_54), .Y(n_1061) );
INVx1_ASAP7_75t_L g1428 ( .A(n_55), .Y(n_1428) );
AOI221xp5_ASAP7_75t_L g1492 ( .A1(n_55), .A2(n_143), .B1(n_925), .B2(n_928), .C(n_1493), .Y(n_1492) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_56), .A2(n_564), .B(n_566), .C(n_567), .Y(n_563) );
INVx1_ASAP7_75t_L g598 ( .A(n_56), .Y(n_598) );
INVxp33_ASAP7_75t_SL g755 ( .A(n_57), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g1582 ( .A1(n_58), .A2(n_120), .B1(n_574), .B2(n_578), .Y(n_1582) );
XNOR2xp5_ASAP7_75t_L g650 ( .A(n_60), .B(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_60), .A2(n_112), .B1(n_1197), .B2(n_1203), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_61), .A2(n_162), .B1(n_613), .B2(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_61), .A2(n_162), .B1(n_727), .B2(n_922), .Y(n_921) );
INVxp33_ASAP7_75t_SL g762 ( .A(n_62), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_62), .A2(n_63), .B1(n_425), .B2(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g757 ( .A(n_63), .Y(n_757) );
INVx1_ASAP7_75t_L g1051 ( .A(n_64), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g1080 ( .A1(n_64), .A2(n_85), .B1(n_784), .B2(n_1081), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g993 ( .A(n_65), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_66), .A2(n_70), .B1(n_417), .B2(n_419), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_66), .A2(n_70), .B1(n_451), .B2(n_454), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_67), .A2(n_237), .B1(n_613), .B2(n_682), .Y(n_715) );
INVx1_ASAP7_75t_L g742 ( .A(n_67), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_68), .A2(n_93), .B1(n_495), .B2(n_561), .Y(n_943) );
INVx1_ASAP7_75t_L g961 ( .A(n_68), .Y(n_961) );
INVxp33_ASAP7_75t_L g1148 ( .A(n_69), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_69), .A2(n_100), .B1(n_385), .B2(n_432), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g1469 ( .A(n_71), .Y(n_1469) );
INVxp33_ASAP7_75t_SL g767 ( .A(n_72), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_72), .A2(n_156), .B1(n_532), .B2(n_781), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g950 ( .A1(n_73), .A2(n_260), .B1(n_498), .B2(n_562), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_73), .A2(n_260), .B1(n_451), .B2(n_915), .C(n_960), .Y(n_959) );
AOI222xp33_ASAP7_75t_L g1420 ( .A1(n_74), .A2(n_1421), .B1(n_1523), .B2(n_1525), .C1(n_1588), .C2(n_1590), .Y(n_1420) );
AOI22xp5_ASAP7_75t_L g1423 ( .A1(n_74), .A2(n_1424), .B1(n_1521), .B2(n_1522), .Y(n_1423) );
INVx1_ASAP7_75t_L g1521 ( .A(n_74), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_75), .A2(n_219), .B1(n_516), .B2(n_520), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_75), .A2(n_239), .B1(n_542), .B2(n_544), .Y(n_541) );
INVx1_ASAP7_75t_L g1572 ( .A(n_76), .Y(n_1572) );
OAI211xp5_ASAP7_75t_SL g1586 ( .A1(n_76), .A2(n_358), .B(n_621), .C(n_1587), .Y(n_1586) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_77), .A2(n_129), .B1(n_1197), .B2(n_1203), .Y(n_1220) );
INVx1_ASAP7_75t_L g660 ( .A(n_78), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_79), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_79), .A2(n_141), .B1(n_535), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_80), .A2(n_254), .B1(n_451), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_80), .A2(n_254), .B1(n_925), .B2(n_928), .Y(n_924) );
INVx1_ASAP7_75t_L g1145 ( .A(n_82), .Y(n_1145) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_83), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_83), .A2(n_167), .B1(n_419), .B2(n_866), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g1010 ( .A1(n_84), .A2(n_278), .B1(n_460), .B2(n_710), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_84), .A2(n_278), .B1(n_418), .B2(n_720), .Y(n_1021) );
OAI222xp33_ASAP7_75t_L g1045 ( .A1(n_85), .A2(n_173), .B1(n_266), .B2(n_1046), .C1(n_1047), .C2(n_1049), .Y(n_1045) );
INVx1_ASAP7_75t_L g891 ( .A(n_86), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g1580 ( .A(n_87), .Y(n_1580) );
INVxp33_ASAP7_75t_SL g375 ( .A(n_88), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_88), .A2(n_259), .B1(n_459), .B2(n_461), .Y(n_458) );
AO22x2_ASAP7_75t_L g1137 ( .A1(n_89), .A2(n_1138), .B1(n_1173), .B2(n_1174), .Y(n_1137) );
INVx1_ASAP7_75t_L g1173 ( .A(n_89), .Y(n_1173) );
INVx1_ASAP7_75t_L g1459 ( .A(n_91), .Y(n_1459) );
INVxp33_ASAP7_75t_SL g1097 ( .A(n_92), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_92), .A2(n_178), .B1(n_535), .B2(n_685), .Y(n_1120) );
INVx1_ASAP7_75t_L g980 ( .A(n_93), .Y(n_980) );
AO22x2_ASAP7_75t_L g985 ( .A1(n_94), .A2(n_986), .B1(n_1028), .B2(n_1029), .Y(n_985) );
INVxp67_ASAP7_75t_L g1028 ( .A(n_94), .Y(n_1028) );
INVx1_ASAP7_75t_L g748 ( .A(n_95), .Y(n_748) );
INVx1_ASAP7_75t_L g406 ( .A(n_96), .Y(n_406) );
INVx1_ASAP7_75t_L g1479 ( .A(n_96), .Y(n_1479) );
INVx1_ASAP7_75t_L g737 ( .A(n_97), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_98), .A2(n_174), .B1(n_424), .B2(n_427), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_98), .A2(n_174), .B1(n_328), .B2(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_99), .A2(n_114), .B1(n_531), .B2(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_99), .A2(n_114), .B1(n_788), .B2(n_791), .Y(n_787) );
INVx1_ASAP7_75t_L g1144 ( .A(n_100), .Y(n_1144) );
INVxp67_ASAP7_75t_SL g813 ( .A(n_102), .Y(n_813) );
INVx1_ASAP7_75t_L g955 ( .A(n_103), .Y(n_955) );
INVxp33_ASAP7_75t_SL g1096 ( .A(n_104), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g1435 ( .A(n_105), .Y(n_1435) );
INVx1_ASAP7_75t_L g1055 ( .A(n_106), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_107), .A2(n_132), .B1(n_1197), .B2(n_1203), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_108), .A2(n_224), .B1(n_1197), .B2(n_1203), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_109), .A2(n_158), .B1(n_418), .B2(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_109), .A2(n_158), .B1(n_574), .B2(n_578), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_110), .A2(n_127), .B1(n_315), .B2(n_680), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_110), .A2(n_127), .B1(n_419), .B2(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g989 ( .A(n_111), .Y(n_989) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_111), .A2(n_245), .B1(n_934), .B2(n_935), .Y(n_1027) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_113), .A2(n_147), .B1(n_1182), .B2(n_1207), .Y(n_1206) );
CKINVDCx5p33_ASAP7_75t_R g1581 ( .A(n_115), .Y(n_1581) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_116), .A2(n_152), .B1(n_1071), .B2(n_1075), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_116), .A2(n_152), .B1(n_524), .B2(n_526), .Y(n_1082) );
INVx1_ASAP7_75t_L g1226 ( .A(n_117), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_118), .A2(n_220), .B1(n_682), .B2(n_1012), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_118), .A2(n_220), .B1(n_428), .B2(n_631), .Y(n_1020) );
CKINVDCx5p33_ASAP7_75t_R g1432 ( .A(n_119), .Y(n_1432) );
INVx1_ASAP7_75t_L g1546 ( .A(n_120), .Y(n_1546) );
INVxp33_ASAP7_75t_SL g319 ( .A(n_121), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_121), .A2(n_258), .B1(n_417), .B2(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g758 ( .A(n_122), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_123), .A2(n_146), .B1(n_495), .B2(n_498), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_123), .A2(n_146), .B1(n_531), .B2(n_532), .Y(n_530) );
OAI211xp5_ASAP7_75t_L g579 ( .A1(n_125), .A2(n_350), .B(n_580), .C(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g624 ( .A(n_125), .Y(n_624) );
INVx1_ASAP7_75t_L g1568 ( .A(n_126), .Y(n_1568) );
OAI22xp5_ASAP7_75t_L g1584 ( .A1(n_126), .A2(n_150), .B1(n_495), .B2(n_498), .Y(n_1584) );
INVx1_ASAP7_75t_L g1058 ( .A(n_128), .Y(n_1058) );
INVx1_ASAP7_75t_L g287 ( .A(n_130), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_131), .A2(n_195), .B1(n_495), .B2(n_498), .Y(n_570) );
INVx1_ASAP7_75t_L g588 ( .A(n_131), .Y(n_588) );
AO22x1_ASAP7_75t_SL g1223 ( .A1(n_133), .A2(n_230), .B1(n_1197), .B2(n_1203), .Y(n_1223) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_134), .A2(n_218), .B1(n_459), .B2(n_953), .C(n_954), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_134), .A2(n_218), .B1(n_934), .B2(n_935), .Y(n_969) );
INVx1_ASAP7_75t_L g949 ( .A(n_135), .Y(n_949) );
INVx1_ASAP7_75t_L g1266 ( .A(n_136), .Y(n_1266) );
AO221x2_ASAP7_75t_L g1237 ( .A1(n_137), .A2(n_267), .B1(n_1218), .B2(n_1238), .C(n_1239), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_138), .A2(n_206), .B1(n_296), .B2(n_349), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_138), .A2(n_237), .B1(n_495), .B2(n_561), .Y(n_747) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_139), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_140), .Y(n_997) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_141), .Y(n_662) );
CKINVDCx5p33_ASAP7_75t_R g1461 ( .A(n_142), .Y(n_1461) );
INVx1_ASAP7_75t_L g1437 ( .A(n_143), .Y(n_1437) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_145), .A2(n_183), .B1(n_1538), .B2(n_1540), .Y(n_1537) );
INVx1_ASAP7_75t_L g1554 ( .A(n_145), .Y(n_1554) );
CKINVDCx5p33_ASAP7_75t_R g1468 ( .A(n_148), .Y(n_1468) );
INVx1_ASAP7_75t_L g882 ( .A(n_149), .Y(n_882) );
INVx1_ASAP7_75t_L g1565 ( .A(n_150), .Y(n_1565) );
CKINVDCx14_ASAP7_75t_R g940 ( .A(n_151), .Y(n_940) );
INVx1_ASAP7_75t_L g948 ( .A(n_153), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_154), .A2(n_239), .B1(n_524), .B2(n_526), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_154), .A2(n_219), .B1(n_547), .B2(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g1149 ( .A(n_155), .Y(n_1149) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_156), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_157), .A2(n_165), .B1(n_594), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_157), .A2(n_165), .B1(n_694), .B2(n_720), .Y(n_719) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_159), .A2(n_202), .B1(n_495), .B2(n_561), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_159), .A2(n_236), .B1(n_687), .B2(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g759 ( .A(n_160), .Y(n_759) );
INVxp33_ASAP7_75t_L g897 ( .A(n_161), .Y(n_897) );
INVxp33_ASAP7_75t_L g1142 ( .A(n_163), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_163), .A2(n_170), .B1(n_694), .B2(n_724), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1234 ( .A1(n_164), .A2(n_265), .B1(n_1182), .B2(n_1207), .Y(n_1234) );
INVx1_ASAP7_75t_L g1103 ( .A(n_166), .Y(n_1103) );
INVxp33_ASAP7_75t_L g1113 ( .A(n_167), .Y(n_1113) );
INVx1_ASAP7_75t_L g1146 ( .A(n_168), .Y(n_1146) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_169), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_169), .A2(n_213), .B1(n_914), .B2(n_915), .Y(n_913) );
INVxp33_ASAP7_75t_L g1141 ( .A(n_170), .Y(n_1141) );
INVxp33_ASAP7_75t_L g1156 ( .A(n_171), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_172), .A2(n_241), .B1(n_613), .B2(n_1122), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_172), .A2(n_241), .B1(n_718), .B2(n_1024), .Y(n_1166) );
INVx1_ASAP7_75t_L g1062 ( .A(n_173), .Y(n_1062) );
INVx1_ASAP7_75t_L g886 ( .A(n_175), .Y(n_886) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_176), .Y(n_289) );
AND3x2_ASAP7_75t_L g1185 ( .A(n_176), .B(n_287), .C(n_1186), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_176), .B(n_287), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_177), .A2(n_235), .B1(n_561), .B2(n_562), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_177), .A2(n_207), .B1(n_296), .B2(n_349), .Y(n_584) );
INVxp33_ASAP7_75t_SL g1100 ( .A(n_178), .Y(n_1100) );
INVxp33_ASAP7_75t_SL g1116 ( .A(n_179), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_179), .A2(n_246), .B1(n_385), .B2(n_1131), .Y(n_1134) );
INVxp33_ASAP7_75t_L g1157 ( .A(n_180), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_180), .A2(n_187), .B1(n_613), .B2(n_682), .Y(n_1164) );
INVx1_ASAP7_75t_L g658 ( .A(n_181), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_182), .A2(n_251), .B1(n_1182), .B2(n_1218), .Y(n_1221) );
INVx1_ASAP7_75t_L g1559 ( .A(n_183), .Y(n_1559) );
INVx2_ASAP7_75t_L g300 ( .A(n_184), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_185), .A2(n_751), .B1(n_802), .B2(n_803), .Y(n_750) );
INVxp67_ASAP7_75t_L g802 ( .A(n_185), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g1585 ( .A1(n_186), .A2(n_249), .B1(n_561), .B2(n_562), .Y(n_1585) );
INVx1_ASAP7_75t_L g1152 ( .A(n_187), .Y(n_1152) );
INVxp33_ASAP7_75t_SL g766 ( .A(n_189), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_191), .A2(n_211), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_191), .A2(n_211), .B1(n_694), .B2(n_695), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g1480 ( .A(n_192), .Y(n_1480) );
INVx1_ASAP7_75t_L g1227 ( .A(n_193), .Y(n_1227) );
INVx1_ASAP7_75t_L g596 ( .A(n_195), .Y(n_596) );
AOI21xp33_ASAP7_75t_L g840 ( .A1(n_196), .A2(n_538), .B(n_841), .Y(n_840) );
INVxp67_ASAP7_75t_SL g864 ( .A(n_196), .Y(n_864) );
INVx1_ASAP7_75t_L g1186 ( .A(n_197), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g887 ( .A(n_198), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_198), .A2(n_234), .B1(n_932), .B2(n_935), .Y(n_931) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_199), .A2(n_350), .B(n_669), .C(n_670), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_199), .A2(n_279), .B1(n_692), .B2(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g854 ( .A(n_200), .Y(n_854) );
INVx1_ASAP7_75t_L g763 ( .A(n_201), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_202), .A2(n_279), .B1(n_296), .B2(n_349), .Y(n_673) );
INVxp33_ASAP7_75t_SL g510 ( .A(n_203), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_203), .A2(n_261), .B1(n_549), .B2(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g1006 ( .A(n_204), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_204), .A2(n_250), .B1(n_685), .B2(n_1016), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_205), .A2(n_270), .B1(n_574), .B2(n_578), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_205), .A2(n_270), .B1(n_626), .B2(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g620 ( .A(n_207), .Y(n_620) );
INVx1_ASAP7_75t_L g971 ( .A(n_208), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g1240 ( .A(n_209), .Y(n_1240) );
INVx1_ASAP7_75t_L g302 ( .A(n_210), .Y(n_302) );
INVx2_ASAP7_75t_L g314 ( .A(n_210), .Y(n_314) );
OAI211xp5_ASAP7_75t_L g944 ( .A1(n_212), .A2(n_566), .B(n_945), .C(n_947), .Y(n_944) );
INVx1_ASAP7_75t_L g964 ( .A(n_212), .Y(n_964) );
INVxp67_ASAP7_75t_SL g900 ( .A(n_213), .Y(n_900) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_214), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_214), .A2(n_262), .B1(n_445), .B2(n_451), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g804 ( .A(n_215), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g992 ( .A(n_217), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_217), .A2(n_276), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
OAI211xp5_ASAP7_75t_L g1032 ( .A1(n_217), .A2(n_350), .B(n_580), .C(n_1033), .Y(n_1032) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_221), .Y(n_889) );
INVx1_ASAP7_75t_L g852 ( .A(n_222), .Y(n_852) );
INVx1_ASAP7_75t_L g957 ( .A(n_223), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_225), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_226), .A2(n_227), .B1(n_1180), .B2(n_1264), .C(n_1265), .Y(n_1263) );
INVx1_ASAP7_75t_L g347 ( .A(n_228), .Y(n_347) );
INVx1_ASAP7_75t_L g569 ( .A(n_229), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_230), .A2(n_558), .B1(n_642), .B2(n_643), .Y(n_557) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_230), .Y(n_643) );
INVx1_ASAP7_75t_L g1004 ( .A(n_231), .Y(n_1004) );
OAI211xp5_ASAP7_75t_L g1037 ( .A1(n_231), .A2(n_564), .B(n_566), .C(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g327 ( .A(n_232), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_232), .A2(n_256), .B1(n_384), .B2(n_419), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g1534 ( .A(n_233), .Y(n_1534) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_234), .Y(n_894) );
INVx1_ASAP7_75t_L g592 ( .A(n_235), .Y(n_592) );
INVx1_ASAP7_75t_L g655 ( .A(n_236), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g1465 ( .A(n_240), .Y(n_1465) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_242), .A2(n_307), .B1(n_308), .B2(n_470), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_242), .Y(n_307) );
INVx1_ASAP7_75t_L g746 ( .A(n_243), .Y(n_746) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_244), .Y(n_890) );
INVx1_ASAP7_75t_L g990 ( .A(n_245), .Y(n_990) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_246), .Y(n_1108) );
XOR2x2_ASAP7_75t_L g1092 ( .A(n_247), .B(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1184 ( .A(n_248), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_248), .B(n_1200), .Y(n_1205) );
INVx1_ASAP7_75t_L g1571 ( .A(n_249), .Y(n_1571) );
INVx1_ASAP7_75t_L g1001 ( .A(n_250), .Y(n_1001) );
INVx1_ASAP7_75t_L g1455 ( .A(n_252), .Y(n_1455) );
INVx1_ASAP7_75t_L g736 ( .A(n_253), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_255), .Y(n_994) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_256), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_257), .Y(n_842) );
INVxp33_ASAP7_75t_SL g345 ( .A(n_258), .Y(n_345) );
INVx1_ASAP7_75t_L g383 ( .A(n_259), .Y(n_383) );
INVxp33_ASAP7_75t_L g509 ( .A(n_261), .Y(n_509) );
INVxp33_ASAP7_75t_SL g395 ( .A(n_262), .Y(n_395) );
INVx2_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_264), .Y(n_633) );
INVx1_ASAP7_75t_L g1063 ( .A(n_266), .Y(n_1063) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_268), .Y(n_820) );
XOR2xp5_ASAP7_75t_L g474 ( .A(n_269), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g487 ( .A(n_271), .Y(n_487) );
INVx1_ASAP7_75t_L g333 ( .A(n_272), .Y(n_333) );
BUFx3_ASAP7_75t_L g366 ( .A(n_274), .Y(n_366) );
INVx1_ASAP7_75t_L g381 ( .A(n_274), .Y(n_381) );
BUFx3_ASAP7_75t_L g367 ( .A(n_275), .Y(n_367) );
INVx1_ASAP7_75t_L g403 ( .A(n_275), .Y(n_403) );
INVx1_ASAP7_75t_L g996 ( .A(n_276), .Y(n_996) );
INVx1_ASAP7_75t_L g972 ( .A(n_277), .Y(n_972) );
INVx1_ASAP7_75t_L g816 ( .A(n_280), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_303), .B(n_1178), .Y(n_281) );
INVx3_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x4_ASAP7_75t_L g1524 ( .A(n_285), .B(n_291), .Y(n_1524) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g1589 ( .A(n_286), .Y(n_1589) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_286), .B(n_288), .Y(n_1595) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_288), .B(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x6_ASAP7_75t_L g354 ( .A(n_293), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g512 ( .A(n_293), .B(n_355), .Y(n_512) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g443 ( .A(n_294), .B(n_302), .Y(n_443) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g615 ( .A(n_295), .B(n_313), .Y(n_615) );
INVx8_ASAP7_75t_L g346 ( .A(n_296), .Y(n_346) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
OR2x6_ASAP7_75t_L g349 ( .A(n_297), .B(n_312), .Y(n_349) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_297), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g841 ( .A1(n_297), .A2(n_443), .B(n_842), .Y(n_841) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_297), .Y(n_956) );
INVx2_ASAP7_75t_SL g963 ( .A(n_297), .Y(n_963) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_297), .B(n_1444), .Y(n_1473) );
INVx2_ASAP7_75t_SL g1562 ( .A(n_297), .Y(n_1562) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
AND2x4_ASAP7_75t_L g323 ( .A(n_299), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g332 ( .A(n_299), .Y(n_332) );
INVx1_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
AND2x2_ASAP7_75t_L g449 ( .A(n_299), .B(n_300), .Y(n_449) );
INVx1_ASAP7_75t_L g318 ( .A(n_300), .Y(n_318) );
INVx2_ASAP7_75t_L g324 ( .A(n_300), .Y(n_324) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
INVx1_ASAP7_75t_L g506 ( .A(n_300), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_300), .B(n_316), .Y(n_577) );
AND2x4_ASAP7_75t_L g334 ( .A(n_301), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g507 ( .A(n_302), .B(n_339), .Y(n_507) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_302), .B(n_339), .Y(n_1111) );
XNOR2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_982), .Y(n_303) );
XOR2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_647), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_471), .B1(n_472), .B2(n_646), .Y(n_305) );
INVx2_ASAP7_75t_SL g646 ( .A(n_306), .Y(n_646) );
INVx1_ASAP7_75t_L g470 ( .A(n_308), .Y(n_470) );
AOI221x1_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_353), .B1(n_356), .B2(n_404), .C(n_409), .Y(n_308) );
NAND4xp25_ASAP7_75t_L g309 ( .A(n_310), .B(n_326), .C(n_344), .D(n_350), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_319), .B1(n_320), .B2(n_325), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_311), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_311), .A2(n_320), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_311), .A2(n_348), .B1(n_886), .B2(n_887), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g988 ( .A1(n_311), .A2(n_320), .B1(n_989), .B2(n_990), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_311), .A2(n_320), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_311), .A2(n_511), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_311), .A2(n_511), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
AND2x4_ASAP7_75t_L g320 ( .A(n_312), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g511 ( .A(n_312), .B(n_321), .Y(n_511) );
INVx1_ASAP7_75t_L g575 ( .A(n_312), .Y(n_575) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_315), .Y(n_453) );
INVx1_ASAP7_75t_L g525 ( .A(n_315), .Y(n_525) );
INVx1_ASAP7_75t_L g533 ( .A(n_315), .Y(n_533) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_315), .Y(n_685) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_315), .Y(n_710) );
AND2x2_ASAP7_75t_L g821 ( .A(n_315), .B(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g914 ( .A(n_315), .Y(n_914) );
BUFx2_ASAP7_75t_L g953 ( .A(n_315), .Y(n_953) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g838 ( .A(n_316), .Y(n_838) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx5_ASAP7_75t_SL g578 ( .A(n_320), .Y(n_578) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx3_ASAP7_75t_L g456 ( .A(n_323), .Y(n_456) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_323), .Y(n_460) );
INVx1_ASAP7_75t_L g529 ( .A(n_323), .Y(n_529) );
AND2x4_ASAP7_75t_L g331 ( .A(n_324), .B(n_332), .Y(n_331) );
AOI222xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_333), .B2(n_334), .C1(n_336), .C2(n_337), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g1060 ( .A1(n_328), .A2(n_583), .B1(n_760), .B2(n_1061), .C1(n_1062), .C2(n_1063), .Y(n_1060) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI222xp33_ASAP7_75t_L g1143 ( .A1(n_330), .A2(n_671), .B1(n_760), .B2(n_1144), .C1(n_1145), .C2(n_1146), .Y(n_1143) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g351 ( .A(n_331), .B(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_331), .Y(n_461) );
BUFx3_ASAP7_75t_L g522 ( .A(n_331), .Y(n_522) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_331), .Y(n_538) );
BUFx3_ASAP7_75t_L g978 ( .A(n_331), .Y(n_978) );
INVx1_ASAP7_75t_L g1013 ( .A(n_331), .Y(n_1013) );
AOI222xp33_ASAP7_75t_L g382 ( .A1(n_333), .A2(n_336), .B1(n_383), .B2(n_384), .C1(n_387), .C2(n_392), .Y(n_382) );
INVx2_ASAP7_75t_L g503 ( .A(n_334), .Y(n_503) );
INVx2_ASAP7_75t_L g672 ( .A(n_334), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_334), .A2(n_337), .B1(n_736), .B2(n_737), .Y(n_735) );
AOI222xp33_ASAP7_75t_L g756 ( .A1(n_334), .A2(n_538), .B1(n_757), .B2(n_758), .C1(n_759), .C2(n_760), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g976 ( .A1(n_334), .A2(n_337), .B1(n_948), .B2(n_949), .C1(n_972), .C2(n_977), .Y(n_976) );
INVx2_ASAP7_75t_L g1110 ( .A(n_334), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_334), .A2(n_337), .B1(n_1580), .B2(n_1581), .Y(n_1579) );
INVx1_ASAP7_75t_L g832 ( .A(n_335), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_337), .A2(n_568), .B1(n_569), .B2(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_337), .A2(n_658), .B1(n_660), .B2(n_671), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g888 ( .A1(n_337), .A2(n_583), .B1(n_778), .B2(n_889), .C1(n_890), .C2(n_891), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_337), .A2(n_671), .B1(n_993), .B2(n_994), .Y(n_1033) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
AND2x4_ASAP7_75t_L g760 ( .A(n_338), .B(n_341), .Y(n_760) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g505 ( .A(n_340), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_340), .B(n_506), .Y(n_1578) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g352 ( .A(n_342), .Y(n_352) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_343), .B(n_469), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_347), .B2(n_348), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_346), .A2(n_348), .B1(n_762), .B2(n_763), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_346), .A2(n_511), .B1(n_893), .B2(n_894), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_346), .A2(n_348), .B1(n_971), .B2(n_980), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_346), .A2(n_348), .B1(n_996), .B2(n_997), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_346), .A2(n_348), .B1(n_1054), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_346), .A2(n_1099), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_346), .A2(n_1117), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_347), .A2(n_369), .B1(n_375), .B2(n_376), .Y(n_368) );
INVx4_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx5_ASAP7_75t_L g1117 ( .A(n_349), .Y(n_1117) );
NAND4xp25_ASAP7_75t_L g752 ( .A(n_350), .B(n_753), .C(n_756), .D(n_761), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g884 ( .A(n_350), .B(n_885), .C(n_888), .D(n_892), .Y(n_884) );
NAND3xp33_ASAP7_75t_L g975 ( .A(n_350), .B(n_976), .C(n_979), .Y(n_975) );
NAND4xp25_ASAP7_75t_L g987 ( .A(n_350), .B(n_988), .C(n_991), .D(n_995), .Y(n_987) );
NAND4xp25_ASAP7_75t_SL g1056 ( .A(n_350), .B(n_1057), .C(n_1060), .D(n_1064), .Y(n_1056) );
NAND4xp25_ASAP7_75t_L g1139 ( .A(n_350), .B(n_1140), .C(n_1143), .D(n_1147), .Y(n_1139) );
CKINVDCx11_ASAP7_75t_R g350 ( .A(n_351), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_351), .B(n_501), .C(n_502), .Y(n_500) );
AOI211xp5_ASAP7_75t_L g1106 ( .A1(n_351), .A2(n_1107), .B(n_1108), .C(n_1109), .Y(n_1106) );
OAI31xp33_ASAP7_75t_L g572 ( .A1(n_353), .A2(n_573), .A3(n_579), .B(n_584), .Y(n_572) );
OAI31xp33_ASAP7_75t_L g666 ( .A1(n_353), .A2(n_667), .A3(n_668), .B(n_673), .Y(n_666) );
OAI31xp33_ASAP7_75t_SL g729 ( .A1(n_353), .A2(n_730), .A3(n_731), .B(n_738), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_353), .A2(n_404), .B1(n_752), .B2(n_764), .C(n_772), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_353), .A2(n_884), .B1(n_895), .B2(n_903), .C(n_905), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g974 ( .A1(n_353), .A2(n_975), .B(n_981), .Y(n_974) );
AOI221x1_ASAP7_75t_L g986 ( .A1(n_353), .A2(n_571), .B1(n_987), .B2(n_998), .C(n_1007), .Y(n_986) );
OAI31xp33_ASAP7_75t_L g1030 ( .A1(n_353), .A2(n_1031), .A3(n_1032), .B(n_1034), .Y(n_1030) );
AOI221x1_ASAP7_75t_L g1042 ( .A1(n_353), .A2(n_571), .B1(n_1043), .B2(n_1056), .C(n_1066), .Y(n_1042) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_353), .A2(n_404), .B1(n_1094), .B2(n_1105), .C(n_1118), .Y(n_1093) );
AOI221x1_ASAP7_75t_L g1138 ( .A1(n_353), .A2(n_404), .B1(n_1139), .B2(n_1150), .C(n_1158), .Y(n_1138) );
OAI31xp33_ASAP7_75t_SL g1573 ( .A1(n_353), .A2(n_1574), .A3(n_1575), .B(n_1582), .Y(n_1573) );
CKINVDCx16_ASAP7_75t_R g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g436 ( .A(n_355), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g704 ( .A(n_355), .B(n_437), .Y(n_704) );
AND2x4_ASAP7_75t_L g1475 ( .A(n_355), .B(n_1476), .Y(n_1475) );
NAND4xp25_ASAP7_75t_SL g356 ( .A(n_357), .B(n_368), .C(n_382), .D(n_394), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND4xp25_ASAP7_75t_L g806 ( .A(n_358), .B(n_807), .C(n_811), .D(n_814), .Y(n_806) );
NAND4xp25_ASAP7_75t_L g895 ( .A(n_358), .B(n_896), .C(n_899), .D(n_901), .Y(n_895) );
NAND4xp25_ASAP7_75t_L g998 ( .A(n_358), .B(n_999), .C(n_1002), .D(n_1005), .Y(n_998) );
INVx5_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_SL g478 ( .A(n_359), .B(n_479), .Y(n_478) );
CKINVDCx8_ASAP7_75t_R g566 ( .A(n_359), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g1044 ( .A(n_359), .B(n_1045), .Y(n_1044) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_359), .A2(n_369), .B1(n_376), .B2(n_1149), .C(n_1154), .Y(n_1153) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x6_ASAP7_75t_L g401 ( .A(n_361), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g496 ( .A(n_361), .Y(n_496) );
AND2x2_ASAP7_75t_L g946 ( .A(n_361), .B(n_718), .Y(n_946) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x6_ASAP7_75t_L g392 ( .A(n_362), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_363), .Y(n_371) );
INVx1_ASAP7_75t_L g378 ( .A(n_363), .Y(n_378) );
AND2x2_ASAP7_75t_L g414 ( .A(n_363), .B(n_406), .Y(n_414) );
INVx2_ASAP7_75t_L g438 ( .A(n_363), .Y(n_438) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_364), .Y(n_718) );
INVx2_ASAP7_75t_L g728 ( .A(n_364), .Y(n_728) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_364), .Y(n_792) );
INVx1_ASAP7_75t_L g1026 ( .A(n_364), .Y(n_1026) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_365), .Y(n_386) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx2_ASAP7_75t_L g373 ( .A(n_366), .Y(n_373) );
AND2x4_ASAP7_75t_L g402 ( .A(n_366), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g374 ( .A(n_367), .Y(n_374) );
AND2x4_ASAP7_75t_L g380 ( .A(n_367), .B(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_369), .A2(n_376), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx4_ASAP7_75t_L g561 ( .A(n_369), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_369), .A2(n_376), .B1(n_763), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_369), .A2(n_376), .B1(n_812), .B2(n_813), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_369), .A2(n_376), .B1(n_886), .B2(n_900), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_369), .A2(n_376), .B1(n_997), .B2(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_369), .A2(n_376), .B1(n_1054), .B2(n_1055), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_369), .A2(n_376), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
AND2x4_ASAP7_75t_L g388 ( .A(n_370), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_SL g659 ( .A(n_370), .B(n_389), .Y(n_659) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx6_ASAP7_75t_L g399 ( .A(n_372), .Y(n_399) );
INVx2_ASAP7_75t_L g433 ( .A(n_372), .Y(n_433) );
BUFx2_ASAP7_75t_L g631 ( .A(n_372), .Y(n_631) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_372), .B(n_1477), .Y(n_1476) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g393 ( .A(n_373), .Y(n_393) );
INVx1_ASAP7_75t_L g391 ( .A(n_374), .Y(n_391) );
INVx4_ASAP7_75t_L g562 ( .A(n_376), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_376), .A2(n_401), .B1(n_662), .B2(n_663), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_376), .A2(n_401), .B1(n_745), .B2(n_746), .Y(n_744) );
AND2x6_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
AND2x4_ASAP7_75t_L g397 ( .A(n_377), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g809 ( .A(n_377), .B(n_398), .Y(n_809) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g488 ( .A(n_378), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g628 ( .A(n_379), .Y(n_628) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_379), .Y(n_724) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_379), .Y(n_935) );
INVx1_ASAP7_75t_L g1169 ( .A(n_379), .Y(n_1169) );
INVx1_ASAP7_75t_L g1512 ( .A(n_379), .Y(n_1512) );
INVx2_ASAP7_75t_L g1541 ( .A(n_379), .Y(n_1541) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g422 ( .A(n_380), .Y(n_422) );
INVx1_ASAP7_75t_L g550 ( .A(n_380), .Y(n_550) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_380), .Y(n_696) );
INVx1_ASAP7_75t_L g721 ( .A(n_380), .Y(n_721) );
INVx1_ASAP7_75t_L g484 ( .A(n_381), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_384), .A2(n_387), .B1(n_392), .B2(n_889), .C1(n_891), .C2(n_902), .Y(n_901) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx4f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_386), .Y(n_428) );
INVx2_ASAP7_75t_SL g545 ( .A(n_386), .Y(n_545) );
INVx1_ASAP7_75t_L g657 ( .A(n_386), .Y(n_657) );
BUFx3_ASAP7_75t_L g797 ( .A(n_386), .Y(n_797) );
AND2x4_ASAP7_75t_L g1502 ( .A(n_386), .B(n_1484), .Y(n_1502) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_387), .A2(n_392), .B1(n_993), .B2(n_994), .C1(n_1003), .C2(n_1004), .Y(n_1002) );
BUFx4f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_388), .A2(n_392), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_388), .A2(n_392), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g1038 ( .A1(n_388), .A2(n_392), .B1(n_993), .B2(n_994), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1587 ( .A1(n_388), .A2(n_392), .B1(n_1580), .B2(n_1581), .Y(n_1587) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g489 ( .A(n_390), .Y(n_489) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g637 ( .A(n_391), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_392), .A2(n_487), .B1(n_488), .B2(n_490), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_392), .A2(n_655), .B1(n_656), .B2(n_658), .C1(n_659), .C2(n_660), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g741 ( .A1(n_392), .A2(n_488), .B1(n_736), .B2(n_737), .C1(n_742), .C2(n_743), .Y(n_741) );
AOI222xp33_ASAP7_75t_L g770 ( .A1(n_392), .A2(n_659), .B1(n_727), .B2(n_758), .C1(n_759), .C2(n_771), .Y(n_770) );
AOI222xp33_ASAP7_75t_L g814 ( .A1(n_392), .A2(n_659), .B1(n_797), .B2(n_815), .C1(n_816), .C2(n_817), .Y(n_814) );
INVx3_ASAP7_75t_L g1049 ( .A(n_392), .Y(n_1049) );
AOI222xp33_ASAP7_75t_L g1101 ( .A1(n_392), .A2(n_659), .B1(n_791), .B2(n_1102), .C1(n_1103), .C2(n_1104), .Y(n_1101) );
AOI222xp33_ASAP7_75t_L g1151 ( .A1(n_392), .A2(n_659), .B1(n_791), .B2(n_1145), .C1(n_1146), .C2(n_1152), .Y(n_1151) );
BUFx3_ASAP7_75t_L g639 ( .A(n_393), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_400), .B2(n_401), .Y(n_394) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_397), .A2(n_401), .B1(n_766), .B2(n_767), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_397), .A2(n_401), .B1(n_897), .B2(n_898), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_397), .A2(n_401), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g426 ( .A(n_399), .Y(n_426) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_399), .Y(n_548) );
INVx1_ASAP7_75t_L g726 ( .A(n_399), .Y(n_726) );
INVx2_ASAP7_75t_SL g790 ( .A(n_399), .Y(n_790) );
INVx2_ASAP7_75t_L g923 ( .A(n_399), .Y(n_923) );
CKINVDCx6p67_ASAP7_75t_R g498 ( .A(n_401), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_401), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
AOI22xp5_ASAP7_75t_SL g999 ( .A1(n_401), .A2(n_809), .B1(n_1000), .B2(n_1001), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_401), .A2(n_809), .B1(n_1051), .B2(n_1052), .Y(n_1050) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_401), .A2(n_809), .B1(n_1156), .B2(n_1157), .Y(n_1155) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_402), .Y(n_418) );
BUFx2_ASAP7_75t_L g554 ( .A(n_402), .Y(n_554) );
BUFx2_ASAP7_75t_L g626 ( .A(n_402), .Y(n_626) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_402), .Y(n_694) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_402), .Y(n_867) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_402), .Y(n_927) );
BUFx3_ASAP7_75t_L g934 ( .A(n_402), .Y(n_934) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_402), .Y(n_1075) );
INVx2_ASAP7_75t_SL g1505 ( .A(n_402), .Y(n_1505) );
INVx1_ASAP7_75t_L g485 ( .A(n_403), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_404), .A2(n_477), .B(n_494), .Y(n_476) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_404), .Y(n_571) );
INVx1_ASAP7_75t_L g904 ( .A(n_404), .Y(n_904) );
OAI31xp33_ASAP7_75t_SL g1583 ( .A1(n_404), .A2(n_1584), .A3(n_1585), .B(n_1586), .Y(n_1583) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
AND2x4_ASAP7_75t_L g665 ( .A(n_405), .B(n_407), .Y(n_665) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g437 ( .A(n_406), .B(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g415 ( .A(n_408), .Y(n_415) );
OR2x6_ASAP7_75t_L g614 ( .A(n_408), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_439), .Y(n_409) );
AOI33xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_416), .A3(n_423), .B1(n_429), .B2(n_430), .B3(n_434), .Y(n_410) );
AOI33xp33_ASAP7_75t_L g540 ( .A1(n_411), .A2(n_541), .A3(n_546), .B1(n_551), .B2(n_553), .B3(n_555), .Y(n_540) );
INVx1_ASAP7_75t_L g868 ( .A(n_411), .Y(n_868) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_412), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_412), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_412), .A2(n_435), .B1(n_1533), .B2(n_1542), .Y(n_1532) );
OR2x6_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
OR2x2_ASAP7_75t_L g966 ( .A(n_413), .B(n_415), .Y(n_966) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g699 ( .A(n_414), .Y(n_699) );
INVx1_ASAP7_75t_L g1508 ( .A(n_414), .Y(n_1508) );
AND2x4_ASAP7_75t_L g442 ( .A(n_415), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g514 ( .A(n_415), .B(n_443), .Y(n_514) );
OR2x2_ASAP7_75t_L g698 ( .A(n_415), .B(n_699), .Y(n_698) );
BUFx2_ASAP7_75t_L g861 ( .A(n_415), .Y(n_861) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_415), .B(n_848), .Y(n_1018) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g543 ( .A(n_418), .Y(n_543) );
INVx1_ASAP7_75t_L g1549 ( .A(n_418), .Y(n_1549) );
INVx2_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g1071 ( .A(n_420), .Y(n_1071) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g1520 ( .A(n_422), .B(n_1485), .Y(n_1520) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g938 ( .A(n_428), .Y(n_938) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g702 ( .A(n_433), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g930 ( .A(n_434), .B(n_931), .C(n_936), .Y(n_930) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g965 ( .A1(n_435), .A2(n_966), .B1(n_967), .B2(n_970), .Y(n_965) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_436), .Y(n_555) );
BUFx4f_ASAP7_75t_L g801 ( .A(n_436), .Y(n_801) );
INVx2_ASAP7_75t_L g1498 ( .A(n_437), .Y(n_1498) );
AND2x4_ASAP7_75t_L g1477 ( .A(n_438), .B(n_1478), .Y(n_1477) );
AOI33xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_444), .A3(n_450), .B1(n_457), .B2(n_458), .B3(n_462), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_440), .B(n_907), .C(n_910), .Y(n_906) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_442), .B(n_676), .C(n_681), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_442), .B(n_709), .C(n_711), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g773 ( .A(n_442), .B(n_774), .C(n_777), .Y(n_773) );
BUFx3_ASAP7_75t_L g958 ( .A(n_442), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_442), .B(n_1010), .C(n_1011), .Y(n_1009) );
AOI33xp33_ASAP7_75t_L g1076 ( .A1(n_442), .A2(n_464), .A3(n_1077), .B1(n_1080), .B2(n_1082), .B3(n_1083), .Y(n_1076) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_442), .B(n_1124), .C(n_1126), .Y(n_1123) );
NAND3xp33_ASAP7_75t_L g1159 ( .A(n_442), .B(n_1160), .C(n_1161), .Y(n_1159) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g612 ( .A(n_448), .Y(n_612) );
BUFx2_ASAP7_75t_L g687 ( .A(n_448), .Y(n_687) );
AND2x4_ASAP7_75t_L g855 ( .A(n_448), .B(n_822), .Y(n_855) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g519 ( .A(n_449), .Y(n_519) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_453), .B(n_1431), .Y(n_1438) );
CKINVDCx5p33_ASAP7_75t_R g1467 ( .A(n_454), .Y(n_1467) );
BUFx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g909 ( .A(n_455), .Y(n_909) );
AND2x4_ASAP7_75t_L g1430 ( .A(n_455), .B(n_1431), .Y(n_1430) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_456), .Y(n_536) );
INVx3_ASAP7_75t_L g680 ( .A(n_456), .Y(n_680) );
BUFx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_SL g916 ( .A(n_460), .Y(n_916) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_461), .Y(n_778) );
INVx2_ASAP7_75t_SL g919 ( .A(n_461), .Y(n_919) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI33xp33_ASAP7_75t_L g1450 ( .A1(n_463), .A2(n_614), .A3(n_1451), .B1(n_1454), .B2(n_1460), .B3(n_1466), .Y(n_1450) );
OAI33xp33_ASAP7_75t_L g1550 ( .A1(n_463), .A2(n_1551), .A3(n_1553), .B1(n_1560), .B2(n_1564), .B3(n_1569), .Y(n_1550) );
CKINVDCx8_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_464), .B(n_684), .C(n_686), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_464), .B(n_780), .C(n_783), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g912 ( .A(n_464), .B(n_913), .C(n_917), .Y(n_912) );
NAND3xp33_ASAP7_75t_L g1119 ( .A(n_464), .B(n_1120), .C(n_1121), .Y(n_1119) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx6_ASAP7_75t_L g539 ( .A(n_465), .Y(n_539) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g1431 ( .A(n_467), .B(n_822), .Y(n_1431) );
INVx2_ASAP7_75t_L g848 ( .A(n_468), .Y(n_848) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_556), .B1(n_644), .B2(n_645), .Y(n_472) );
INVx1_ASAP7_75t_L g645 ( .A(n_473), .Y(n_645) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_476), .B(n_499), .C(n_513), .D(n_540), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_491), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g1533 ( .A1(n_480), .A2(n_1534), .B1(n_1535), .B2(n_1536), .C(n_1537), .Y(n_1533) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g565 ( .A(n_483), .Y(n_565) );
INVx2_ASAP7_75t_L g623 ( .A(n_483), .Y(n_623) );
BUFx2_ASAP7_75t_L g874 ( .A(n_483), .Y(n_874) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
OR2x2_ASAP7_75t_L g497 ( .A(n_484), .B(n_485), .Y(n_497) );
INVx2_ASAP7_75t_L g1046 ( .A(n_488), .Y(n_1046) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g619 ( .A(n_497), .Y(n_619) );
INVx1_ASAP7_75t_L g641 ( .A(n_497), .Y(n_641) );
INVx1_ASAP7_75t_L g1496 ( .A(n_497), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1518 ( .A(n_497), .B(n_1485), .Y(n_1518) );
BUFx2_ASAP7_75t_L g1535 ( .A(n_497), .Y(n_1535) );
AO21x1_ASAP7_75t_SL g499 ( .A1(n_500), .A2(n_508), .B(n_512), .Y(n_499) );
INVx1_ASAP7_75t_L g583 ( .A(n_503), .Y(n_583) );
INVx1_ASAP7_75t_L g581 ( .A(n_504), .Y(n_581) );
OAI21xp5_ASAP7_75t_SL g845 ( .A1(n_504), .A2(n_815), .B(n_846), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_504), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_954) );
OAI22xp33_ASAP7_75t_SL g960 ( .A1(n_504), .A2(n_961), .B1(n_962), .B2(n_964), .Y(n_960) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g600 ( .A(n_505), .Y(n_600) );
INVx2_ASAP7_75t_L g734 ( .A(n_505), .Y(n_734) );
AOI33xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .A3(n_523), .B1(n_530), .B2(n_534), .B3(n_539), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_518), .Y(n_1084) );
INVx1_ASAP7_75t_L g1128 ( .A(n_518), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1436 ( .A(n_518), .B(n_1431), .Y(n_1436) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g531 ( .A(n_519), .Y(n_531) );
INVx2_ASAP7_75t_SL g785 ( .A(n_519), .Y(n_785) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g1085 ( .A(n_521), .Y(n_1085) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
AND2x4_ASAP7_75t_L g853 ( .A(n_522), .B(n_825), .Y(n_853) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g782 ( .A(n_528), .Y(n_782) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g827 ( .A(n_529), .Y(n_827) );
BUFx3_ASAP7_75t_L g911 ( .A(n_531), .Y(n_911) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g677 ( .A(n_533), .Y(n_677) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g594 ( .A(n_536), .Y(n_594) );
INVx2_ASAP7_75t_L g608 ( .A(n_536), .Y(n_608) );
INVx2_ASAP7_75t_L g714 ( .A(n_536), .Y(n_714) );
INVx3_ASAP7_75t_L g1016 ( .A(n_536), .Y(n_1016) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g689 ( .A(n_538), .Y(n_689) );
HB1xp67_ASAP7_75t_L g1081 ( .A(n_538), .Y(n_1081) );
INVx2_ASAP7_75t_L g601 ( .A(n_539), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_539), .B(n_713), .C(n_715), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g951 ( .A1(n_539), .A2(n_952), .B1(n_958), .B2(n_959), .C(n_965), .Y(n_951) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g692 ( .A(n_545), .Y(n_692) );
INVx1_ASAP7_75t_L g1069 ( .A(n_545), .Y(n_1069) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g552 ( .A(n_548), .Y(n_552) );
INVx1_ASAP7_75t_L g1024 ( .A(n_548), .Y(n_1024) );
INVx2_ASAP7_75t_L g1131 ( .A(n_548), .Y(n_1131) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g928 ( .A(n_550), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_555), .Y(n_616) );
AOI33xp33_ASAP7_75t_L g1067 ( .A1(n_555), .A2(n_697), .A3(n_1068), .B1(n_1070), .B2(n_1072), .B3(n_1074), .Y(n_1067) );
INVx1_ASAP7_75t_L g644 ( .A(n_556), .Y(n_644) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g642 ( .A(n_558), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_572), .C(n_585), .Y(n_558) );
OAI31xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .A3(n_570), .B(n_571), .Y(n_559) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g1048 ( .A(n_565), .Y(n_1048) );
NAND3xp33_ASAP7_75t_SL g653 ( .A(n_566), .B(n_654), .C(n_661), .Y(n_653) );
NAND3xp33_ASAP7_75t_SL g740 ( .A(n_566), .B(n_741), .C(n_744), .Y(n_740) );
NAND4xp25_ASAP7_75t_SL g764 ( .A(n_566), .B(n_765), .C(n_768), .D(n_770), .Y(n_764) );
NAND4xp25_ASAP7_75t_L g1094 ( .A(n_566), .B(n_1095), .C(n_1098), .D(n_1101), .Y(n_1094) );
AOI221x1_ASAP7_75t_L g805 ( .A1(n_571), .A2(n_806), .B1(n_818), .B2(n_859), .C(n_862), .Y(n_805) );
OAI31xp33_ASAP7_75t_L g1035 ( .A1(n_571), .A2(n_1036), .A3(n_1037), .B(n_1039), .Y(n_1035) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g605 ( .A(n_576), .Y(n_605) );
BUFx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g591 ( .A(n_577), .Y(n_591) );
INVx1_ASAP7_75t_L g1464 ( .A(n_577), .Y(n_1464) );
OAI22xp33_ASAP7_75t_L g1451 ( .A1(n_580), .A2(n_962), .B1(n_1452), .B2(n_1453), .Y(n_1451) );
OAI22xp33_ASAP7_75t_L g1466 ( .A1(n_580), .A2(n_1467), .B1(n_1468), .B2(n_1469), .Y(n_1466) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g1563 ( .A(n_581), .Y(n_1563) );
AOI222xp33_ASAP7_75t_L g991 ( .A1(n_583), .A2(n_613), .B1(n_760), .B2(n_992), .C1(n_993), .C2(n_994), .Y(n_991) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_602), .C(n_629), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_595), .C(n_601), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_592), .B2(n_593), .Y(n_587) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
HB1xp67_ASAP7_75t_L g1567 ( .A(n_591), .Y(n_1567) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI22xp33_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_597), .B1(n_598), .B2(n_599), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g1460 ( .A1(n_597), .A2(n_1461), .B1(n_1462), .B2(n_1465), .Y(n_1460) );
OAI22xp33_ASAP7_75t_L g1569 ( .A1(n_599), .A2(n_1570), .B1(n_1571), .B2(n_1572), .Y(n_1569) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g669 ( .A(n_600), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_614), .B1(n_616), .B2(n_617), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_607), .B2(n_609), .C(n_610), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g1454 ( .A1(n_604), .A2(n_1455), .B1(n_1456), .B2(n_1459), .Y(n_1454) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_SL g682 ( .A(n_612), .Y(n_682) );
INVx2_ASAP7_75t_L g1122 ( .A(n_612), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_613), .Y(n_1107) );
INVx1_ASAP7_75t_L g1552 ( .A(n_614), .Y(n_1552) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_616), .A2(n_863), .B1(n_868), .B2(n_869), .Y(n_862) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B1(n_621), .B2(n_624), .C(n_625), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_618), .A2(n_955), .B1(n_957), .B2(n_968), .C(n_969), .Y(n_967) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_618), .A2(n_968), .B1(n_971), .B2(n_972), .C(n_973), .Y(n_970) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_619), .Y(n_871) );
OAI21xp33_ASAP7_75t_SL g632 ( .A1(n_621), .A2(n_633), .B(n_634), .Y(n_632) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI221xp5_ASAP7_75t_SL g863 ( .A1(n_623), .A2(n_640), .B1(n_842), .B2(n_864), .C(n_865), .Y(n_863) );
BUFx3_ASAP7_75t_L g968 ( .A(n_623), .Y(n_968) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g876 ( .A(n_628), .Y(n_876) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g1489 ( .A(n_637), .Y(n_1489) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_639), .B(n_1477), .Y(n_1491) );
BUFx2_ASAP7_75t_L g1543 ( .A(n_640), .Y(n_1543) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
XOR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_879), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_749), .B1(n_877), .B2(n_878), .Y(n_648) );
INVx2_ASAP7_75t_L g877 ( .A(n_649), .Y(n_877) );
XOR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_705), .Y(n_649) );
NAND3x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_666), .C(n_674), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_664), .B(n_665), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g743 ( .A(n_657), .Y(n_743) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_665), .A2(n_740), .B(n_747), .Y(n_739) );
OAI31xp33_ASAP7_75t_L g942 ( .A1(n_665), .A2(n_943), .A3(n_944), .B(n_950), .Y(n_942) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND4x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_683), .C(n_690), .D(n_700), .Y(n_674) );
INVx1_ASAP7_75t_L g1570 ( .A(n_678), .Y(n_1570) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g776 ( .A(n_680), .Y(n_776) );
INVx1_ASAP7_75t_L g1458 ( .A(n_680), .Y(n_1458) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .C(n_697), .Y(n_690) );
BUFx3_ASAP7_75t_L g799 ( .A(n_694), .Y(n_799) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx3_ASAP7_75t_L g800 ( .A(n_696), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_697), .B(n_717), .C(n_719), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g1019 ( .A(n_697), .B(n_1020), .C(n_1021), .Y(n_1019) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_697), .B(n_1130), .C(n_1132), .Y(n_1129) );
NAND3xp33_ASAP7_75t_L g1165 ( .A(n_697), .B(n_1166), .C(n_1167), .Y(n_1165) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .C(n_704), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g722 ( .A(n_704), .B(n_723), .C(n_725), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_704), .B(n_1023), .C(n_1027), .Y(n_1022) );
NAND3xp33_ASAP7_75t_L g1133 ( .A(n_704), .B(n_1134), .C(n_1135), .Y(n_1133) );
NAND3xp33_ASAP7_75t_L g1170 ( .A(n_704), .B(n_1171), .C(n_1172), .Y(n_1170) );
XOR2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_748), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_729), .C(n_739), .Y(n_706) );
AND4x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .C(n_716), .D(n_722), .Y(n_707) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_718), .Y(n_1003) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g1545 ( .A(n_724), .Y(n_1545) );
HB1xp67_ASAP7_75t_L g1510 ( .A(n_726), .Y(n_1510) );
INVx1_ASAP7_75t_L g1507 ( .A(n_727), .Y(n_1507) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx3_ASAP7_75t_L g1073 ( .A(n_728), .Y(n_1073) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR2x6_ASAP7_75t_L g850 ( .A(n_734), .B(n_834), .Y(n_850) );
INVx1_ASAP7_75t_L g878 ( .A(n_749), .Y(n_878) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_804), .Y(n_749) );
INVx1_ASAP7_75t_L g803 ( .A(n_751), .Y(n_803) );
NAND4xp25_ASAP7_75t_SL g772 ( .A(n_773), .B(n_779), .C(n_786), .D(n_795), .Y(n_772) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
BUFx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_785), .B(n_858), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_793), .C(n_794), .Y(n_786) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AND2x4_ASAP7_75t_L g1513 ( .A(n_792), .B(n_1514), .Y(n_1513) );
NAND3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .C(n_801), .Y(n_795) );
AOI222xp33_ASAP7_75t_L g851 ( .A1(n_812), .A2(n_852), .B1(n_853), .B2(n_854), .C1(n_855), .C2(n_856), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_828), .C(n_851), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_821), .B1(n_823), .B2(n_824), .Y(n_819) );
INVx2_ASAP7_75t_L g826 ( .A(n_822), .Y(n_826) );
AND2x4_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1079 ( .A(n_827), .Y(n_1079) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_844), .C(n_849), .Y(n_828) );
NAND2x1p5_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .Y(n_830) );
NAND2x1_ASAP7_75t_SL g1442 ( .A(n_831), .B(n_1443), .Y(n_1442) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OR2x6_ASAP7_75t_L g837 ( .A(n_834), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g858 ( .A(n_834), .Y(n_858) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g1447 ( .A(n_838), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI221xp5_ASAP7_75t_SL g869 ( .A1(n_852), .A2(n_854), .B1(n_870), .B2(n_872), .C(n_875), .Y(n_869) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
AOI31xp33_ASAP7_75t_L g1481 ( .A1(n_859), .A2(n_1482), .A3(n_1499), .B(n_1516), .Y(n_1481) );
INVx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
CKINVDCx8_ASAP7_75t_R g860 ( .A(n_861), .Y(n_860) );
BUFx4f_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_SL g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g1494 ( .A(n_874), .Y(n_1494) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
XNOR2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_939), .Y(n_880) );
XNOR2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
NAND4xp25_ASAP7_75t_L g905 ( .A(n_906), .B(n_912), .C(n_920), .D(n_930), .Y(n_905) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVxp67_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_924), .C(n_929), .Y(n_920) );
BUFx3_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
AND2x4_ASAP7_75t_L g1483 ( .A(n_927), .B(n_1484), .Y(n_1483) );
INVx2_ASAP7_75t_SL g1539 ( .A(n_927), .Y(n_1539) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx2_ASAP7_75t_SL g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
XNOR2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
NAND3x1_ASAP7_75t_SL g941 ( .A(n_942), .B(n_951), .C(n_974), .Y(n_941) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx3_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
BUFx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AND2x6_ASAP7_75t_L g1433 ( .A(n_978), .B(n_1431), .Y(n_1433) );
NAND2x1p5_ASAP7_75t_L g1449 ( .A(n_978), .B(n_1443), .Y(n_1449) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_1089), .B1(n_1176), .B2(n_1177), .Y(n_982) );
INVx1_ASAP7_75t_L g1177 ( .A(n_983), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_1040), .B1(n_1087), .B2(n_1088), .Y(n_984) );
INVx1_ASAP7_75t_L g1087 ( .A(n_985), .Y(n_1087) );
INVx1_ASAP7_75t_L g1034 ( .A(n_988), .Y(n_1034) );
INVx1_ASAP7_75t_L g1031 ( .A(n_995), .Y(n_1031) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_999), .Y(n_1036) );
INVxp67_ASAP7_75t_L g1039 ( .A(n_1005), .Y(n_1039) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1029 ( .A(n_1008), .B(n_1030), .C(n_1035), .Y(n_1029) );
AND4x1_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1014), .C(n_1019), .D(n_1022), .Y(n_1008) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
NAND3xp33_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1017), .C(n_1018), .Y(n_1014) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_1018), .B(n_1163), .C(n_1164), .Y(n_1162) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1040), .Y(n_1088) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
NAND3xp33_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1050), .C(n_1053), .Y(n_1043) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1076), .Y(n_1066) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1079), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1265 ( .A1(n_1086), .A2(n_1266), .B1(n_1267), .B2(n_1268), .Y(n_1265) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1089), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1136), .B1(n_1137), .B2(n_1175), .Y(n_1091) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1092), .Y(n_1175) );
NAND3xp33_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1112), .C(n_1115), .Y(n_1105) );
NAND4xp25_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1123), .C(n_1129), .D(n_1133), .Y(n_1118) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1138), .Y(n_1174) );
NAND3xp33_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1153), .C(n_1155), .Y(n_1150) );
NAND4xp25_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1162), .C(n_1165), .D(n_1170), .Y(n_1158) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
OAI21xp33_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1187), .B(n_1420), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
OAI22xp5_ASAP7_75t_SL g1224 ( .A1(n_1181), .A2(n_1225), .B1(n_1226), .B2(n_1227), .Y(n_1224) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1181), .Y(n_1238) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1185), .Y(n_1182) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1183), .Y(n_1208) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1184), .B(n_1200), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1185), .B(n_1208), .Y(n_1207) );
AND2x4_ASAP7_75t_L g1218 ( .A(n_1185), .B(n_1208), .Y(n_1218) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1186), .Y(n_1200) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1352), .Y(n_1187) );
OAI211xp5_ASAP7_75t_L g1188 ( .A1(n_1189), .A2(n_1296), .B(n_1323), .C(n_1339), .Y(n_1188) );
AOI21xp33_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1271), .B(n_1272), .Y(n_1189) );
AOI21xp5_ASAP7_75t_L g1296 ( .A1(n_1190), .A2(n_1297), .B(n_1322), .Y(n_1296) );
OAI211xp5_ASAP7_75t_L g1190 ( .A1(n_1191), .A2(n_1212), .B(n_1228), .C(n_1253), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1381 ( .A(n_1191), .B(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1209), .Y(n_1192) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1193), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1193), .B(n_1209), .Y(n_1315) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1194), .B(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1194), .B(n_1232), .Y(n_1258) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1195), .B(n_1250), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1195), .B(n_1232), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1206), .Y(n_1195) );
AND2x4_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1201), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1199), .B(n_1202), .Y(n_1242) );
HB1xp67_ASAP7_75t_L g1594 ( .A(n_1200), .Y(n_1594) );
AND2x4_ASAP7_75t_L g1203 ( .A(n_1201), .B(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1202), .B(n_1205), .Y(n_1245) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1592 ( .A(n_1208), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1209), .B(n_1236), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1209), .B(n_1249), .Y(n_1248) );
CKINVDCx5p33_ASAP7_75t_R g1260 ( .A(n_1209), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1209), .B(n_1279), .Y(n_1278) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1209), .B(n_1279), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1209), .B(n_1232), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1209), .B(n_1258), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1333 ( .A(n_1209), .B(n_1313), .Y(n_1333) );
NOR2xp33_ASAP7_75t_L g1342 ( .A(n_1209), .B(n_1312), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1209), .B(n_1230), .Y(n_1387) );
AND2x4_ASAP7_75t_SL g1209 ( .A(n_1210), .B(n_1211), .Y(n_1209) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1212), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1212), .B(n_1351), .Y(n_1350) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1222), .Y(n_1212) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1213), .Y(n_1356) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1213), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1219), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1214), .B(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1215), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1215), .B(n_1256), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1215), .B(n_1219), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1215), .B(n_1222), .Y(n_1321) );
BUFx6f_ASAP7_75t_L g1329 ( .A(n_1215), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1217), .Y(n_1215) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1218), .Y(n_1225) );
BUFx3_ASAP7_75t_L g1264 ( .A(n_1218), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1219), .B(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1219), .Y(n_1256) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1219), .Y(n_1295) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1219), .Y(n_1319) );
AOI321xp33_ASAP7_75t_L g1339 ( .A1(n_1219), .A2(n_1340), .A3(n_1343), .B1(n_1345), .B2(n_1347), .C(n_1350), .Y(n_1339) );
NAND2xp5_ASAP7_75t_SL g1345 ( .A(n_1219), .B(n_1346), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1221), .Y(n_1219) );
CKINVDCx6p67_ASAP7_75t_R g1247 ( .A(n_1222), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1222), .B(n_1262), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1222), .B(n_1252), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1222), .B(n_1318), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g1322 ( .A(n_1222), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1397 ( .A(n_1222), .B(n_1252), .Y(n_1397) );
OR2x6_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1402 ( .A(n_1223), .B(n_1224), .Y(n_1402) );
AOI22xp5_ASAP7_75t_L g1228 ( .A1(n_1229), .A2(n_1246), .B1(n_1248), .B2(n_1251), .Y(n_1228) );
O2A1O1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1229), .A2(n_1281), .B(n_1285), .C(n_1286), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1235), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1230), .B(n_1358), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1230), .B(n_1260), .Y(n_1378) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVxp67_ASAP7_75t_SL g1250 ( .A(n_1232), .Y(n_1250) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1232), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1234), .Y(n_1232) );
AOI211xp5_ASAP7_75t_L g1300 ( .A1(n_1235), .A2(n_1287), .B(n_1301), .C(n_1305), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1235), .B(n_1249), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1235), .B(n_1258), .Y(n_1385) );
INVx2_ASAP7_75t_SL g1277 ( .A(n_1236), .Y(n_1277) );
BUFx2_ASAP7_75t_L g1283 ( .A(n_1236), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1303 ( .A(n_1236), .B(n_1256), .Y(n_1303) );
BUFx3_ASAP7_75t_L g1310 ( .A(n_1236), .Y(n_1310) );
INVx2_ASAP7_75t_SL g1236 ( .A(n_1237), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1237), .B(n_1260), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1237), .B(n_1256), .Y(n_1401) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_1240), .A2(n_1241), .B1(n_1243), .B2(n_1244), .Y(n_1239) );
BUFx3_ASAP7_75t_L g1267 ( .A(n_1241), .Y(n_1267) );
BUFx6f_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
HB1xp67_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1245), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_1246), .A2(n_1291), .B1(n_1394), .B2(n_1396), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1247), .B(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1247), .B(n_1261), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1247), .B(n_1274), .Y(n_1405) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1248), .Y(n_1351) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1249), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1249), .B(n_1260), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1249), .B(n_1259), .Y(n_1417) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1251), .Y(n_1346) );
AOI21xp33_ASAP7_75t_SL g1398 ( .A1(n_1251), .A2(n_1294), .B(n_1399), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1252), .B(n_1261), .Y(n_1344) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1252), .Y(n_1412) );
A2O1A1Ixp33_ASAP7_75t_SL g1253 ( .A1(n_1254), .A2(n_1257), .B(n_1261), .C(n_1270), .Y(n_1253) );
NOR2xp33_ASAP7_75t_L g1418 ( .A(n_1254), .B(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1255), .B(n_1277), .Y(n_1361) );
OAI21xp33_ASAP7_75t_L g1386 ( .A1(n_1255), .A2(n_1324), .B(n_1387), .Y(n_1386) );
OAI21xp5_ASAP7_75t_L g1390 ( .A1(n_1255), .A2(n_1375), .B(n_1391), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1259), .Y(n_1257) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1258), .Y(n_1287) );
OAI21xp5_ASAP7_75t_SL g1334 ( .A1(n_1258), .A2(n_1335), .B(n_1336), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1258), .B(n_1277), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1260), .B(n_1282), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1260), .B(n_1325), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1260), .B(n_1349), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1260), .B(n_1304), .Y(n_1364) );
INVx2_ASAP7_75t_L g1338 ( .A(n_1261), .Y(n_1338) );
A2O1A1Ixp33_ASAP7_75t_L g1362 ( .A1(n_1261), .A2(n_1328), .B(n_1363), .C(n_1365), .Y(n_1362) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1270), .Y(n_1406) );
OAI211xp5_ASAP7_75t_SL g1272 ( .A1(n_1273), .A2(n_1275), .B(n_1280), .C(n_1290), .Y(n_1272) );
A2O1A1Ixp33_ASAP7_75t_L g1354 ( .A1(n_1273), .A2(n_1275), .B(n_1292), .C(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1274), .B(n_1283), .Y(n_1289) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
NOR2xp33_ASAP7_75t_L g1305 ( .A(n_1277), .B(n_1284), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1277), .B(n_1315), .Y(n_1314) );
NOR2x1p5_ASAP7_75t_L g1325 ( .A(n_1277), .B(n_1287), .Y(n_1325) );
HB1xp67_ASAP7_75t_L g1377 ( .A(n_1277), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1278), .B(n_1310), .Y(n_1392) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1283), .B(n_1293), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1332 ( .A(n_1283), .B(n_1333), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1283), .B(n_1342), .Y(n_1341) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1283), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1283), .B(n_1412), .Y(n_1411) );
NOR2xp33_ASAP7_75t_L g1359 ( .A(n_1284), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1285), .Y(n_1309) );
AOI21xp33_ASAP7_75t_SL g1286 ( .A1(n_1287), .A2(n_1288), .B(n_1289), .Y(n_1286) );
OAI21xp33_ASAP7_75t_L g1394 ( .A1(n_1288), .A2(n_1367), .B(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1289), .Y(n_1336) );
OAI21xp5_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1294), .B(n_1295), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1293), .Y(n_1409) );
NAND2xp67_ASAP7_75t_L g1371 ( .A(n_1295), .B(n_1372), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1295), .B(n_1417), .Y(n_1416) );
OAI211xp5_ASAP7_75t_L g1297 ( .A1(n_1298), .A2(n_1300), .B(n_1306), .C(n_1307), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1304), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1303), .B(n_1378), .Y(n_1380) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1304), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1404 ( .A(n_1304), .B(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1306), .Y(n_1327) );
A2O1A1Ixp33_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1311), .B(n_1314), .C(n_1316), .Y(n_1307) );
NOR2xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1310), .Y(n_1308) );
O2A1O1Ixp33_ASAP7_75t_SL g1330 ( .A1(n_1309), .A2(n_1331), .B(n_1334), .C(n_1337), .Y(n_1330) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1310), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1310), .B(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1320), .Y(n_1316) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1318), .Y(n_1369) );
INVx3_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
AOI31xp33_ASAP7_75t_L g1373 ( .A1(n_1322), .A2(n_1374), .A3(n_1384), .B(n_1386), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1326), .B1(n_1327), .B2(n_1328), .C(n_1330), .Y(n_1323) );
AOI211xp5_ASAP7_75t_L g1374 ( .A1(n_1328), .A2(n_1375), .B(n_1379), .C(n_1381), .Y(n_1374) );
CKINVDCx14_ASAP7_75t_R g1328 ( .A(n_1329), .Y(n_1328) );
OAI21xp33_ASAP7_75t_L g1384 ( .A1(n_1329), .A2(n_1370), .B(n_1385), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g1407 ( .A1(n_1329), .A2(n_1363), .B1(n_1408), .B2(n_1410), .C(n_1413), .Y(n_1407) );
INVxp67_ASAP7_75t_SL g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1335), .Y(n_1395) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_1337), .A2(n_1356), .B(n_1357), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1388 ( .A1(n_1337), .A2(n_1389), .B1(n_1406), .B2(n_1407), .Y(n_1388) );
INVx3_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1342), .B(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1388), .Y(n_1352) );
O2A1O1Ixp33_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1359), .B(n_1362), .C(n_1373), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1358), .B(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1364), .Y(n_1419) );
AOI21xp5_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1368), .B(n_1370), .Y(n_1365) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1369), .Y(n_1414) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1378), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1408 ( .A(n_1378), .B(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
AOI211xp5_ASAP7_75t_SL g1413 ( .A1(n_1385), .A2(n_1414), .B(n_1415), .C(n_1418), .Y(n_1413) );
NAND4xp25_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1393), .C(n_1398), .D(n_1404), .Y(n_1389) );
INVxp67_ASAP7_75t_SL g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
NOR3xp33_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1402), .C(n_1403), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1424), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1470), .Y(n_1424) );
NOR3xp33_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1439), .C(n_1450), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1434), .Y(n_1426) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_1428), .A2(n_1429), .B1(n_1432), .B2(n_1433), .Y(n_1427) );
BUFx2_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
OAI221xp5_ASAP7_75t_L g1493 ( .A1(n_1432), .A2(n_1435), .B1(n_1494), .B2(n_1495), .C(n_1497), .Y(n_1493) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_1435), .A2(n_1436), .B1(n_1437), .B2(n_1438), .Y(n_1434) );
INVx2_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx2_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
NAND2x1p5_ASAP7_75t_L g1446 ( .A(n_1443), .B(n_1447), .Y(n_1446) );
INVx3_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
BUFx4f_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
BUFx2_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx2_ASAP7_75t_SL g1456 ( .A(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1458), .Y(n_1558) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_1461), .A2(n_1468), .B1(n_1517), .B2(n_1519), .Y(n_1516) );
BUFx2_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
BUFx3_ASAP7_75t_L g1556 ( .A(n_1464), .Y(n_1556) );
AOI211xp5_ASAP7_75t_L g1482 ( .A1(n_1465), .A2(n_1483), .B(n_1486), .C(n_1492), .Y(n_1482) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_1469), .A2(n_1500), .B1(n_1503), .B2(n_1509), .C(n_1513), .Y(n_1499) );
AOI21xp5_ASAP7_75t_L g1470 ( .A1(n_1471), .A2(n_1480), .B(n_1481), .Y(n_1470) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
AND2x4_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1474), .Y(n_1472) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
AND2x4_ASAP7_75t_L g1488 ( .A(n_1477), .B(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1477), .Y(n_1515) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx2_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx2_ASAP7_75t_SL g1490 ( .A(n_1491), .Y(n_1490) );
INVx2_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
INVx2_ASAP7_75t_SL g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_SL g1514 ( .A(n_1515), .Y(n_1514) );
INVx6_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
INVx4_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
BUFx2_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVxp67_ASAP7_75t_SL g1525 ( .A(n_1526), .Y(n_1525) );
HB1xp67_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
HB1xp67_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
NAND3xp33_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1573), .C(n_1583), .Y(n_1530) );
NOR2xp33_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1550), .Y(n_1531) );
OAI22xp33_ASAP7_75t_L g1560 ( .A1(n_1534), .A2(n_1536), .B1(n_1561), .B2(n_1563), .Y(n_1560) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
OAI221xp5_ASAP7_75t_L g1542 ( .A1(n_1543), .A2(n_1544), .B1(n_1545), .B2(n_1546), .C(n_1547), .Y(n_1542) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
OAI22xp5_ASAP7_75t_L g1553 ( .A1(n_1554), .A2(n_1555), .B1(n_1557), .B2(n_1559), .Y(n_1553) );
INVx2_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
OAI22xp33_ASAP7_75t_L g1564 ( .A1(n_1561), .A2(n_1565), .B1(n_1566), .B2(n_1568), .Y(n_1564) );
INVx2_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
BUFx3_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
BUFx6f_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
A2O1A1Ixp33_ASAP7_75t_L g1590 ( .A1(n_1589), .A2(n_1591), .B(n_1593), .C(n_1595), .Y(n_1590) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
endmodule