module fake_netlist_5_127_n_1230 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1230);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1230;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_171;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1121;
wire n_314;
wire n_604;
wire n_368;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_1010;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_829;
wire n_361;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_174;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_210;
wire n_774;
wire n_1059;
wire n_176;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_177;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_181;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1026;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_101),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_65),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_109),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_13),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_57),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_122),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_123),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_69),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_77),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_99),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_112),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_102),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_52),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_155),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_38),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_45),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_104),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_6),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_76),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_27),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_45),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_61),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_74),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_57),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_170),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_58),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_35),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_61),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_25),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_16),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_18),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_47),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_145),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_56),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_82),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_48),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_160),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_163),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_110),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_23),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_124),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_148),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_41),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_35),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_91),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_129),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_157),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_85),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_97),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_159),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_167),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_111),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_13),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_162),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_84),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_21),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_150),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_87),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_152),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_63),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_92),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_64),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_42),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_48),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_73),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_169),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_16),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_139),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_25),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_29),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_134),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_153),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_158),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_46),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_140),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_12),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_165),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_34),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_67),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_55),
.Y(n_285)
);

BUFx8_ASAP7_75t_SL g286 ( 
.A(n_19),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_7),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_103),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_18),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_51),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_219),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_181),
.B(n_0),
.Y(n_293)
);

INVxp33_ASAP7_75t_SL g294 ( 
.A(n_182),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_200),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_182),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_272),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_183),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_286),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_203),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_183),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_189),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_0),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_191),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_209),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_206),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_192),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_228),
.B(n_1),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_265),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_174),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_207),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_193),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_210),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_231),
.B(n_1),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_265),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_174),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_252),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_231),
.B(n_2),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_218),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_220),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_229),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_234),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_287),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_196),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_198),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_202),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_243),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_287),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_204),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_287),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_184),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_194),
.B(n_2),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_241),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_246),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_287),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_205),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_174),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_211),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_247),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_187),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_256),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_267),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_212),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_213),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_187),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_173),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_217),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_197),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_268),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_221),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_271),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_273),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_222),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_276),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_175),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_291),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_225),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_276),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_184),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_227),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_194),
.B(n_3),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_230),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_274),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_274),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_254),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_254),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_180),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_377),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_176),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_296),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_353),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_171),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_305),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_171),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_337),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_305),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

CKINVDCx8_ASAP7_75t_R g403 ( 
.A(n_292),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_315),
.B(n_180),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_302),
.B(n_201),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_303),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_304),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_306),
.B(n_307),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_313),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_319),
.B(n_201),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_172),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g417 ( 
.A(n_318),
.B(n_224),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_325),
.B(n_326),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_333),
.A2(n_244),
.B(n_224),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_334),
.B(n_172),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_340),
.B(n_177),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_301),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_301),
.B(n_244),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_313),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_345),
.B(n_371),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_375),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_314),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_323),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_310),
.Y(n_440)
);

BUFx8_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_324),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_329),
.B(n_276),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_293),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_316),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_295),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_311),
.B(n_177),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_321),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_321),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_330),
.B(n_185),
.Y(n_451)
);

INVxp33_ASAP7_75t_SL g452 ( 
.A(n_300),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_423),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_R g456 ( 
.A(n_397),
.B(n_330),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_417),
.A2(n_290),
.B1(n_232),
.B2(n_259),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_387),
.B(n_331),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_383),
.B(n_331),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_178),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_L g466 ( 
.A1(n_445),
.A2(n_355),
.B1(n_327),
.B2(n_376),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_423),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_387),
.B(n_332),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_383),
.B(n_332),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_383),
.B(n_335),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_389),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_417),
.B(n_261),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_391),
.B(n_294),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

AOI21x1_ASAP7_75t_L g480 ( 
.A1(n_418),
.A2(n_190),
.B(n_179),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_391),
.B(n_320),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_397),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_299),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_423),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_309),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_445),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_445),
.A2(n_290),
.B1(n_282),
.B2(n_283),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_411),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_410),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_417),
.A2(n_259),
.B1(n_197),
.B2(n_232),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_390),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_199),
.C(n_195),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_445),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_390),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_413),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_413),
.Y(n_502)
);

INVx4_ASAP7_75t_SL g503 ( 
.A(n_411),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_312),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_411),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_424),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_446),
.B(n_317),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_445),
.A2(n_282),
.B1(n_283),
.B2(n_278),
.Y(n_514)
);

INVx8_ASAP7_75t_L g515 ( 
.A(n_445),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_387),
.B(n_335),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_446),
.B(n_351),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_394),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_394),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_394),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_449),
.B(n_351),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_491),
.B(n_499),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_475),
.A2(n_445),
.B1(n_383),
.B2(n_415),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_505),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_484),
.B(n_430),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_491),
.B(n_415),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_476),
.B(n_485),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_507),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_507),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_490),
.B(n_449),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_454),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_484),
.B(n_392),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_516),
.B(n_403),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_501),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_463),
.A2(n_449),
.B1(n_450),
.B2(n_339),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_499),
.B(n_383),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_461),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_444),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_461),
.B(n_438),
.Y(n_545)
);

A2O1A1Ixp33_ASAP7_75t_L g546 ( 
.A1(n_498),
.A2(n_450),
.B(n_422),
.C(n_421),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_515),
.A2(n_418),
.B(n_421),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_457),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_468),
.B(n_450),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_460),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_475),
.B(n_444),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_460),
.B(n_444),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_468),
.B(n_450),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_515),
.A2(n_494),
.B(n_481),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_483),
.B(n_450),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_438),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_462),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_470),
.A2(n_343),
.B1(n_344),
.B2(n_322),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_469),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_469),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_516),
.B(n_403),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_458),
.A2(n_422),
.B1(n_427),
.B2(n_414),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_474),
.B(n_444),
.Y(n_564)
);

O2A1O1Ixp5_ASAP7_75t_L g565 ( 
.A1(n_498),
.A2(n_385),
.B(n_399),
.C(n_395),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_496),
.A2(n_506),
.B1(n_493),
.B2(n_494),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_474),
.B(n_444),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_472),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_471),
.A2(n_399),
.B1(n_405),
.B2(n_392),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_517),
.B(n_441),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_466),
.B(n_441),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_479),
.B(n_395),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_501),
.B(n_438),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_479),
.B(n_448),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_504),
.B(n_441),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_506),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_489),
.B(n_448),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_512),
.B(n_441),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_489),
.B(n_385),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_492),
.A2(n_427),
.B1(n_407),
.B2(n_414),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_502),
.B(n_439),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_495),
.B(n_442),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_L g585 ( 
.A(n_518),
.B(n_412),
.C(n_401),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_495),
.B(n_515),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_523),
.B(n_347),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_502),
.B(n_441),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_457),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_481),
.B(n_384),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_515),
.B(n_442),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_506),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

BUFx5_ASAP7_75t_L g594 ( 
.A(n_508),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_522),
.B(n_401),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_477),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_515),
.A2(n_404),
.B(n_407),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_519),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_477),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_522),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_521),
.A2(n_427),
.B1(n_407),
.B2(n_414),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_514),
.B(n_412),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_455),
.B(n_405),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_473),
.B(n_354),
.Y(n_604)
);

AND2x4_ASAP7_75t_SL g605 ( 
.A(n_516),
.B(n_447),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_519),
.B(n_404),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_493),
.A2(n_407),
.B1(n_414),
.B2(n_404),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_457),
.B(n_261),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_455),
.B(n_439),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_467),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_520),
.B(n_407),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_467),
.B(n_389),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_457),
.B(n_459),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_520),
.B(n_414),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_481),
.A2(n_427),
.B1(n_443),
.B2(n_435),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_521),
.B(n_427),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_488),
.B(n_508),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_481),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_488),
.B(n_432),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_494),
.A2(n_443),
.B1(n_435),
.B2(n_214),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_513),
.B(n_435),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_577),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_554),
.A2(n_494),
.B(n_459),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_531),
.B(n_513),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_568),
.B(n_543),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_536),
.B(n_543),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_577),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_597),
.A2(n_459),
.B(n_457),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_568),
.B(n_503),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_565),
.A2(n_464),
.B(n_432),
.C(n_509),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_538),
.B(n_352),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_592),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_604),
.B(n_300),
.C(n_352),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_613),
.A2(n_459),
.B(n_457),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_613),
.A2(n_465),
.B(n_459),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_538),
.B(n_297),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_592),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_524),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_573),
.B(n_575),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_590),
.A2(n_465),
.B(n_459),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_590),
.A2(n_465),
.B(n_486),
.Y(n_641)
);

OAI21xp33_ASAP7_75t_L g642 ( 
.A1(n_574),
.A2(n_382),
.B(n_381),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_608),
.A2(n_480),
.B(n_464),
.Y(n_643)
);

A2O1A1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_546),
.A2(n_509),
.B(n_511),
.C(n_510),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_542),
.A2(n_465),
.B(n_486),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_526),
.A2(n_465),
.B1(n_215),
.B2(n_298),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_548),
.A2(n_465),
.B(n_486),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_544),
.A2(n_510),
.B(n_509),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_578),
.B(n_510),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_589),
.A2(n_487),
.B(n_486),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_524),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_530),
.B(n_511),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_527),
.A2(n_511),
.B1(n_251),
.B2(n_216),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_600),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_527),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_551),
.A2(n_547),
.B(n_606),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_525),
.A2(n_487),
.B(n_486),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_555),
.A2(n_275),
.B(n_208),
.C(n_277),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_534),
.B(n_482),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_529),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_534),
.B(n_482),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_598),
.B(n_482),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_608),
.A2(n_487),
.B(n_486),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_586),
.A2(n_487),
.B(n_478),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_549),
.A2(n_456),
.B1(n_361),
.B2(n_365),
.Y(n_667)
);

AOI21x1_ASAP7_75t_L g668 ( 
.A1(n_617),
.A2(n_480),
.B(n_478),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_563),
.A2(n_478),
.B(n_477),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_598),
.A2(n_250),
.B(n_226),
.C(n_239),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_609),
.B(n_482),
.Y(n_671)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_574),
.A2(n_382),
.B(n_381),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_563),
.A2(n_566),
.B(n_611),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_618),
.A2(n_487),
.B(n_497),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_535),
.B(n_497),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_529),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_618),
.A2(n_614),
.B(n_616),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_540),
.B(n_356),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_581),
.A2(n_556),
.B(n_545),
.C(n_582),
.Y(n_679)
);

O2A1O1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_553),
.A2(n_437),
.B(n_439),
.C(n_431),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_582),
.B(n_497),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_533),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_533),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_618),
.A2(n_487),
.B(n_500),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_537),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_503),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

AOI21xp33_ASAP7_75t_L g688 ( 
.A1(n_570),
.A2(n_235),
.B(n_437),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_607),
.A2(n_591),
.B(n_552),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_535),
.B(n_500),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_541),
.B(n_556),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_564),
.A2(n_500),
.B(n_400),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_550),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_587),
.A2(n_362),
.B1(n_368),
.B2(n_503),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_550),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_602),
.A2(n_431),
.B(n_436),
.C(n_238),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_557),
.B(n_503),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_609),
.B(n_357),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_600),
.B(n_516),
.Y(n_699)
);

AND2x4_ASAP7_75t_SL g700 ( 
.A(n_583),
.B(n_436),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_567),
.A2(n_400),
.B(n_398),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_610),
.A2(n_400),
.B(n_398),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_558),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_610),
.B(n_357),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_558),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_583),
.B(n_403),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_615),
.A2(n_400),
.B(n_398),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_621),
.A2(n_400),
.B(n_408),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_528),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_601),
.A2(n_416),
.B(n_408),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_605),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_601),
.A2(n_416),
.B(n_408),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_528),
.B(n_503),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_571),
.A2(n_367),
.B1(n_359),
.B2(n_374),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_557),
.B(n_394),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_569),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_595),
.B(n_452),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_682),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_SL g719 ( 
.A(n_636),
.B(n_539),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_709),
.B(n_631),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_639),
.A2(n_673),
.B1(n_572),
.B2(n_681),
.Y(n_721)
);

OAI21xp33_ASAP7_75t_L g722 ( 
.A1(n_642),
.A2(n_360),
.B(n_359),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_698),
.B(n_559),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_682),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_654),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_629),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_711),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_679),
.A2(n_561),
.B1(n_560),
.B2(n_579),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_700),
.B(n_585),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_706),
.B(n_584),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_655),
.B(n_562),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_655),
.B(n_594),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_626),
.B(n_612),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_655),
.B(n_594),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_629),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_704),
.Y(n_736)
);

AOI21x1_ASAP7_75t_L g737 ( 
.A1(n_668),
.A2(n_561),
.B(n_560),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_672),
.B(n_691),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_703),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_646),
.A2(n_576),
.B1(n_588),
.B2(n_619),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_624),
.B(n_638),
.Y(n_741)
);

INVx3_ASAP7_75t_SL g742 ( 
.A(n_699),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_640),
.A2(n_620),
.B(n_603),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_678),
.B(n_360),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_628),
.A2(n_580),
.B(n_569),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_624),
.B(n_594),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_R g747 ( 
.A(n_717),
.B(n_367),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_703),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_651),
.B(n_594),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_667),
.B(n_605),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_659),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_686),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_634),
.A2(n_593),
.B(n_580),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_688),
.A2(n_236),
.B(n_289),
.C(n_599),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_658),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_659),
.Y(n_756)
);

NOR2xp67_ASAP7_75t_L g757 ( 
.A(n_694),
.B(n_369),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_625),
.B(n_594),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_625),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_635),
.A2(n_596),
.B(n_593),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_646),
.B(n_369),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_714),
.B(n_370),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_659),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_686),
.A2(n_594),
.B1(n_370),
.B2(n_374),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_SL g765 ( 
.A1(n_688),
.A2(n_436),
.B(n_428),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_681),
.A2(n_261),
.B1(n_596),
.B2(n_599),
.Y(n_766)
);

O2A1O1Ixp5_ASAP7_75t_L g767 ( 
.A1(n_643),
.A2(n_425),
.B(n_433),
.C(n_429),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_649),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_623),
.A2(n_420),
.B(n_416),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_716),
.Y(n_770)
);

OA22x2_ASAP7_75t_L g771 ( 
.A1(n_713),
.A2(n_278),
.B1(n_285),
.B2(n_288),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_641),
.A2(n_420),
.B(n_594),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_622),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_652),
.B(n_594),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_662),
.B(n_425),
.Y(n_775)
);

OAI22x1_ASAP7_75t_L g776 ( 
.A1(n_676),
.A2(n_285),
.B1(n_188),
.B2(n_288),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_647),
.A2(n_420),
.B(n_261),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_677),
.A2(n_656),
.B(n_645),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_630),
.A2(n_433),
.B(n_429),
.C(n_428),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_683),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_627),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_670),
.A2(n_384),
.B(n_386),
.C(n_393),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_761),
.A2(n_633),
.B(n_660),
.C(n_696),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_773),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_755),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_741),
.B(n_652),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_737),
.A2(n_666),
.B(n_665),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_778),
.A2(n_689),
.B(n_650),
.Y(n_788)
);

OA22x2_ASAP7_75t_L g789 ( 
.A1(n_740),
.A2(n_687),
.B1(n_637),
.B2(n_632),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_781),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_745),
.A2(n_657),
.B(n_669),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_772),
.A2(n_648),
.B(n_692),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_727),
.Y(n_793)
);

OA21x2_ASAP7_75t_L g794 ( 
.A1(n_767),
.A2(n_644),
.B(n_675),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_725),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_721),
.A2(n_697),
.B1(n_671),
.B2(n_685),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_746),
.A2(n_684),
.B(n_674),
.Y(n_797)
);

INVx3_ASAP7_75t_SL g798 ( 
.A(n_725),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_773),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_753),
.A2(n_712),
.B(n_710),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_723),
.B(n_680),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_747),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_721),
.A2(n_715),
.B(n_707),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_770),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_738),
.A2(n_715),
.B(n_681),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_723),
.A2(n_761),
.B1(n_719),
.B2(n_744),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_SL g807 ( 
.A(n_726),
.B(n_693),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_770),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_738),
.B(n_695),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_751),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_780),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_SL g812 ( 
.A(n_747),
.B(n_279),
.C(n_186),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_718),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_775),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_730),
.B(n_705),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_718),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_774),
.A2(n_690),
.B(n_675),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_728),
.A2(n_690),
.B(n_697),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_760),
.A2(n_701),
.B(n_708),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_724),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_736),
.B(n_744),
.Y(n_821)
);

O2A1O1Ixp5_ASAP7_75t_L g822 ( 
.A1(n_731),
.A2(n_664),
.B(n_663),
.C(n_661),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_731),
.B(n_661),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_743),
.A2(n_664),
.B(n_663),
.Y(n_824)
);

AOI21xp33_ASAP7_75t_L g825 ( 
.A1(n_762),
.A2(n_653),
.B(n_281),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_759),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_766),
.A2(n_702),
.B(n_681),
.Y(n_827)
);

AO31x2_ASAP7_75t_L g828 ( 
.A1(n_754),
.A2(n_681),
.A3(n_434),
.B(n_426),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_766),
.A2(n_435),
.B(n_233),
.Y(n_829)
);

AO31x2_ASAP7_75t_L g830 ( 
.A1(n_754),
.A2(n_426),
.A3(n_434),
.B(n_386),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_751),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_752),
.B(n_724),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_732),
.A2(n_435),
.B(n_237),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_775),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_732),
.A2(n_262),
.B(n_240),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_733),
.A2(n_394),
.B(n_393),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_739),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_806),
.A2(n_757),
.B1(n_771),
.B2(n_733),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_784),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_785),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_801),
.A2(n_771),
.B1(n_750),
.B2(n_776),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_821),
.A2(n_764),
.B1(n_729),
.B2(n_742),
.Y(n_842)
);

INVx6_ASAP7_75t_L g843 ( 
.A(n_831),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_790),
.Y(n_844)
);

INVx5_ASAP7_75t_L g845 ( 
.A(n_831),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_815),
.B(n_720),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_799),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_802),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_784),
.Y(n_849)
);

INVx6_ASAP7_75t_L g850 ( 
.A(n_831),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_826),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_799),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_808),
.Y(n_853)
);

CKINVDCx11_ASAP7_75t_R g854 ( 
.A(n_798),
.Y(n_854)
);

BUFx10_ASAP7_75t_L g855 ( 
.A(n_802),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_825),
.A2(n_722),
.B1(n_742),
.B2(n_768),
.Y(n_856)
);

BUFx10_ASAP7_75t_L g857 ( 
.A(n_811),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_786),
.A2(n_752),
.B1(n_751),
.B2(n_756),
.Y(n_858)
);

CKINVDCx11_ASAP7_75t_R g859 ( 
.A(n_798),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_795),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_815),
.B(n_726),
.Y(n_861)
);

BUFx4f_ASAP7_75t_SL g862 ( 
.A(n_795),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_831),
.B(n_751),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_786),
.A2(n_756),
.B1(n_763),
.B2(n_749),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_793),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_814),
.B(n_735),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_805),
.A2(n_756),
.B1(n_763),
.B2(n_758),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_804),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_804),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_816),
.Y(n_870)
);

INVx6_ASAP7_75t_L g871 ( 
.A(n_831),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_834),
.A2(n_756),
.B1(n_763),
.B2(n_735),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_812),
.A2(n_765),
.B1(n_763),
.B2(n_734),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_789),
.A2(n_748),
.B1(n_739),
.B2(n_734),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_793),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_826),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_823),
.B(n_748),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_823),
.B(n_779),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_832),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_783),
.A2(n_279),
.B1(n_281),
.B2(n_284),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_813),
.Y(n_882)
);

BUFx8_ASAP7_75t_L g883 ( 
.A(n_832),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_837),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_816),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_789),
.A2(n_809),
.B1(n_803),
.B2(n_827),
.Y(n_886)
);

INVx8_ASAP7_75t_L g887 ( 
.A(n_810),
.Y(n_887)
);

BUFx4f_ASAP7_75t_SL g888 ( 
.A(n_810),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_810),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_789),
.A2(n_284),
.B1(n_434),
.B2(n_426),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_809),
.A2(n_223),
.B1(n_242),
.B2(n_245),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_820),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_820),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_830),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_807),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_894),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_847),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_879),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_852),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_845),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_876),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_882),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_868),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_869),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_853),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_845),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_838),
.A2(n_796),
.B1(n_836),
.B2(n_818),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_885),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_893),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_886),
.A2(n_788),
.B(n_824),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_886),
.B(n_817),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_839),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_840),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_849),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_838),
.A2(n_794),
.B1(n_829),
.B2(n_835),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_874),
.B(n_828),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_874),
.B(n_828),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_890),
.A2(n_787),
.B(n_819),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_878),
.B(n_828),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_890),
.A2(n_787),
.B(n_819),
.Y(n_920)
);

AO31x2_ASAP7_75t_L g921 ( 
.A1(n_864),
.A2(n_797),
.A3(n_828),
.B(n_777),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_883),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_870),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_892),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_867),
.A2(n_792),
.B(n_791),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_841),
.B(n_828),
.Y(n_926)
);

BUFx2_ASAP7_75t_R g927 ( 
.A(n_865),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_841),
.A2(n_794),
.B1(n_791),
.B2(n_248),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_844),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_884),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_845),
.B(n_830),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_884),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_858),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_916),
.B(n_830),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_898),
.A2(n_856),
.B1(n_881),
.B2(n_842),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_910),
.A2(n_792),
.B(n_800),
.Y(n_936)
);

INVx5_ASAP7_75t_SL g937 ( 
.A(n_931),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_916),
.B(n_917),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_907),
.A2(n_856),
.B(n_891),
.C(n_873),
.Y(n_939)
);

OA21x2_ASAP7_75t_L g940 ( 
.A1(n_910),
.A2(n_800),
.B(n_822),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_927),
.B(n_846),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_898),
.B(n_830),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_896),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_916),
.B(n_830),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_907),
.B(n_891),
.C(n_895),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_907),
.A2(n_877),
.B(n_861),
.C(n_875),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_898),
.B(n_895),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_924),
.B(n_929),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_916),
.B(n_880),
.Y(n_949)
);

NOR2x1_ASAP7_75t_SL g950 ( 
.A(n_900),
.B(n_845),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_928),
.A2(n_862),
.B1(n_851),
.B2(n_866),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_922),
.B(n_848),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_924),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_931),
.Y(n_954)
);

INVx5_ASAP7_75t_SL g955 ( 
.A(n_931),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_SL g956 ( 
.A1(n_930),
.A2(n_872),
.B(n_854),
.C(n_859),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_931),
.B(n_883),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_924),
.B(n_857),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_915),
.A2(n_833),
.B(n_769),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_917),
.B(n_794),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_917),
.B(n_889),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_927),
.B(n_855),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_917),
.B(n_889),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_L g964 ( 
.A(n_928),
.B(n_860),
.C(n_253),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_896),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_929),
.B(n_857),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_922),
.B(n_855),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_915),
.A2(n_782),
.B(n_863),
.Y(n_968)
);

AND2x2_ASAP7_75t_SL g969 ( 
.A(n_911),
.B(n_860),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_910),
.A2(n_887),
.B(n_263),
.C(n_260),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_931),
.B(n_62),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_929),
.B(n_843),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_SL g973 ( 
.A1(n_930),
.A2(n_862),
.B(n_888),
.C(n_6),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_954),
.B(n_931),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_938),
.B(n_925),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_938),
.B(n_925),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_948),
.B(n_911),
.Y(n_977)
);

INVxp33_ASAP7_75t_L g978 ( 
.A(n_952),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_939),
.A2(n_926),
.B1(n_922),
.B2(n_911),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_947),
.B(n_930),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_954),
.B(n_925),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_954),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_943),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_943),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_943),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_947),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_965),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_965),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_960),
.B(n_929),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_960),
.B(n_913),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_945),
.A2(n_964),
.B1(n_935),
.B2(n_969),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_954),
.B(n_925),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_972),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_953),
.B(n_913),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_972),
.B(n_931),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_934),
.B(n_897),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_953),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_953),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_993),
.B(n_937),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_974),
.B(n_950),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_991),
.A2(n_964),
.B1(n_969),
.B2(n_945),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_982),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_974),
.B(n_950),
.Y(n_1003)
);

AOI211xp5_ASAP7_75t_L g1004 ( 
.A1(n_979),
.A2(n_973),
.B(n_951),
.C(n_956),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_993),
.B(n_937),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_987),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_987),
.Y(n_1007)
);

AOI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_979),
.A2(n_951),
.B(n_970),
.C(n_946),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_982),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_991),
.A2(n_969),
.B1(n_949),
.B2(n_941),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_987),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_974),
.B(n_971),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_980),
.B(n_986),
.C(n_977),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_993),
.B(n_937),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_986),
.Y(n_1015)
);

AOI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_980),
.A2(n_949),
.B1(n_966),
.B2(n_958),
.C(n_913),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_989),
.B(n_942),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_978),
.A2(n_971),
.B1(n_957),
.B2(n_967),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_975),
.B(n_937),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1000),
.B(n_975),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_1015),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1007),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_1013),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1007),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_1010),
.B(n_978),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1006),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1017),
.B(n_977),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1016),
.B(n_990),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1000),
.B(n_975),
.Y(n_1029)
);

NOR2xp67_ASAP7_75t_L g1030 ( 
.A(n_1009),
.B(n_984),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_1025),
.A2(n_1001),
.B(n_1010),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1020),
.B(n_1000),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1021),
.B(n_976),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1023),
.B(n_989),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_1023),
.B(n_990),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_1020),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1026),
.Y(n_1037)
);

OAI21xp33_ASAP7_75t_L g1038 ( 
.A1(n_1031),
.A2(n_1025),
.B(n_1028),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1031),
.B(n_1027),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1032),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1036),
.B(n_1029),
.Y(n_1041)
);

AOI31xp33_ASAP7_75t_L g1042 ( 
.A1(n_1038),
.A2(n_1004),
.A3(n_1008),
.B(n_962),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1039),
.B(n_1035),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1039),
.A2(n_1040),
.B(n_1034),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1041),
.A2(n_1018),
.B1(n_1033),
.B2(n_1030),
.Y(n_1045)
);

AOI21xp33_ASAP7_75t_SL g1046 ( 
.A1(n_1038),
.A2(n_1018),
.B(n_1037),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1039),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1038),
.A2(n_1000),
.B1(n_1003),
.B2(n_1012),
.Y(n_1048)
);

AOI211xp5_ASAP7_75t_SL g1049 ( 
.A1(n_1038),
.A2(n_971),
.B(n_1003),
.C(n_926),
.Y(n_1049)
);

NAND2xp33_ASAP7_75t_SL g1050 ( 
.A(n_1039),
.B(n_1002),
.Y(n_1050)
);

AOI222xp33_ASAP7_75t_L g1051 ( 
.A1(n_1038),
.A2(n_922),
.B1(n_976),
.B2(n_1002),
.C1(n_1003),
.C2(n_1029),
.Y(n_1051)
);

AOI222xp33_ASAP7_75t_L g1052 ( 
.A1(n_1038),
.A2(n_976),
.B1(n_1003),
.B2(n_959),
.C1(n_1012),
.C2(n_1009),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1047),
.B(n_1022),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1043),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1042),
.B(n_1022),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_SL g1056 ( 
.A1(n_1046),
.A2(n_1012),
.B(n_971),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_1045),
.B(n_1009),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_1050),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1044),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1052),
.A2(n_1012),
.B(n_1019),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_1048),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1051),
.A2(n_957),
.B1(n_1019),
.B2(n_992),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1049),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1047),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_1042),
.A2(n_992),
.B(n_981),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1042),
.A2(n_1024),
.B1(n_997),
.B2(n_998),
.C(n_1011),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_1047),
.B(n_887),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_1047),
.B(n_887),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1058),
.A2(n_959),
.B(n_994),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1061),
.A2(n_957),
.B1(n_981),
.B2(n_992),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1054),
.B(n_1064),
.Y(n_1072)
);

AOI21xp33_ASAP7_75t_L g1073 ( 
.A1(n_1055),
.A2(n_4),
.B(n_5),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1053),
.Y(n_1074)
);

OAI21xp33_ASAP7_75t_SL g1075 ( 
.A1(n_1057),
.A2(n_1005),
.B(n_999),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1067),
.B(n_999),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_1067),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1063),
.B(n_1005),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1056),
.B(n_1014),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_1068),
.Y(n_1080)
);

OAI221xp5_ASAP7_75t_L g1081 ( 
.A1(n_1060),
.A2(n_1062),
.B1(n_1066),
.B2(n_1065),
.C(n_1068),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1059),
.B(n_1014),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1058),
.A2(n_957),
.B1(n_981),
.B2(n_1009),
.Y(n_1083)
);

OAI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1058),
.A2(n_1009),
.B(n_968),
.C(n_926),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1064),
.Y(n_1085)
);

XOR2x2_ASAP7_75t_L g1086 ( 
.A(n_1058),
.B(n_4),
.Y(n_1086)
);

NOR2x1p5_ASAP7_75t_L g1087 ( 
.A(n_1059),
.B(n_932),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1073),
.B(n_1006),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_1077),
.B(n_968),
.C(n_932),
.Y(n_1089)
);

OAI211xp5_ASAP7_75t_SL g1090 ( 
.A1(n_1080),
.A2(n_1073),
.B(n_1074),
.C(n_1081),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1085),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1086),
.B(n_1011),
.Y(n_1092)
);

NOR3x1_ASAP7_75t_L g1093 ( 
.A(n_1078),
.B(n_982),
.C(n_997),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_L g1094 ( 
.A(n_1072),
.B(n_5),
.Y(n_1094)
);

NOR4xp25_ASAP7_75t_L g1095 ( 
.A(n_1084),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_L g1096 ( 
.A(n_1071),
.B(n_1009),
.C(n_932),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1076),
.B(n_995),
.Y(n_1097)
);

NAND3xp33_ASAP7_75t_SL g1098 ( 
.A(n_1083),
.B(n_255),
.C(n_249),
.Y(n_1098)
);

NAND4xp75_ASAP7_75t_L g1099 ( 
.A(n_1069),
.B(n_906),
.C(n_900),
.D(n_998),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_SL g1100 ( 
.A(n_1070),
.B(n_258),
.C(n_257),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1082),
.B(n_995),
.Y(n_1101)
);

NAND4xp25_ASAP7_75t_SL g1102 ( 
.A(n_1075),
.B(n_994),
.C(n_926),
.D(n_963),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1079),
.B(n_932),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_1087),
.B(n_266),
.C(n_264),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1095),
.A2(n_269),
.B1(n_933),
.B2(n_905),
.C(n_988),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_SL g1106 ( 
.A(n_1094),
.B(n_888),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1092),
.Y(n_1107)
);

AOI322xp5_ASAP7_75t_L g1108 ( 
.A1(n_1091),
.A2(n_961),
.A3(n_963),
.B1(n_996),
.B2(n_974),
.C1(n_944),
.C2(n_934),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_L g1109 ( 
.A1(n_1090),
.A2(n_933),
.B1(n_905),
.B2(n_988),
.C(n_985),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_L g1110 ( 
.A(n_1104),
.B(n_10),
.Y(n_1110)
);

NAND4xp75_ASAP7_75t_L g1111 ( 
.A(n_1093),
.B(n_900),
.C(n_906),
.D(n_12),
.Y(n_1111)
);

OAI211xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1103),
.A2(n_10),
.B(n_11),
.C(n_14),
.Y(n_1112)
);

AOI211xp5_ASAP7_75t_L g1113 ( 
.A1(n_1100),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_1113)
);

NOR3xp33_ASAP7_75t_L g1114 ( 
.A(n_1098),
.B(n_933),
.C(n_15),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1096),
.A2(n_955),
.B1(n_937),
.B2(n_974),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1088),
.A2(n_905),
.B(n_906),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_1088),
.A2(n_17),
.B(n_19),
.Y(n_1117)
);

NAND4xp25_ASAP7_75t_L g1118 ( 
.A(n_1089),
.B(n_1101),
.C(n_1097),
.D(n_1102),
.Y(n_1118)
);

AOI211xp5_ASAP7_75t_L g1119 ( 
.A1(n_1099),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1090),
.A2(n_906),
.B(n_900),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1090),
.B(n_20),
.Y(n_1121)
);

OAI211xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1091),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1094),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1090),
.B(n_24),
.Y(n_1124)
);

AOI211x1_ASAP7_75t_SL g1125 ( 
.A1(n_1090),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_1125)
);

AOI31xp33_ASAP7_75t_L g1126 ( 
.A1(n_1094),
.A2(n_863),
.A3(n_28),
.B(n_29),
.Y(n_1126)
);

OAI31xp33_ASAP7_75t_L g1127 ( 
.A1(n_1090),
.A2(n_26),
.A3(n_30),
.B(n_31),
.Y(n_1127)
);

NAND4xp25_ASAP7_75t_L g1128 ( 
.A(n_1090),
.B(n_942),
.C(n_995),
.D(n_961),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1123),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1121),
.A2(n_30),
.B(n_31),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1124),
.A2(n_957),
.B1(n_955),
.B2(n_944),
.Y(n_1131)
);

AO22x2_ASAP7_75t_SL g1132 ( 
.A1(n_1114),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1132)
);

OAI211xp5_ASAP7_75t_L g1133 ( 
.A1(n_1127),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_1133)
);

AO22x2_ASAP7_75t_L g1134 ( 
.A1(n_1107),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1134)
);

AO22x1_ASAP7_75t_L g1135 ( 
.A1(n_1125),
.A2(n_957),
.B1(n_40),
.B2(n_41),
.Y(n_1135)
);

AOI211xp5_ASAP7_75t_L g1136 ( 
.A1(n_1105),
.A2(n_39),
.B(n_40),
.C(n_43),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1117),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1106),
.A2(n_957),
.B1(n_995),
.B2(n_996),
.Y(n_1138)
);

CKINVDCx6p67_ASAP7_75t_R g1139 ( 
.A(n_1126),
.Y(n_1139)
);

AOI211xp5_ASAP7_75t_L g1140 ( 
.A1(n_1112),
.A2(n_43),
.B(n_44),
.C(n_46),
.Y(n_1140)
);

NOR2x1p5_ASAP7_75t_L g1141 ( 
.A(n_1111),
.B(n_44),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1117),
.Y(n_1142)
);

AOI222xp33_ASAP7_75t_L g1143 ( 
.A1(n_1109),
.A2(n_1122),
.B1(n_1110),
.B2(n_1115),
.C1(n_1128),
.C2(n_1119),
.Y(n_1143)
);

OA22x2_ASAP7_75t_L g1144 ( 
.A1(n_1118),
.A2(n_984),
.B1(n_995),
.B2(n_985),
.Y(n_1144)
);

AOI211xp5_ASAP7_75t_L g1145 ( 
.A1(n_1120),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1113),
.A2(n_955),
.B1(n_983),
.B2(n_996),
.Y(n_1146)
);

OAI211xp5_ASAP7_75t_L g1147 ( 
.A1(n_1116),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1108),
.Y(n_1148)
);

OAI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1127),
.A2(n_983),
.B1(n_54),
.B2(n_55),
.C(n_56),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_L g1150 ( 
.A(n_1127),
.B(n_53),
.C(n_58),
.Y(n_1150)
);

OAI211xp5_ASAP7_75t_SL g1151 ( 
.A1(n_1127),
.A2(n_59),
.B(n_60),
.C(n_919),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1127),
.B(n_59),
.C(n_60),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_L g1153 ( 
.A(n_1142),
.B(n_899),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_1137),
.B(n_66),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1137),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1139),
.B(n_996),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1134),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1131),
.A2(n_955),
.B1(n_899),
.B2(n_901),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1135),
.B(n_996),
.Y(n_1159)
);

NAND4xp75_ASAP7_75t_L g1160 ( 
.A(n_1129),
.B(n_940),
.C(n_901),
.D(n_899),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1141),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1132),
.B(n_901),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_1134),
.Y(n_1163)
);

AND2x2_ASAP7_75t_SL g1164 ( 
.A(n_1148),
.B(n_940),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1140),
.B(n_1130),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1144),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1133),
.B(n_897),
.Y(n_1167)
);

NOR2x1p5_ASAP7_75t_L g1168 ( 
.A(n_1150),
.B(n_903),
.Y(n_1168)
);

AND3x4_ASAP7_75t_L g1169 ( 
.A(n_1151),
.B(n_897),
.C(n_902),
.Y(n_1169)
);

NOR2x1_ASAP7_75t_L g1170 ( 
.A(n_1152),
.B(n_70),
.Y(n_1170)
);

XNOR2x1_ASAP7_75t_L g1171 ( 
.A(n_1146),
.B(n_71),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_1147),
.B(n_72),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1149),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1138),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1163),
.B(n_1143),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1157),
.B(n_1145),
.Y(n_1176)
);

AOI221xp5_ASAP7_75t_L g1177 ( 
.A1(n_1166),
.A2(n_1136),
.B1(n_903),
.B2(n_904),
.C(n_897),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1161),
.B(n_902),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1154),
.B(n_1155),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1170),
.B(n_955),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_L g1181 ( 
.A(n_1173),
.B(n_919),
.C(n_904),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1157),
.B(n_902),
.Y(n_1182)
);

NOR3x1_ASAP7_75t_L g1183 ( 
.A(n_1165),
.B(n_78),
.C(n_79),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1156),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1172),
.B(n_902),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1153),
.Y(n_1186)
);

OAI211xp5_ASAP7_75t_L g1187 ( 
.A1(n_1174),
.A2(n_904),
.B(n_903),
.C(n_940),
.Y(n_1187)
);

NOR2x1p5_ASAP7_75t_L g1188 ( 
.A(n_1162),
.B(n_909),
.Y(n_1188)
);

OAI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1159),
.A2(n_1167),
.B1(n_1171),
.B2(n_1158),
.C(n_1169),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1175),
.B(n_1164),
.C(n_1168),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1176),
.A2(n_1160),
.B(n_908),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1179),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1184),
.B(n_909),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1180),
.A2(n_843),
.B1(n_850),
.B2(n_871),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1189),
.A2(n_908),
.B(n_909),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1177),
.A2(n_909),
.B1(n_908),
.B2(n_896),
.C(n_912),
.Y(n_1196)
);

XOR2xp5_ASAP7_75t_L g1197 ( 
.A(n_1179),
.B(n_80),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1186),
.A2(n_843),
.B1(n_850),
.B2(n_871),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1183),
.Y(n_1199)
);

OAI221xp5_ASAP7_75t_L g1200 ( 
.A1(n_1182),
.A2(n_850),
.B1(n_871),
.B2(n_908),
.C(n_919),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1178),
.A2(n_919),
.B1(n_923),
.B2(n_914),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1188),
.A2(n_923),
.B1(n_914),
.B2(n_912),
.Y(n_1202)
);

AO22x2_ASAP7_75t_L g1203 ( 
.A1(n_1185),
.A2(n_923),
.B1(n_914),
.B2(n_912),
.Y(n_1203)
);

NAND4xp25_ASAP7_75t_L g1204 ( 
.A(n_1181),
.B(n_81),
.C(n_83),
.D(n_86),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1192),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1190),
.A2(n_1187),
.B1(n_923),
.B2(n_914),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1199),
.A2(n_912),
.B1(n_940),
.B2(n_936),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_1197),
.A2(n_88),
.B1(n_89),
.B2(n_94),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1193),
.Y(n_1209)
);

AO22x2_ASAP7_75t_L g1210 ( 
.A1(n_1198),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_1210)
);

OAI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1204),
.A2(n_1191),
.B1(n_1194),
.B2(n_1195),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1200),
.A2(n_936),
.B1(n_920),
.B2(n_918),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1196),
.A2(n_936),
.B1(n_920),
.B2(n_918),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1201),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_1214)
);

XNOR2xp5_ASAP7_75t_L g1215 ( 
.A(n_1205),
.B(n_1203),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1209),
.A2(n_1202),
.B(n_1203),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1208),
.A2(n_108),
.B(n_114),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1211),
.B(n_921),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1210),
.B(n_115),
.Y(n_1219)
);

XOR2xp5_ASAP7_75t_L g1220 ( 
.A(n_1214),
.B(n_116),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1217),
.Y(n_1221)
);

AO22x2_ASAP7_75t_L g1222 ( 
.A1(n_1220),
.A2(n_1206),
.B1(n_1212),
.B2(n_1207),
.Y(n_1222)
);

XOR2xp5_ASAP7_75t_L g1223 ( 
.A(n_1220),
.B(n_1213),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1215),
.A2(n_117),
.B(n_119),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1221),
.A2(n_1219),
.B(n_1216),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1225),
.A2(n_1224),
.B(n_1223),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1226),
.A2(n_1218),
.B(n_1222),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1227),
.A2(n_120),
.B(n_121),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1228),
.A2(n_127),
.B1(n_128),
.B2(n_132),
.C(n_133),
.Y(n_1229)
);

AOI211xp5_ASAP7_75t_L g1230 ( 
.A1(n_1229),
.A2(n_135),
.B(n_137),
.C(n_144),
.Y(n_1230)
);


endmodule