module fake_jpeg_20993_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_39),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_41),
.B(n_46),
.Y(n_105)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_53),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx6p67_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_7),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_67),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_23),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_7),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_9),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_40),
.A2(n_28),
.B1(n_36),
.B2(n_35),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_83),
.A2(n_101),
.B1(n_103),
.B2(n_109),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_28),
.B1(n_36),
.B2(n_23),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_102),
.B1(n_67),
.B2(n_68),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_28),
.B1(n_36),
.B2(n_32),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_92),
.A2(n_106),
.B1(n_39),
.B2(n_46),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_28),
.B1(n_36),
.B2(n_35),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_23),
.B1(n_35),
.B2(n_34),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_37),
.B1(n_34),
.B2(n_26),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_38),
.A2(n_37),
.B1(n_34),
.B2(n_26),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_56),
.A2(n_14),
.B(n_13),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_87),
.B(n_79),
.C(n_105),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_53),
.A2(n_37),
.B1(n_26),
.B2(n_29),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_115),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_49),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_116),
.B(n_119),
.Y(n_177)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_152),
.Y(n_157)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_127),
.Y(n_156)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_23),
.B1(n_104),
.B2(n_29),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_126),
.B(n_140),
.Y(n_188)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_70),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_133),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_59),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_132),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_107),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_57),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_42),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_76),
.C(n_50),
.Y(n_161)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_149),
.B1(n_155),
.B2(n_78),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_86),
.B(n_29),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_94),
.A2(n_31),
.B(n_33),
.C(n_25),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_50),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_90),
.B(n_31),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_78),
.B1(n_30),
.B2(n_21),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_80),
.A2(n_47),
.B1(n_69),
.B2(n_65),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_74),
.A2(n_31),
.B1(n_33),
.B2(n_25),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_74),
.B(n_33),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_153),
.A2(n_154),
.B1(n_78),
.B2(n_86),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_77),
.B(n_50),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_80),
.A2(n_69),
.B1(n_66),
.B2(n_65),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_113),
.B1(n_85),
.B2(n_95),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_167),
.B1(n_174),
.B2(n_182),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_10),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_193),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_165),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_100),
.B1(n_77),
.B2(n_95),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_168),
.B(n_135),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_117),
.A2(n_113),
.B1(n_85),
.B2(n_96),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_179),
.A2(n_186),
.B1(n_139),
.B2(n_136),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_43),
.B1(n_66),
.B2(n_64),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_117),
.A2(n_51),
.B1(n_64),
.B2(n_43),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_191),
.B1(n_14),
.B2(n_1),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_128),
.A2(n_30),
.B1(n_21),
.B2(n_96),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_189),
.B1(n_137),
.B2(n_123),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_44),
.C(n_51),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_155),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_140),
.B1(n_130),
.B2(n_150),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_143),
.A2(n_30),
.B1(n_21),
.B2(n_55),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_129),
.A2(n_119),
.B1(n_126),
.B2(n_134),
.Y(n_191)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_52),
.B1(n_44),
.B2(n_111),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_195),
.A2(n_200),
.B1(n_202),
.B2(n_204),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_197),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_156),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_164),
.A2(n_149),
.B1(n_127),
.B2(n_142),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_148),
.B(n_135),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_206),
.B(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_124),
.B1(n_137),
.B2(n_118),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_209),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_120),
.B1(n_52),
.B2(n_121),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_208),
.A2(n_214),
.B1(n_220),
.B2(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_121),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_191),
.B(n_161),
.CI(n_172),
.CON(n_210),
.SN(n_210)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_210),
.B(n_212),
.Y(n_266)
);

AO21x2_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_151),
.B(n_131),
.Y(n_211)
);

AO21x2_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_166),
.B(n_183),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_188),
.B(n_11),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_115),
.B(n_114),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_157),
.A2(n_193),
.B1(n_185),
.B2(n_167),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_135),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_221),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_32),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_225),
.B1(n_175),
.B2(n_159),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_162),
.A2(n_9),
.B(n_13),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_218),
.A2(n_219),
.B(n_222),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_178),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_6),
.B1(n_12),
.B2(n_10),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_5),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_9),
.B(n_12),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_SL g223 ( 
.A(n_170),
.B(n_4),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_228),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_169),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_158),
.A2(n_4),
.B1(n_10),
.B2(n_12),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_233),
.B1(n_187),
.B2(n_181),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_169),
.B(n_0),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_0),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_0),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_174),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

AO21x2_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_211),
.B(n_208),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_192),
.C(n_173),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_246),
.C(n_253),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g239 ( 
.A(n_223),
.B(n_159),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_265),
.C(n_219),
.Y(n_279)
);

NAND2x1_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_180),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_202),
.B(n_226),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_203),
.B1(n_207),
.B2(n_211),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_245),
.B1(n_262),
.B2(n_233),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_192),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_252),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_198),
.A2(n_206),
.B1(n_187),
.B2(n_217),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_196),
.B1(n_222),
.B2(n_166),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_173),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_190),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_180),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_264),
.C(n_228),
.Y(n_298)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_207),
.A2(n_181),
.B1(n_166),
.B2(n_2),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_199),
.B(n_166),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_225),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_224),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_269),
.A2(n_236),
.B(n_267),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_211),
.B1(n_214),
.B2(n_195),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_288),
.B1(n_297),
.B2(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_275),
.A2(n_282),
.B1(n_293),
.B2(n_257),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_277),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_215),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_279),
.A2(n_265),
.B1(n_218),
.B2(n_249),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_281),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_232),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_220),
.B1(n_211),
.B2(n_197),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_240),
.B(n_221),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_285),
.Y(n_301)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_291),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_261),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_287),
.Y(n_309)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_212),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_263),
.B1(n_241),
.B2(n_254),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_229),
.Y(n_294)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_259),
.A2(n_211),
.B1(n_228),
.B2(n_227),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_302),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_236),
.B(n_267),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_285),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_316),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_317),
.B1(n_319),
.B2(n_323),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_264),
.C(n_246),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_312),
.C(n_320),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_311),
.B(n_319),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_298),
.C(n_252),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_255),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_289),
.A2(n_237),
.B1(n_266),
.B2(n_238),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_237),
.B1(n_260),
.B2(n_250),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_276),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_282),
.A2(n_266),
.B1(n_235),
.B2(n_256),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_278),
.B(n_256),
.C(n_1),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_275),
.A2(n_1),
.B1(n_2),
.B2(n_293),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_277),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_326),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_280),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_327),
.A2(n_303),
.B(n_301),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_274),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_336),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_291),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_337),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_341),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_297),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_311),
.B(n_281),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_343),
.A2(n_315),
.B1(n_276),
.B2(n_273),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_318),
.B(n_300),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_349),
.B(n_350),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_317),
.C(n_320),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_355),
.C(n_344),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_310),
.C(n_315),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_356),
.Y(n_362)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_299),
.B1(n_300),
.B2(n_292),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_306),
.Y(n_366)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_360),
.Y(n_365)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_346),
.C(n_344),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_345),
.B(n_325),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_364),
.B(n_351),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_366),
.A2(n_356),
.B1(n_354),
.B2(n_352),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_349),
.A2(n_330),
.B1(n_324),
.B2(n_314),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_371),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_331),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_347),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_350),
.A2(n_292),
.B(n_341),
.Y(n_371)
);

XOR2x2_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_335),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_355),
.Y(n_377)
);

INVx11_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_361),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_376),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_379),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_370),
.A2(n_354),
.B(n_352),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_378),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_363),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_305),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_383),
.B(n_371),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_381),
.B(n_385),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_384),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_276),
.B1(n_334),
.B2(n_360),
.Y(n_384)
);

AOI21x1_ASAP7_75t_SL g398 ( 
.A1(n_387),
.A2(n_365),
.B(n_362),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_346),
.C(n_368),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_390),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_380),
.A2(n_369),
.B(n_374),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_382),
.A2(n_365),
.B1(n_373),
.B2(n_369),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_367),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_389),
.B(n_358),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_397),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_276),
.B(n_386),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_388),
.B(n_353),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_399),
.A2(n_391),
.B(n_392),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_362),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_386),
.C(n_387),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_401),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_402),
.A2(n_403),
.B(n_396),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_405),
.A2(n_404),
.B1(n_398),
.B2(n_329),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_406),
.B(n_323),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_329),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_2),
.Y(n_410)
);


endmodule