module fake_netlist_6_2316_n_1764 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1764);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1764;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_34),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_24),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_32),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_37),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_45),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_55),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_93),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_123),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_40),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_51),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_37),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_78),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_127),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_79),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_24),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_148),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_75),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_99),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_3),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_28),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_18),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_48),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_100),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_53),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_50),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_18),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_48),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_88),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_92),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_105),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_110),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_134),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_122),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_44),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_63),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_89),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_66),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_83),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_41),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_91),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_47),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_46),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_107),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_74),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_82),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_65),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_46),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_14),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_7),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_87),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_104),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_146),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_121),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_60),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_84),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_43),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_31),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_62),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_85),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_80),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_5),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_109),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_4),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_14),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_40),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_41),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_86),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_59),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_54),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_50),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_28),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_95),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_67),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_139),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_23),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_117),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_51),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_35),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_64),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_33),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_30),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_3),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_17),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_10),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_7),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_25),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_9),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_58),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_126),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_2),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_23),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_152),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_124),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_76),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_20),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_6),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_17),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_15),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_57),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_138),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_6),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_25),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_90),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_34),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_118),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_72),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_33),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_111),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_130),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_9),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_4),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_115),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_133),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_71),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_184),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_159),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_201),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_0),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_188),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_201),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_185),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_201),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_162),
.B(n_178),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_201),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_201),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_276),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_172),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_179),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_217),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_187),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_226),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_193),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_218),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_190),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_226),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_194),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_198),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_199),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_226),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_205),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_214),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_193),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_0),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_206),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_208),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_209),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_226),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_210),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_221),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_160),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_160),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_179),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_259),
.B(n_1),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_219),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_251),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_196),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_211),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_213),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_261),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_212),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_174),
.B(n_1),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_263),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_196),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_227),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_235),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_301),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_174),
.B(n_8),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_212),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_232),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_232),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_295),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_234),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_163),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_177),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_245),
.B(n_8),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_245),
.B(n_10),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_236),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_256),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_197),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_223),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_250),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_255),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_256),
.B(n_11),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_155),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_237),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_310),
.B(n_216),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_315),
.A2(n_270),
.B(n_260),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_216),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_335),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_318),
.B(n_266),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_157),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_326),
.B(n_336),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_157),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_381),
.B(n_179),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_161),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_333),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_341),
.B(n_362),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_376),
.B(n_166),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_358),
.B(n_173),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_311),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_350),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_311),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_371),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_347),
.B(n_179),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_358),
.B(n_191),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_364),
.B(n_165),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_368),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_337),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_377),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_312),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_364),
.B(n_165),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_365),
.B(n_204),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_319),
.B(n_309),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_380),
.B(n_347),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_388),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_441),
.B(n_348),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_390),
.B(n_179),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_308),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_404),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_412),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_412),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_398),
.B(n_314),
.Y(n_464)
);

INVxp33_ASAP7_75t_SL g465 ( 
.A(n_448),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_405),
.B(n_356),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_398),
.B(n_348),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_405),
.B(n_324),
.Y(n_468)
);

OR2x2_ASAP7_75t_SL g469 ( 
.A(n_426),
.B(n_361),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_437),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_409),
.A2(n_287),
.B1(n_268),
.B2(n_277),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_426),
.B(n_361),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_389),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_413),
.B(n_328),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_413),
.B(n_330),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_407),
.B(n_331),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_389),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_407),
.B(n_332),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_390),
.A2(n_374),
.B1(n_373),
.B2(n_283),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_413),
.B(n_334),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_413),
.B(n_338),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_400),
.B(n_339),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_413),
.B(n_340),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_413),
.B(n_342),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_390),
.B(n_352),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_390),
.B(n_215),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_384),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_429),
.B(n_353),
.Y(n_502)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_415),
.Y(n_503)
);

BUFx4f_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_409),
.A2(n_383),
.B1(n_375),
.B2(n_359),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_415),
.B(n_170),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_400),
.B(n_366),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_448),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_384),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_415),
.B(n_229),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_384),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_386),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_386),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_386),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_387),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_415),
.B(n_215),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_421),
.B(n_281),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_399),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_423),
.B(n_433),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_387),
.Y(n_521)
);

AO22x2_ASAP7_75t_L g522 ( 
.A1(n_421),
.A2(n_249),
.B1(n_282),
.B2(n_274),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_389),
.Y(n_523)
);

AND3x2_ASAP7_75t_L g524 ( 
.A(n_429),
.B(n_304),
.C(n_228),
.Y(n_524)
);

AND3x2_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_207),
.C(n_248),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_423),
.B(n_366),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_423),
.B(n_367),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_421),
.B(n_306),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_421),
.A2(n_289),
.B1(n_278),
.B2(n_230),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_432),
.B(n_215),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_389),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_387),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_391),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_391),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_418),
.B(n_238),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_418),
.B(n_240),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_432),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_431),
.B(n_439),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_423),
.B(n_380),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_439),
.B(n_367),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_392),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_432),
.B(n_215),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_394),
.B(n_164),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_394),
.B(n_369),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_392),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_392),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_418),
.B(n_432),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_399),
.B(n_215),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_435),
.B(n_164),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_397),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_433),
.A2(n_239),
.B1(n_230),
.B2(n_298),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_397),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_389),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_435),
.B(n_164),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_448),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_397),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_401),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_389),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_399),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_443),
.B(n_369),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_438),
.B(n_230),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_401),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_389),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_433),
.A2(n_230),
.B1(n_239),
.B2(n_298),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_401),
.Y(n_567)
);

INVx8_ASAP7_75t_L g568 ( 
.A(n_432),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_406),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_432),
.B(n_230),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_406),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_438),
.B(n_239),
.Y(n_572)
);

INVx6_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_444),
.B(n_370),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_406),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_408),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_444),
.A2(n_239),
.B1(n_298),
.B2(n_370),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_408),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_443),
.B(n_202),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_444),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_444),
.B(n_243),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_451),
.B(n_202),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_447),
.B(n_202),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_408),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_451),
.B(n_225),
.Y(n_586)
);

BUFx4f_ASAP7_75t_L g587 ( 
.A(n_438),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_452),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_410),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_410),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_410),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_450),
.A2(n_239),
.B1(n_298),
.B2(n_299),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_SL g593 ( 
.A(n_452),
.B(n_181),
.C(n_303),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_411),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_452),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_451),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_389),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_438),
.B(n_225),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_450),
.A2(n_449),
.B1(n_436),
.B2(n_442),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_411),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_411),
.Y(n_601)
);

BUFx8_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

INVx8_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_573),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_470),
.B(n_320),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_490),
.B(n_167),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_519),
.B(n_450),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_481),
.B(n_167),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_560),
.B(n_450),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_503),
.B(n_450),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_573),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_509),
.B(n_156),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_486),
.A2(n_343),
.B1(n_323),
.B2(n_354),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_450),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_459),
.B(n_168),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_573),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_453),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_573),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_596),
.B(n_327),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_503),
.B(n_438),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_468),
.B(n_168),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_453),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_507),
.B(n_438),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_498),
.B(n_169),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_508),
.B(n_156),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_464),
.B(n_349),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_538),
.B(n_298),
.Y(n_630)
);

BUFx5_ASAP7_75t_L g631 ( 
.A(n_456),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_456),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_538),
.B(n_438),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_506),
.B(n_511),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_548),
.B(n_438),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_473),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_SL g637 ( 
.A(n_538),
.B(n_473),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_520),
.B(n_416),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_581),
.B(n_436),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_517),
.B(n_244),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_545),
.B(n_169),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_581),
.A2(n_357),
.B1(n_254),
.B2(n_257),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_522),
.A2(n_449),
.B1(n_442),
.B2(n_436),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_535),
.B(n_171),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_454),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_454),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_520),
.B(n_416),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_518),
.B(n_171),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_561),
.B(n_416),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_537),
.B(n_417),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_466),
.B(n_417),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_466),
.B(n_478),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_466),
.B(n_417),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_455),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_501),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_466),
.B(n_430),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_540),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_564),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_479),
.B(n_430),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_488),
.B(n_430),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_528),
.A2(n_264),
.B1(n_307),
.B2(n_175),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_510),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_576),
.B(n_457),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_489),
.A2(n_497),
.B1(n_494),
.B2(n_540),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_540),
.B(n_430),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_502),
.B(n_175),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_526),
.B(n_434),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_526),
.B(n_434),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_455),
.Y(n_670)
);

AND2x6_ASAP7_75t_SL g671 ( 
.A(n_465),
.B(n_275),
.Y(n_671)
);

BUFx8_ASAP7_75t_L g672 ( 
.A(n_463),
.Y(n_672)
);

AND2x6_ASAP7_75t_L g673 ( 
.A(n_474),
.B(n_296),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_517),
.B(n_176),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_505),
.B(n_176),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_527),
.B(n_574),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_584),
.B(n_463),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_460),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_584),
.B(n_442),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_510),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_472),
.B(n_182),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_564),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_517),
.B(n_182),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_527),
.B(n_434),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_593),
.B(n_449),
.C(n_183),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_460),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_550),
.B(n_183),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_582),
.B(n_269),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_574),
.B(n_434),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_555),
.B(n_269),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_580),
.B(n_280),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_474),
.B(n_440),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_477),
.B(n_440),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_477),
.B(n_440),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_564),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_515),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_568),
.A2(n_385),
.B(n_445),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_483),
.B(n_485),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_461),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_522),
.A2(n_424),
.B1(n_425),
.B2(n_158),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_525),
.B(n_424),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_483),
.B(n_440),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_471),
.B(n_271),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_467),
.B(n_280),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_521),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_485),
.B(n_491),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_487),
.A2(n_286),
.B1(n_302),
.B2(n_284),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_517),
.B(n_284),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_461),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_521),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_462),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_476),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_583),
.B(n_424),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_462),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_529),
.A2(n_302),
.B1(n_286),
.B2(n_292),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_586),
.B(n_285),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_471),
.B(n_285),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_517),
.A2(n_292),
.B1(n_305),
.B2(n_446),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_517),
.A2(n_305),
.B1(n_445),
.B2(n_446),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_491),
.B(n_428),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_524),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_544),
.B(n_225),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_469),
.B(n_186),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_517),
.A2(n_446),
.B1(n_445),
.B2(n_385),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_532),
.B(n_445),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_532),
.B(n_446),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_522),
.A2(n_385),
.B1(n_425),
.B2(n_293),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_480),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_547),
.B(n_428),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_480),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_568),
.B(n_293),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_469),
.B(n_189),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_547),
.B(n_192),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_563),
.B(n_428),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_556),
.Y(n_735)
);

AND2x6_ASAP7_75t_SL g736 ( 
.A(n_465),
.B(n_271),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_599),
.A2(n_425),
.B1(n_258),
.B2(n_195),
.C(n_200),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_484),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_563),
.B(n_428),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_567),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_567),
.B(n_428),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_522),
.A2(n_293),
.B1(n_427),
.B2(n_422),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_569),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_569),
.B(n_203),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_575),
.B(n_220),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_575),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_579),
.B(n_428),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_579),
.B(n_222),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_585),
.B(n_224),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_598),
.B(n_420),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_588),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_578),
.B(n_552),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_476),
.B(n_588),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_504),
.A2(n_395),
.B(n_403),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_495),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_484),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_594),
.B(n_428),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_594),
.B(n_512),
.Y(n_759)
);

BUFx12f_ASAP7_75t_SL g760 ( 
.A(n_476),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_492),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_549),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_475),
.B(n_393),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_458),
.B(n_566),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_595),
.B(n_158),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_458),
.B(n_428),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_592),
.A2(n_601),
.B1(n_600),
.B2(n_512),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_513),
.B(n_233),
.Y(n_768)
);

AND2x4_ASAP7_75t_SL g769 ( 
.A(n_513),
.B(n_271),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_514),
.B(n_428),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_514),
.B(n_427),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_634),
.B(n_516),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_635),
.A2(n_587),
.B(n_504),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_605),
.B(n_595),
.Y(n_774)
);

AO21x1_ASAP7_75t_L g775 ( 
.A1(n_653),
.A2(n_549),
.B(n_562),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_665),
.A2(n_499),
.B1(n_530),
.B2(n_543),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_645),
.B(n_516),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_616),
.B(n_533),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_645),
.B(n_642),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_642),
.B(n_533),
.Y(n_780)
);

BUFx8_ASAP7_75t_L g781 ( 
.A(n_751),
.Y(n_781)
);

OR2x2_ASAP7_75t_SL g782 ( 
.A(n_765),
.B(n_470),
.Y(n_782)
);

AOI21x1_ASAP7_75t_L g783 ( 
.A1(n_637),
.A2(n_601),
.B(n_600),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_627),
.B(n_180),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_639),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_605),
.B(n_534),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_679),
.B(n_534),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_698),
.A2(n_504),
.B(n_587),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_677),
.B(n_180),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_639),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_641),
.B(n_231),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_631),
.B(n_587),
.Y(n_792)
);

NOR2x2_ASAP7_75t_L g793 ( 
.A(n_703),
.B(n_536),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_611),
.A2(n_562),
.B(n_572),
.Y(n_794)
);

AOI21xp33_ASAP7_75t_L g795 ( 
.A1(n_641),
.A2(n_241),
.B(n_242),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_632),
.A2(n_553),
.B1(n_591),
.B2(n_590),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_658),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_658),
.Y(n_798)
);

AOI33xp33_ASAP7_75t_L g799 ( 
.A1(n_735),
.A2(n_273),
.A3(n_272),
.B1(n_279),
.B2(n_288),
.B3(n_290),
.Y(n_799)
);

AOI21x1_ASAP7_75t_L g800 ( 
.A1(n_633),
.A2(n_551),
.B(n_591),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_615),
.A2(n_572),
.B(n_482),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_604),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_660),
.A2(n_523),
.B(n_475),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_700),
.A2(n_632),
.B1(n_636),
.B2(n_676),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_636),
.B(n_536),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_604),
.B(n_542),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_656),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_661),
.A2(n_475),
.B(n_482),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_664),
.B(n_542),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_622),
.A2(n_482),
.B(n_523),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_608),
.A2(n_523),
.B(n_531),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_610),
.A2(n_531),
.B(n_565),
.Y(n_812)
);

BUFx4f_ASAP7_75t_L g813 ( 
.A(n_659),
.Y(n_813)
);

OAI21xp33_ASAP7_75t_L g814 ( 
.A1(n_704),
.A2(n_231),
.B(n_272),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_706),
.A2(n_531),
.B(n_565),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_663),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_755),
.A2(n_565),
.B(n_495),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_607),
.A2(n_558),
.B(n_590),
.C(n_589),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_626),
.A2(n_551),
.B(n_589),
.C(n_577),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_697),
.A2(n_597),
.B(n_495),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_664),
.B(n_546),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_626),
.B(n_546),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_720),
.A2(n_553),
.B(n_577),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_692),
.A2(n_597),
.B(n_495),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_650),
.B(n_557),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_680),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_612),
.B(n_557),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_693),
.A2(n_597),
.B(n_495),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_651),
.B(n_558),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_696),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_613),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_609),
.A2(n_571),
.B(n_500),
.C(n_493),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_694),
.A2(n_597),
.B(n_554),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_616),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_631),
.B(n_571),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_702),
.A2(n_597),
.B(n_554),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_621),
.B(n_246),
.Y(n_837)
);

NOR2x2_ASAP7_75t_L g838 ( 
.A(n_717),
.B(n_273),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_628),
.B(n_279),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_631),
.B(n_554),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_SL g841 ( 
.A1(n_764),
.A2(n_500),
.B(n_496),
.C(n_493),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_618),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_672),
.Y(n_843)
);

CKINVDCx8_ASAP7_75t_R g844 ( 
.A(n_736),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_631),
.B(n_499),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_631),
.B(n_499),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_756),
.A2(n_554),
.B(n_559),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_705),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_769),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_620),
.A2(n_499),
.B1(n_570),
.B2(n_543),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_631),
.B(n_616),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_672),
.Y(n_852)
);

AND2x2_ASAP7_75t_SL g853 ( 
.A(n_700),
.B(n_554),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_756),
.A2(n_559),
.B(n_492),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_616),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_720),
.A2(n_496),
.B(n_403),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_633),
.A2(n_559),
.B(n_395),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_710),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_740),
.B(n_499),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_629),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_743),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_762),
.A2(n_499),
.B(n_543),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_746),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_752),
.B(n_499),
.Y(n_864)
);

O2A1O1Ixp5_ASAP7_75t_L g865 ( 
.A1(n_625),
.A2(n_422),
.B(n_420),
.C(n_427),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_666),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_SL g867 ( 
.A(n_760),
.B(n_294),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_768),
.B(n_570),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_668),
.A2(n_559),
.B(n_402),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_SL g870 ( 
.A1(n_630),
.A2(n_395),
.B(n_396),
.C(n_402),
.Y(n_870)
);

INVx11_ASAP7_75t_L g871 ( 
.A(n_602),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_652),
.A2(n_420),
.B(n_422),
.C(n_427),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_629),
.B(n_559),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_701),
.B(n_420),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_669),
.A2(n_559),
.B(n_403),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_629),
.Y(n_876)
);

NAND2x1_ASAP7_75t_L g877 ( 
.A(n_629),
.B(n_570),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_617),
.B(n_247),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_603),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_684),
.A2(n_403),
.B(n_395),
.Y(n_880)
);

OAI21xp33_ASAP7_75t_L g881 ( 
.A1(n_704),
.A2(n_290),
.B(n_294),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_768),
.B(n_570),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_754),
.B(n_291),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_733),
.B(n_570),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_667),
.A2(n_252),
.B(n_253),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_681),
.B(n_667),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_619),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_753),
.A2(n_570),
.B1(n_543),
.B2(n_530),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_603),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_657),
.B(n_393),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_701),
.B(n_422),
.Y(n_891)
);

AOI33xp33_ASAP7_75t_L g892 ( 
.A1(n_644),
.A2(n_721),
.A3(n_707),
.B1(n_614),
.B2(n_727),
.B3(n_682),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_689),
.B(n_393),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_638),
.A2(n_396),
.B(n_402),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_648),
.A2(n_396),
.B(n_402),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_713),
.B(n_654),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_606),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_L g898 ( 
.A(n_603),
.B(n_543),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_762),
.A2(n_543),
.B(n_530),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_723),
.B(n_262),
.C(n_265),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_602),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_624),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_759),
.A2(n_267),
.B1(n_288),
.B2(n_291),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_646),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_673),
.A2(n_570),
.B1(n_543),
.B2(n_530),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_733),
.B(n_530),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_673),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_767),
.A2(n_530),
.B(n_396),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_713),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_712),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_644),
.B(n_393),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_759),
.A2(n_393),
.B(n_530),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_744),
.Y(n_913)
);

INVx8_ASAP7_75t_L g914 ( 
.A(n_673),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_673),
.B(n_393),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_647),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_744),
.B(n_393),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_655),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_681),
.B(n_11),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_649),
.A2(n_12),
.B(n_15),
.C(n_16),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_745),
.B(n_393),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_695),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_716),
.A2(n_393),
.B1(n_151),
.B2(n_145),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_670),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_673),
.A2(n_12),
.B1(n_16),
.B2(n_19),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_745),
.B(n_19),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_748),
.B(n_20),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_623),
.B(n_21),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_678),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_687),
.B(n_22),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_675),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_716),
.A2(n_136),
.B1(n_132),
.B2(n_119),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_766),
.A2(n_116),
.B(n_114),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_630),
.A2(n_113),
.B(n_108),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_742),
.B(n_102),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_725),
.B(n_98),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_671),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_726),
.A2(n_97),
.B(n_77),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_686),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_723),
.B(n_22),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_748),
.B(n_26),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_732),
.B(n_26),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_699),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_729),
.A2(n_73),
.B(n_29),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_732),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_734),
.A2(n_27),
.B(n_35),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_709),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_739),
.A2(n_36),
.B(n_38),
.Y(n_948)
);

AO21x1_ASAP7_75t_L g949 ( 
.A1(n_687),
.A2(n_36),
.B(n_38),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_741),
.A2(n_39),
.B(n_42),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_749),
.B(n_39),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_747),
.A2(n_42),
.B(n_44),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_758),
.A2(n_45),
.B(n_49),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_749),
.B(n_52),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_771),
.A2(n_52),
.B(n_770),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_688),
.A2(n_731),
.B(n_719),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_691),
.B(n_730),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_643),
.B(n_691),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_711),
.A2(n_761),
.B(n_757),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_714),
.B(n_738),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_807),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_886),
.A2(n_722),
.B1(n_690),
.B2(n_662),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_913),
.B(n_685),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_913),
.B(n_685),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_779),
.B(n_958),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_852),
.B(n_843),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_909),
.Y(n_967)
);

AOI21xp33_ASAP7_75t_L g968 ( 
.A1(n_958),
.A2(n_715),
.B(n_737),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_792),
.A2(n_640),
.B(n_674),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_940),
.A2(n_683),
.B1(n_708),
.B2(n_750),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_791),
.A2(n_718),
.B(n_724),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_786),
.B(n_728),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_827),
.Y(n_973)
);

AOI222xp33_ASAP7_75t_L g974 ( 
.A1(n_940),
.A2(n_750),
.B1(n_763),
.B2(n_942),
.C1(n_881),
.C2(n_814),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_774),
.B(n_750),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_909),
.B(n_763),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_774),
.B(n_763),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_792),
.A2(n_763),
.B(n_835),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_800),
.A2(n_763),
.B(n_783),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_788),
.A2(n_773),
.B(n_845),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_789),
.B(n_839),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_786),
.B(n_809),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_879),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_809),
.B(n_821),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_831),
.B(n_896),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_879),
.B(n_867),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_831),
.B(n_896),
.Y(n_987)
);

NAND3xp33_ASAP7_75t_SL g988 ( 
.A(n_900),
.B(n_942),
.C(n_927),
.Y(n_988)
);

INVx3_ASAP7_75t_SL g989 ( 
.A(n_793),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_926),
.A2(n_954),
.B(n_941),
.C(n_951),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_879),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_781),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_816),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_821),
.B(n_780),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_879),
.Y(n_995)
);

CKINVDCx14_ASAP7_75t_R g996 ( 
.A(n_937),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_871),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_919),
.A2(n_930),
.B(n_928),
.C(n_878),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_827),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_858),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_846),
.A2(n_840),
.B(n_851),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_840),
.A2(n_851),
.B(n_829),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_826),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_822),
.B(n_866),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_SL g1005 ( 
.A1(n_897),
.A2(n_782),
.B1(n_844),
.B2(n_925),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_917),
.A2(n_921),
.B(n_805),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_795),
.A2(n_885),
.B(n_928),
.C(n_952),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_830),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_878),
.A2(n_837),
.B(n_799),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_822),
.B(n_804),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_892),
.A2(n_900),
.B(n_837),
.C(n_777),
.Y(n_1011)
);

INVx6_ASAP7_75t_L g1012 ( 
.A(n_781),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_848),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_922),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_804),
.A2(n_853),
.B1(n_825),
.B2(n_787),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_817),
.A2(n_824),
.B(n_833),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_861),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_842),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_931),
.B(n_785),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_790),
.B(n_784),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_834),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_863),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_813),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_920),
.A2(n_935),
.B(n_957),
.C(n_949),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_842),
.Y(n_1025)
);

AOI222xp33_ASAP7_75t_L g1026 ( 
.A1(n_925),
.A2(n_903),
.B1(n_883),
.B2(n_935),
.C1(n_901),
.C2(n_853),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_874),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_806),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_874),
.B(n_891),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_884),
.A2(n_906),
.B(n_938),
.C(n_868),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_882),
.A2(n_818),
.B(n_772),
.C(n_797),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_910),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_798),
.B(n_891),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_834),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_806),
.B(n_802),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_828),
.A2(n_836),
.B(n_820),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_916),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_849),
.B(n_802),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_856),
.A2(n_810),
.B(n_812),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_910),
.B(n_813),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_794),
.A2(n_893),
.B(n_801),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_943),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_893),
.A2(n_898),
.B(n_915),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_901),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_945),
.A2(n_923),
.B1(n_932),
.B2(n_946),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_947),
.B(n_939),
.Y(n_1046)
);

OA21x2_ASAP7_75t_L g1047 ( 
.A1(n_865),
.A2(n_819),
.B(n_823),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_947),
.B(n_924),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_887),
.B(n_929),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_890),
.A2(n_815),
.B(n_808),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_834),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_902),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_911),
.A2(n_862),
.B(n_899),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_834),
.B(n_876),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_904),
.B(n_918),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_888),
.A2(n_876),
.B1(n_860),
.B2(n_855),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_960),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_911),
.B(n_956),
.Y(n_1058)
);

O2A1O1Ixp5_ASAP7_75t_L g1059 ( 
.A1(n_775),
.A2(n_936),
.B(n_890),
.C(n_955),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_803),
.A2(n_811),
.B(n_873),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_873),
.A2(n_847),
.B(n_908),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_855),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_956),
.B(n_953),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_778),
.Y(n_1064)
);

BUFx12f_ASAP7_75t_L g1065 ( 
.A(n_855),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_796),
.B(n_876),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_959),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_865),
.A2(n_869),
.B(n_875),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_950),
.B(n_944),
.C(n_936),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_948),
.B(n_855),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_854),
.A2(n_859),
.B(n_864),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_860),
.B(n_876),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_776),
.A2(n_850),
.B1(n_860),
.B2(n_907),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_860),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_914),
.A2(n_912),
.B(n_841),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_914),
.A2(n_841),
.B(n_778),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_888),
.A2(n_907),
.B1(n_914),
.B2(n_889),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_907),
.A2(n_934),
.B1(n_933),
.B2(n_905),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_877),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_889),
.B(n_907),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_832),
.A2(n_872),
.B(n_870),
.C(n_895),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_905),
.B(n_857),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_894),
.B(n_880),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_838),
.B(n_779),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_L g1085 ( 
.A(n_958),
.B(n_886),
.C(n_641),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_779),
.B(n_886),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_886),
.B(n_913),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_779),
.B(n_886),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_909),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_779),
.B(n_886),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_909),
.B(n_874),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_958),
.A2(n_641),
.B(n_886),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_800),
.A2(n_783),
.B(n_856),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_871),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_958),
.A2(n_942),
.B(n_940),
.C(n_927),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_879),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_827),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_958),
.A2(n_940),
.B(n_942),
.C(n_490),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_958),
.A2(n_886),
.B1(n_804),
.B2(n_913),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_827),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_779),
.B(n_886),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_886),
.B(n_913),
.Y(n_1102)
);

INVx4_ASAP7_75t_L g1103 ( 
.A(n_879),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_958),
.A2(n_886),
.B1(n_804),
.B2(n_913),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_779),
.B(n_913),
.Y(n_1105)
);

CKINVDCx8_ASAP7_75t_R g1106 ( 
.A(n_852),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_791),
.B(n_677),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_R g1108 ( 
.A(n_879),
.B(n_470),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1095),
.A2(n_1007),
.B(n_998),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1006),
.A2(n_1030),
.B(n_969),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_961),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_1014),
.Y(n_1112)
);

AO22x2_ASAP7_75t_L g1113 ( 
.A1(n_1099),
.A2(n_1104),
.B1(n_988),
.B2(n_1085),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1092),
.A2(n_965),
.B(n_968),
.C(n_990),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1043),
.A2(n_984),
.B(n_980),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1032),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1098),
.A2(n_988),
.B(n_965),
.C(n_1011),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_979),
.A2(n_1093),
.B(n_1075),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1041),
.A2(n_1036),
.B(n_982),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1009),
.A2(n_1024),
.B(n_962),
.C(n_971),
.Y(n_1120)
);

AOI211x1_ASAP7_75t_L g1121 ( 
.A1(n_1087),
.A2(n_1102),
.B(n_1101),
.C(n_1090),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1010),
.A2(n_975),
.B(n_1045),
.C(n_970),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1039),
.A2(n_1076),
.B(n_1060),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_997),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_993),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_963),
.A2(n_964),
.B(n_1088),
.C(n_1086),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1000),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_1025),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_1045),
.B(n_1026),
.C(n_974),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1016),
.A2(n_1071),
.B(n_1068),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1059),
.A2(n_1015),
.B(n_1053),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_975),
.A2(n_1105),
.B(n_985),
.C(n_987),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_1050),
.A2(n_1083),
.A3(n_1058),
.B(n_1061),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1001),
.A2(n_978),
.B(n_1002),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1083),
.A2(n_1031),
.A3(n_1067),
.B(n_1056),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1081),
.A2(n_1059),
.B(n_1066),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1105),
.B(n_994),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1107),
.B(n_981),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1020),
.B(n_1084),
.C(n_987),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1084),
.A2(n_1020),
.B1(n_985),
.B2(n_1005),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_1012),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1037),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1063),
.A2(n_1082),
.B(n_1069),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1044),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1003),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1025),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1077),
.A2(n_1078),
.B(n_1047),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_986),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1078),
.A2(n_1047),
.B(n_1070),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1073),
.A2(n_1079),
.B(n_1064),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1091),
.B(n_1027),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1089),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1069),
.A2(n_1004),
.B(n_977),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_972),
.A2(n_977),
.B1(n_1042),
.B2(n_1057),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1080),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1072),
.A2(n_1054),
.B(n_1049),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1046),
.A2(n_1048),
.B(n_1035),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_989),
.B(n_967),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1065),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1089),
.B(n_1091),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_967),
.A2(n_989),
.B(n_1042),
.C(n_1018),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1012),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1013),
.A2(n_1017),
.A3(n_1022),
.B(n_1033),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1019),
.B(n_1018),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1074),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1034),
.A2(n_1052),
.B(n_1008),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_1012),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1034),
.A2(n_973),
.B(n_1097),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1029),
.A2(n_1033),
.B(n_1080),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1019),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_976),
.A2(n_999),
.B(n_1100),
.Y(n_1171)
);

OAI22x1_ASAP7_75t_L g1172 ( 
.A1(n_1023),
.A2(n_1038),
.B1(n_1027),
.B2(n_1040),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1028),
.A2(n_1038),
.B1(n_966),
.B2(n_1051),
.Y(n_1173)
);

NAND2xp33_ASAP7_75t_L g1174 ( 
.A(n_986),
.B(n_1108),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1106),
.B(n_996),
.Y(n_1175)
);

CKINVDCx11_ASAP7_75t_R g1176 ( 
.A(n_966),
.Y(n_1176)
);

AOI221x1_ASAP7_75t_L g1177 ( 
.A1(n_1021),
.A2(n_983),
.B1(n_991),
.B2(n_1103),
.C(n_995),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1108),
.B(n_1062),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1021),
.B(n_995),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_983),
.A2(n_991),
.B1(n_1096),
.B2(n_1103),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_983),
.B(n_966),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1094),
.A2(n_992),
.B(n_1006),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_979),
.A2(n_1093),
.B(n_1075),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_965),
.B(n_1086),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_997),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1095),
.A2(n_958),
.B(n_1007),
.C(n_1092),
.Y(n_1189)
);

BUFx10_ASAP7_75t_L g1190 ( 
.A(n_1012),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_965),
.B(n_779),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1080),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1193)
);

AO22x2_ASAP7_75t_L g1194 ( 
.A1(n_1099),
.A2(n_1104),
.B1(n_988),
.B2(n_1085),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_L g1195 ( 
.A(n_988),
.B(n_913),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1107),
.B(n_677),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1030),
.A2(n_775),
.A3(n_1015),
.B(n_980),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_961),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1080),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1032),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_965),
.B(n_1086),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_965),
.B(n_984),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1032),
.Y(n_1204)
);

NAND2x1_ASAP7_75t_L g1205 ( 
.A(n_1021),
.B(n_834),
.Y(n_1205)
);

OAI211xp5_ASAP7_75t_L g1206 ( 
.A1(n_1095),
.A2(n_958),
.B(n_814),
.C(n_881),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1207)
);

INVx5_ASAP7_75t_L g1208 ( 
.A(n_1065),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1065),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1030),
.A2(n_775),
.A3(n_1015),
.B(n_980),
.Y(n_1211)
);

AOI21xp33_ASAP7_75t_L g1212 ( 
.A1(n_1095),
.A2(n_1007),
.B(n_1098),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_961),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_965),
.A2(n_1085),
.B1(n_984),
.B2(n_958),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1107),
.B(n_677),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1065),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_988),
.A2(n_980),
.B(n_1030),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1059),
.A2(n_1030),
.B(n_980),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_965),
.B(n_1086),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_965),
.B(n_1086),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_961),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_961),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1086),
.B(n_735),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1030),
.A2(n_775),
.A3(n_1015),
.B(n_980),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_979),
.A2(n_1093),
.B(n_1075),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_979),
.A2(n_1093),
.B(n_1075),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1030),
.A2(n_775),
.A3(n_1015),
.B(n_980),
.Y(n_1229)
);

AOI221xp5_ASAP7_75t_SL g1230 ( 
.A1(n_1095),
.A2(n_1007),
.B1(n_1104),
.B2(n_1099),
.C(n_1092),
.Y(n_1230)
);

BUFx10_ASAP7_75t_L g1231 ( 
.A(n_1012),
.Y(n_1231)
);

AOI221x1_ASAP7_75t_L g1232 ( 
.A1(n_988),
.A2(n_1092),
.B1(n_998),
.B2(n_942),
.C(n_940),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1092),
.A2(n_958),
.B1(n_886),
.B2(n_942),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1095),
.A2(n_1007),
.B(n_998),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_961),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1095),
.A2(n_958),
.B(n_1007),
.C(n_1092),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_965),
.B(n_1086),
.Y(n_1239)
);

OAI22x1_ASAP7_75t_L g1240 ( 
.A1(n_965),
.A2(n_958),
.B1(n_940),
.B2(n_942),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_965),
.B(n_779),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_L g1242 ( 
.A(n_997),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1030),
.A2(n_775),
.A3(n_1015),
.B(n_980),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_979),
.A2(n_1093),
.B(n_1075),
.Y(n_1244)
);

BUFx4_ASAP7_75t_SL g1245 ( 
.A(n_997),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1025),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1006),
.A2(n_568),
.B(n_1030),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1030),
.A2(n_775),
.A3(n_1015),
.B(n_980),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_979),
.A2(n_1093),
.B(n_1075),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_965),
.B(n_1086),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1032),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1129),
.A2(n_1241),
.B1(n_1191),
.B2(n_1233),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1111),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1125),
.Y(n_1254)
);

CKINVDCx6p67_ASAP7_75t_R g1255 ( 
.A(n_1208),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1245),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1187),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1129),
.A2(n_1233),
.B1(n_1203),
.B2(n_1250),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1240),
.A2(n_1109),
.B1(n_1235),
.B2(n_1214),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1206),
.A2(n_1109),
.B1(n_1235),
.B2(n_1113),
.Y(n_1260)
);

BUFx4_ASAP7_75t_R g1261 ( 
.A(n_1141),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1203),
.A2(n_1221),
.B1(n_1201),
.B2(n_1185),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1124),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1242),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1113),
.A2(n_1194),
.B1(n_1214),
.B2(n_1139),
.Y(n_1265)
);

BUFx4_ASAP7_75t_SL g1266 ( 
.A(n_1148),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1194),
.A2(n_1195),
.B1(n_1139),
.B2(n_1212),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1220),
.B(n_1239),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1195),
.A2(n_1212),
.B1(n_1140),
.B2(n_1216),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1127),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1141),
.Y(n_1271)
);

BUFx8_ASAP7_75t_L g1272 ( 
.A(n_1159),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1140),
.A2(n_1232),
.B(n_1189),
.Y(n_1273)
);

INVx6_ASAP7_75t_L g1274 ( 
.A(n_1167),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1196),
.A2(n_1138),
.B1(n_1170),
.B2(n_1172),
.Y(n_1275)
);

CKINVDCx14_ASAP7_75t_R g1276 ( 
.A(n_1176),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1167),
.Y(n_1277)
);

CKINVDCx11_ASAP7_75t_R g1278 ( 
.A(n_1190),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1155),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1190),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1137),
.B(n_1132),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1114),
.B(n_1238),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1213),
.Y(n_1283)
);

INVx3_ASAP7_75t_SL g1284 ( 
.A(n_1231),
.Y(n_1284)
);

CKINVDCx6p67_ASAP7_75t_R g1285 ( 
.A(n_1208),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1120),
.A2(n_1117),
.B(n_1122),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1170),
.A2(n_1224),
.B1(n_1153),
.B2(n_1151),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1222),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1153),
.A2(n_1151),
.B1(n_1174),
.B2(n_1218),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1218),
.A2(n_1131),
.B1(n_1154),
.B2(n_1158),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1131),
.A2(n_1164),
.B1(n_1143),
.B2(n_1128),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1223),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1165),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1143),
.A2(n_1230),
.B1(n_1154),
.B2(n_1246),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1236),
.Y(n_1295)
);

BUFx5_ASAP7_75t_L g1296 ( 
.A(n_1142),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1145),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1169),
.A2(n_1171),
.B1(n_1160),
.B2(n_1173),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1112),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1121),
.A2(n_1173),
.B1(n_1126),
.B2(n_1146),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1231),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1163),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1178),
.A2(n_1182),
.B1(n_1144),
.B2(n_1162),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1159),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1152),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1209),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1181),
.A2(n_1116),
.B1(n_1171),
.B2(n_1209),
.Y(n_1307)
);

BUFx10_ASAP7_75t_L g1308 ( 
.A(n_1175),
.Y(n_1308)
);

BUFx4_ASAP7_75t_R g1309 ( 
.A(n_1251),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1181),
.A2(n_1209),
.B1(n_1217),
.B2(n_1199),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1217),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1166),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_1200),
.Y(n_1313)
);

BUFx4f_ASAP7_75t_SL g1314 ( 
.A(n_1204),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1150),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1230),
.B(n_1135),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1155),
.A2(n_1192),
.B1(n_1199),
.B2(n_1110),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1161),
.A2(n_1210),
.B(n_1247),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1192),
.A2(n_1115),
.B1(n_1219),
.B2(n_1188),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1135),
.B(n_1136),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1156),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1179),
.B(n_1180),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1219),
.A2(n_1157),
.B1(n_1193),
.B2(n_1237),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1180),
.A2(n_1227),
.B1(n_1202),
.B2(n_1215),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1183),
.A2(n_1234),
.B1(n_1207),
.B2(n_1186),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1168),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1147),
.A2(n_1149),
.B1(n_1119),
.B2(n_1134),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1135),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1205),
.A2(n_1177),
.B1(n_1248),
.B2(n_1243),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1133),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1133),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1130),
.A2(n_1118),
.B1(n_1249),
.B2(n_1244),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1197),
.A2(n_1248),
.B1(n_1243),
.B2(n_1211),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1184),
.A2(n_1226),
.B1(n_1228),
.B2(n_1123),
.Y(n_1334)
);

BUFx2_ASAP7_75t_SL g1335 ( 
.A(n_1133),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1197),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1197),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1248),
.Y(n_1338)
);

INVx6_ASAP7_75t_L g1339 ( 
.A(n_1211),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1225),
.A2(n_1129),
.B1(n_1140),
.B2(n_1233),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1229),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1229),
.A2(n_1129),
.B1(n_958),
.B2(n_886),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1243),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1198),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1129),
.A2(n_958),
.B1(n_886),
.B2(n_988),
.Y(n_1345)
);

INVx6_ASAP7_75t_L g1346 ( 
.A(n_1141),
.Y(n_1346)
);

INVx6_ASAP7_75t_L g1347 ( 
.A(n_1141),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1203),
.B(n_965),
.Y(n_1348)
);

CKINVDCx6p67_ASAP7_75t_R g1349 ( 
.A(n_1208),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1198),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1129),
.A2(n_958),
.B1(n_886),
.B2(n_988),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1198),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1198),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1198),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1129),
.A2(n_958),
.B1(n_886),
.B2(n_988),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1155),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1160),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1129),
.A2(n_958),
.B1(n_886),
.B2(n_988),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1198),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1198),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1198),
.Y(n_1361)
);

BUFx2_ASAP7_75t_SL g1362 ( 
.A(n_1124),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1198),
.Y(n_1363)
);

BUFx4f_ASAP7_75t_L g1364 ( 
.A(n_1159),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1198),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1245),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1129),
.A2(n_958),
.B1(n_886),
.B2(n_988),
.Y(n_1367)
);

BUFx4f_ASAP7_75t_SL g1368 ( 
.A(n_1242),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1160),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1203),
.B(n_965),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1203),
.B(n_965),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1268),
.B(n_1262),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1319),
.A2(n_1323),
.B(n_1334),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1265),
.B(n_1259),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1319),
.A2(n_1332),
.B(n_1325),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1330),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1268),
.B(n_1262),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_SL g1378 ( 
.A(n_1318),
.B(n_1329),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1302),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1271),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1299),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1305),
.Y(n_1382)
);

AO22x1_ASAP7_75t_L g1383 ( 
.A1(n_1252),
.A2(n_1282),
.B1(n_1281),
.B2(n_1258),
.Y(n_1383)
);

BUFx8_ASAP7_75t_L g1384 ( 
.A(n_1304),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1357),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1328),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1337),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1336),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1339),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_SL g1390 ( 
.A(n_1286),
.B(n_1273),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1271),
.Y(n_1391)
);

OAI222xp33_ASAP7_75t_L g1392 ( 
.A1(n_1252),
.A2(n_1260),
.B1(n_1358),
.B2(n_1345),
.C1(n_1367),
.C2(n_1351),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1264),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1338),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1324),
.A2(n_1333),
.B(n_1329),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1342),
.B(n_1290),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1296),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1357),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1341),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1256),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1315),
.A2(n_1321),
.B(n_1312),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1343),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1296),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1316),
.B(n_1320),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1296),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1355),
.A2(n_1258),
.B1(n_1269),
.B2(n_1303),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1320),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1282),
.A2(n_1281),
.B1(n_1336),
.B2(n_1300),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1369),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1348),
.A2(n_1371),
.B1(n_1370),
.B2(n_1275),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1340),
.A2(n_1287),
.B1(n_1289),
.B2(n_1291),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1322),
.A2(n_1300),
.B(n_1326),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1331),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1335),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1291),
.A2(n_1298),
.B1(n_1267),
.B2(n_1294),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1253),
.A2(n_1270),
.B(n_1254),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1283),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1288),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1266),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_SL g1420 ( 
.A(n_1366),
.B(n_1257),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1292),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1369),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1279),
.B(n_1356),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1295),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1293),
.B(n_1371),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1297),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1271),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1370),
.B(n_1348),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1344),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1350),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1352),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1294),
.B(n_1359),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1353),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1317),
.A2(n_1360),
.B(n_1354),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1274),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1363),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1307),
.A2(n_1310),
.B(n_1327),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1361),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1365),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1274),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1327),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1276),
.A2(n_1308),
.B1(n_1356),
.B2(n_1279),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1274),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1346),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_SL g1445 ( 
.A1(n_1261),
.A2(n_1255),
.B(n_1349),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1346),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1346),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1285),
.A2(n_1347),
.B(n_1311),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1347),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1347),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1311),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1311),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1368),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1278),
.Y(n_1454)
);

NOR2x1_ASAP7_75t_R g1455 ( 
.A(n_1277),
.B(n_1301),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1280),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1373),
.A2(n_1308),
.B(n_1309),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1385),
.B(n_1263),
.Y(n_1458)
);

AOI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1390),
.A2(n_1284),
.B1(n_1364),
.B2(n_1362),
.C(n_1313),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1390),
.A2(n_1272),
.B(n_1306),
.C(n_1313),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1389),
.B(n_1272),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1398),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1409),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1393),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1392),
.A2(n_1314),
.B1(n_1383),
.B2(n_1374),
.C(n_1415),
.Y(n_1465)
);

OR2x6_ASAP7_75t_L g1466 ( 
.A(n_1375),
.B(n_1373),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1384),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1400),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1422),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1416),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1417),
.B(n_1421),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1425),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1428),
.B(n_1372),
.Y(n_1473)
);

OAI211xp5_ASAP7_75t_L g1474 ( 
.A1(n_1406),
.A2(n_1411),
.B(n_1408),
.C(n_1374),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1377),
.B(n_1383),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_SL g1476 ( 
.A1(n_1380),
.A2(n_1435),
.B(n_1427),
.C(n_1391),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1421),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1396),
.B(n_1432),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1396),
.B(n_1432),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1410),
.A2(n_1388),
.B(n_1441),
.C(n_1375),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1378),
.A2(n_1395),
.B(n_1437),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1442),
.A2(n_1412),
.B(n_1381),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1420),
.B(n_1419),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1388),
.B(n_1448),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1416),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1412),
.A2(n_1382),
.B(n_1448),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1418),
.B(n_1424),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1426),
.Y(n_1488)
);

NAND4xp25_ASAP7_75t_L g1489 ( 
.A(n_1429),
.B(n_1431),
.C(n_1433),
.D(n_1426),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1388),
.A2(n_1378),
.B(n_1395),
.C(n_1437),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1456),
.B(n_1444),
.Y(n_1491)
);

BUFx2_ASAP7_75t_R g1492 ( 
.A(n_1437),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1395),
.B(n_1407),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1445),
.A2(n_1449),
.B(n_1447),
.C(n_1446),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1376),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1407),
.B(n_1404),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1401),
.A2(n_1414),
.B(n_1402),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_SL g1498 ( 
.A1(n_1427),
.A2(n_1443),
.B(n_1440),
.C(n_1435),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1430),
.B(n_1436),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1454),
.A2(n_1453),
.B1(n_1449),
.B2(n_1440),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1445),
.A2(n_1446),
.B(n_1450),
.C(n_1447),
.Y(n_1501)
);

AO21x1_ASAP7_75t_L g1502 ( 
.A1(n_1413),
.A2(n_1439),
.B(n_1438),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1493),
.B(n_1376),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1497),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1466),
.B(n_1397),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1465),
.A2(n_1454),
.B1(n_1434),
.B2(n_1384),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1475),
.B(n_1450),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1466),
.B(n_1495),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1474),
.A2(n_1434),
.B1(n_1423),
.B2(n_1446),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1484),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1466),
.B(n_1405),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1470),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1497),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1496),
.B(n_1379),
.Y(n_1514)
);

NOR2x1_ASAP7_75t_L g1515 ( 
.A(n_1490),
.B(n_1403),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1485),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1484),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1481),
.B(n_1386),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1484),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1477),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1484),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1471),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1473),
.B(n_1387),
.Y(n_1523)
);

INVxp67_ASAP7_75t_SL g1524 ( 
.A(n_1502),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1510),
.Y(n_1525)
);

AOI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1515),
.A2(n_1457),
.B(n_1486),
.Y(n_1526)
);

NAND4xp25_ASAP7_75t_SL g1527 ( 
.A(n_1506),
.B(n_1490),
.C(n_1459),
.D(n_1480),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1522),
.B(n_1457),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1512),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1513),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1522),
.B(n_1457),
.Y(n_1531)
);

OAI33xp33_ASAP7_75t_L g1532 ( 
.A1(n_1523),
.A2(n_1489),
.A3(n_1472),
.B1(n_1500),
.B2(n_1488),
.B3(n_1458),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1516),
.B(n_1462),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1513),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1512),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1516),
.B(n_1463),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1520),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1505),
.B(n_1499),
.Y(n_1538)
);

OAI33xp33_ASAP7_75t_L g1539 ( 
.A1(n_1523),
.A2(n_1494),
.A3(n_1501),
.B1(n_1387),
.B2(n_1394),
.B3(n_1399),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1520),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1522),
.B(n_1487),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1512),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1508),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1523),
.B(n_1469),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1524),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1487),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1504),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_L g1548 ( 
.A(n_1524),
.B(n_1480),
.C(n_1482),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1516),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1514),
.B(n_1507),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1506),
.A2(n_1492),
.B1(n_1479),
.B2(n_1478),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1514),
.B(n_1477),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1545),
.B(n_1507),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1533),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1545),
.B(n_1503),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1543),
.B(n_1517),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1547),
.B(n_1510),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1532),
.B(n_1548),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1548),
.B(n_1509),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1528),
.B(n_1517),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1517),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1529),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1537),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1529),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1528),
.B(n_1531),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1517),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1529),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1537),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1535),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1531),
.B(n_1508),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1508),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1535),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1538),
.B(n_1508),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1575)
);

INVxp67_ASAP7_75t_SL g1576 ( 
.A(n_1540),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1541),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1541),
.B(n_1511),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1532),
.B(n_1491),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1550),
.B(n_1503),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1550),
.B(n_1503),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1549),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1533),
.B(n_1518),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1535),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1533),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1544),
.B(n_1503),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1542),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1557),
.B(n_1510),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1536),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1588),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1553),
.B(n_1536),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1554),
.B(n_1536),
.Y(n_1593)
);

NAND2x1_ASAP7_75t_L g1594 ( 
.A(n_1557),
.B(n_1515),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1558),
.A2(n_1551),
.B1(n_1509),
.B2(n_1460),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_SL g1596 ( 
.A(n_1558),
.B(n_1467),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1580),
.B(n_1454),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1588),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1578),
.B(n_1525),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1562),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1578),
.B(n_1525),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1544),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1559),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1557),
.B(n_1467),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1583),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1567),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1563),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_1559),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1554),
.B(n_1552),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1581),
.B(n_1454),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1571),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1567),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1562),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1562),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1564),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1571),
.B(n_1525),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1586),
.B(n_1552),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1563),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.B(n_1525),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1581),
.B(n_1541),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1564),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1583),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1564),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1573),
.B(n_1510),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1573),
.B(n_1510),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1569),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1582),
.B(n_1546),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1582),
.B(n_1546),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1587),
.B(n_1546),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1587),
.B(n_1454),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1590),
.B(n_1586),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1596),
.Y(n_1632)
);

NAND2x1_ASAP7_75t_L g1633 ( 
.A(n_1589),
.B(n_1557),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1599),
.B(n_1573),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1603),
.B(n_1579),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1574),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1611),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1607),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1608),
.A2(n_1527),
.B1(n_1551),
.B2(n_1521),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1611),
.B(n_1557),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1600),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1590),
.B(n_1584),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1600),
.Y(n_1644)
);

NOR2x1p5_ASAP7_75t_SL g1645 ( 
.A(n_1605),
.B(n_1583),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1592),
.B(n_1584),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1601),
.B(n_1557),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1592),
.B(n_1584),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1616),
.B(n_1575),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1605),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1597),
.B(n_1579),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1575),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1602),
.B(n_1579),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1619),
.B(n_1575),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1613),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1610),
.B(n_1555),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1622),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1614),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1589),
.B(n_1577),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1589),
.B(n_1577),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1630),
.B(n_1595),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1614),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1624),
.B(n_1577),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1655),
.B(n_1609),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1642),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1650),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1642),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1644),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1632),
.B(n_1647),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1650),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1639),
.B(n_1618),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1663),
.B(n_1609),
.Y(n_1674)
);

OAI32xp33_ASAP7_75t_L g1675 ( 
.A1(n_1636),
.A2(n_1593),
.A3(n_1617),
.B1(n_1555),
.B2(n_1626),
.Y(n_1675)
);

O2A1O1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1631),
.A2(n_1460),
.B(n_1568),
.C(n_1576),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1644),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1654),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1640),
.A2(n_1594),
.B(n_1509),
.C(n_1604),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1652),
.B(n_1617),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1654),
.Y(n_1681)
);

OAI32xp33_ASAP7_75t_L g1682 ( 
.A1(n_1631),
.A2(n_1593),
.A3(n_1591),
.B1(n_1598),
.B2(n_1606),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1633),
.A2(n_1594),
.B1(n_1576),
.B2(n_1568),
.C(n_1612),
.Y(n_1683)
);

OAI21xp33_ASAP7_75t_SL g1684 ( 
.A1(n_1662),
.A2(n_1625),
.B(n_1624),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1657),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1650),
.B(n_1625),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1556),
.Y(n_1687)
);

A2O1A1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1645),
.A2(n_1483),
.B(n_1527),
.C(n_1515),
.Y(n_1688)
);

AO22x1_ASAP7_75t_L g1689 ( 
.A1(n_1647),
.A2(n_1454),
.B1(n_1384),
.B2(n_1468),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1647),
.A2(n_1519),
.B1(n_1521),
.B2(n_1539),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1688),
.B(n_1641),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1686),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1671),
.B(n_1638),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1667),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1688),
.A2(n_1638),
.B1(n_1526),
.B2(n_1633),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1674),
.B(n_1634),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1686),
.A2(n_1641),
.B1(n_1661),
.B2(n_1650),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1686),
.A2(n_1641),
.B1(n_1661),
.B2(n_1662),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1668),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1680),
.A2(n_1641),
.B1(n_1661),
.B2(n_1658),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1670),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1682),
.A2(n_1468),
.B(n_1455),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1673),
.B(n_1634),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1643),
.Y(n_1705)
);

AOI222xp33_ASAP7_75t_L g1706 ( 
.A1(n_1675),
.A2(n_1645),
.B1(n_1539),
.B2(n_1664),
.C1(n_1660),
.C2(n_1657),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1687),
.A2(n_1661),
.B1(n_1637),
.B2(n_1635),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1689),
.B(n_1464),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1668),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_L g1710 ( 
.A(n_1706),
.B(n_1676),
.C(n_1679),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1695),
.B(n_1679),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1708),
.A2(n_1676),
.B(n_1683),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1692),
.B(n_1672),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1692),
.B(n_1672),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1693),
.B(n_1677),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1691),
.B(n_1678),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1703),
.A2(n_1690),
.B(n_1684),
.C(n_1685),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1696),
.B(n_1705),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1704),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1700),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1710),
.A2(n_1701),
.B1(n_1697),
.B2(n_1698),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1719),
.B(n_1709),
.Y(n_1722)
);

AOI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1711),
.A2(n_1695),
.B(n_1702),
.C(n_1699),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1712),
.A2(n_1694),
.B1(n_1681),
.B2(n_1707),
.C(n_1706),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1716),
.B(n_1718),
.Y(n_1725)
);

AO21x1_ASAP7_75t_L g1726 ( 
.A1(n_1713),
.A2(n_1714),
.B(n_1720),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1715),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1717),
.B(n_1646),
.C(n_1643),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1719),
.B(n_1464),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1635),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1725),
.A2(n_1664),
.B(n_1660),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1722),
.B(n_1651),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1724),
.A2(n_1648),
.B1(n_1646),
.B2(n_1637),
.Y(n_1733)
);

AOI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1721),
.A2(n_1455),
.B(n_1648),
.C(n_1656),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1728),
.B(n_1651),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1723),
.A2(n_1656),
.B1(n_1653),
.B2(n_1649),
.Y(n_1736)
);

XOR2x2_ASAP7_75t_L g1737 ( 
.A(n_1734),
.B(n_1729),
.Y(n_1737)
);

AOI322xp5_ASAP7_75t_L g1738 ( 
.A1(n_1735),
.A2(n_1727),
.A3(n_1733),
.B1(n_1732),
.B2(n_1730),
.C1(n_1726),
.C2(n_1649),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1731),
.B(n_1653),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1736),
.A2(n_1659),
.B1(n_1665),
.B2(n_1615),
.C(n_1621),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1733),
.A2(n_1659),
.B1(n_1665),
.B2(n_1615),
.C(n_1621),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1733),
.A2(n_1623),
.B1(n_1622),
.B2(n_1627),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1733),
.A2(n_1623),
.B1(n_1556),
.B2(n_1561),
.C(n_1560),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1737),
.A2(n_1384),
.B1(n_1565),
.B2(n_1560),
.Y(n_1744)
);

NOR2x1_ASAP7_75t_L g1745 ( 
.A(n_1739),
.B(n_1583),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1741),
.A2(n_1565),
.B1(n_1560),
.B2(n_1561),
.C(n_1566),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1742),
.Y(n_1747)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1748 ( 
.A1(n_1738),
.A2(n_1585),
.B(n_1569),
.C(n_1572),
.D(n_1628),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1747),
.B(n_1443),
.Y(n_1749)
);

NOR2x1_ASAP7_75t_L g1750 ( 
.A(n_1745),
.B(n_1585),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1744),
.A2(n_1740),
.B1(n_1743),
.B2(n_1746),
.C(n_1748),
.Y(n_1751)
);

OAI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1750),
.B(n_1749),
.C(n_1526),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1565),
.B1(n_1561),
.B2(n_1566),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1753),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1753),
.A2(n_1566),
.B1(n_1556),
.B2(n_1570),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1754),
.A2(n_1620),
.B(n_1629),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1755),
.A2(n_1461),
.B1(n_1451),
.B2(n_1452),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1756),
.A2(n_1461),
.B(n_1452),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1757),
.Y(n_1759)
);

OAI32xp33_ASAP7_75t_L g1760 ( 
.A1(n_1759),
.A2(n_1585),
.A3(n_1572),
.B1(n_1534),
.B2(n_1530),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1760),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1761),
.Y(n_1762)
);

OAI221xp5_ASAP7_75t_R g1763 ( 
.A1(n_1762),
.A2(n_1758),
.B1(n_1547),
.B2(n_1526),
.C(n_1540),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1498),
.B(n_1476),
.C(n_1461),
.Y(n_1764)
);


endmodule