module fake_jpeg_18478_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_8),
.B(n_29),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_3),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_77),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_84),
.Y(n_87)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_53),
.Y(n_96)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_96),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_68),
.B1(n_67),
.B2(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_93),
.B1(n_67),
.B2(n_63),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_66),
.B1(n_63),
.B2(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_103),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_56),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_78),
.B1(n_75),
.B2(n_52),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_106),
.B1(n_7),
.B2(n_12),
.Y(n_128)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_5),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_50),
.B1(n_55),
.B2(n_70),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_4),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_74),
.B1(n_51),
.B2(n_59),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_61),
.B1(n_64),
.B2(n_62),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_125),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_121),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_73),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_25),
.CI(n_28),
.CON(n_137),
.SN(n_137)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_123),
.B1(n_128),
.B2(n_22),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_4),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_57),
.B1(n_58),
.B2(n_30),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_6),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_7),
.Y(n_127)
);

OR2x4_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_31),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_15),
.C(n_17),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_133),
.Y(n_142)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_135),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_18),
.C(n_20),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_131),
.B(n_139),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_130),
.B(n_137),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_144),
.A2(n_138),
.B(n_141),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_149),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_147),
.B(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_156),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_132),
.B(n_33),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_32),
.B(n_37),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_38),
.B(n_40),
.C(n_46),
.D(n_47),
.Y(n_160)
);

AOI321xp33_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_48),
.A3(n_114),
.B1(n_128),
.B2(n_122),
.C(n_142),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);


endmodule