module fake_jpeg_31083_n_465 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_465);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_465;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_31),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_19),
.A2(n_7),
.B1(n_12),
.B2(n_10),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_17),
.B1(n_16),
.B2(n_43),
.Y(n_143)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_6),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_68),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_28),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_79),
.Y(n_119)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_41),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_95),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_21),
.B(n_6),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_28),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_27),
.B(n_6),
.CON(n_97),
.SN(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_30),
.B(n_46),
.C(n_43),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_23),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_109),
.B(n_116),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_53),
.A2(n_36),
.B1(n_47),
.B2(n_34),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_115),
.A2(n_143),
.B1(n_37),
.B2(n_39),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_33),
.B(n_42),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_135),
.C(n_142),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_41),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_133),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_36),
.B1(n_47),
.B2(n_34),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_72),
.B1(n_74),
.B2(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_48),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_57),
.B(n_48),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_61),
.B(n_17),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_104),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_40),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_83),
.A2(n_47),
.B1(n_36),
.B2(n_30),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_153),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_47),
.B1(n_30),
.B2(n_29),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_29),
.B1(n_43),
.B2(n_46),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_56),
.A2(n_46),
.B1(n_29),
.B2(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_16),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_177),
.Y(n_207)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_160),
.A2(n_196),
.B1(n_138),
.B2(n_118),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_109),
.A2(n_66),
.B(n_78),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_161),
.A2(n_183),
.B(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_130),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_162),
.B(n_181),
.Y(n_218)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_96),
.B1(n_73),
.B2(n_71),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_164),
.A2(n_4),
.B(n_8),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_165),
.B(n_171),
.Y(n_241)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_77),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_119),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_172),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_175),
.B(n_178),
.Y(n_205)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_112),
.B(n_37),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_128),
.A2(n_85),
.B1(n_39),
.B2(n_42),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_188),
.B1(n_189),
.B2(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_54),
.C(n_86),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_155),
.C(n_4),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_77),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_182),
.B(n_184),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_115),
.A2(n_33),
.B1(n_38),
.B2(n_35),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_124),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_5),
.B(n_12),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_123),
.B(n_35),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_200),
.Y(n_209)
);

BUFx2_ASAP7_75t_SL g188 ( 
.A(n_155),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_190),
.B(n_193),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_106),
.A2(n_81),
.B1(n_76),
.B2(n_75),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_197),
.B1(n_198),
.B2(n_138),
.Y(n_232)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_38),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_110),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_111),
.A2(n_49),
.B1(n_67),
.B2(n_93),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_126),
.A2(n_93),
.B1(n_67),
.B2(n_9),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_99),
.A2(n_87),
.B1(n_8),
.B2(n_9),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_202),
.B(n_204),
.Y(n_235)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_203),
.Y(n_228)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_113),
.B(n_5),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_129),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_153),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_211),
.C(n_220),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_146),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_157),
.A2(n_125),
.B1(n_147),
.B2(n_113),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_213),
.A2(n_221),
.B1(n_232),
.B2(n_218),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_242),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_225),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_108),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_181),
.A2(n_108),
.B1(n_140),
.B2(n_103),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_183),
.A2(n_103),
.B1(n_140),
.B2(n_114),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_223),
.A2(n_234),
.B1(n_197),
.B2(n_162),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_161),
.A2(n_141),
.B(n_155),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_237),
.B(n_174),
.Y(n_261)
);

NAND3xp33_ASAP7_75t_SL g225 ( 
.A(n_185),
.B(n_107),
.C(n_144),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_177),
.B(n_144),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_4),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_107),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_160),
.A2(n_110),
.B1(n_130),
.B2(n_12),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_0),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_156),
.B(n_173),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_166),
.B(n_8),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_244),
.B(n_255),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_164),
.B1(n_180),
.B2(n_191),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_245),
.A2(n_248),
.B1(n_253),
.B2(n_259),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_164),
.B1(n_176),
.B2(n_193),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_246),
.A2(n_271),
.B1(n_273),
.B2(n_212),
.Y(n_290)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_210),
.A2(n_173),
.B(n_187),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_276),
.B(n_237),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_163),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_257),
.Y(n_307)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_164),
.B1(n_189),
.B2(n_169),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

AO22x1_ASAP7_75t_SL g257 ( 
.A1(n_211),
.A2(n_201),
.B1(n_200),
.B2(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_218),
.A2(n_159),
.B1(n_168),
.B2(n_158),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_228),
.B(n_202),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_260),
.B(n_264),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_243),
.B(n_242),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_209),
.B(n_235),
.Y(n_297)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_167),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_265),
.B(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_218),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

HAxp5_ASAP7_75t_SL g274 ( 
.A(n_229),
.B(n_14),
.CON(n_274),
.SN(n_274)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_224),
.A2(n_14),
.B(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_227),
.B(n_0),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_220),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_279),
.A2(n_281),
.B(n_296),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_219),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_282),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_288),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_207),
.C(n_209),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_302),
.C(n_306),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_249),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_294),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_295),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_255),
.A2(n_243),
.B1(n_233),
.B2(n_213),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_297),
.A2(n_276),
.B(n_273),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_221),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_245),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_230),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_250),
.B(n_241),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_304),
.B(n_302),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_240),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_271),
.A2(n_234),
.B1(n_214),
.B2(n_240),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_256),
.B1(n_262),
.B2(n_261),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_300),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_316),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_SL g356 ( 
.A1(n_318),
.A2(n_334),
.B(n_247),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_332),
.B1(n_336),
.B2(n_299),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_257),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_325),
.Y(n_349)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_324),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_278),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_327),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_304),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_330),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_256),
.C(n_250),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_333),
.C(n_284),
.Y(n_341)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_263),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_286),
.A2(n_307),
.B1(n_281),
.B2(n_301),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_253),
.C(n_254),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_335),
.B(n_283),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_286),
.A2(n_257),
.B1(n_248),
.B2(n_259),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_299),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_337),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_283),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_347),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_318),
.A2(n_308),
.B1(n_297),
.B2(n_279),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_346),
.B1(n_354),
.B2(n_356),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_342),
.C(n_350),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_294),
.C(n_306),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_315),
.A2(n_257),
.B1(n_293),
.B2(n_300),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_293),
.C(n_267),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_352),
.A2(n_360),
.B1(n_362),
.B2(n_337),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_322),
.A2(n_298),
.B1(n_280),
.B2(n_291),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_269),
.C(n_270),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_311),
.C(n_333),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_280),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_311),
.Y(n_378)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_359),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_303),
.B1(n_275),
.B2(n_272),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_319),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_363),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_275),
.B1(n_272),
.B2(n_216),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_315),
.A2(n_216),
.B1(n_233),
.B2(n_266),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_367),
.B(n_369),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_351),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_382),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_351),
.A2(n_313),
.B(n_333),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_371),
.A2(n_309),
.B(n_334),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_340),
.Y(n_372)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_372),
.Y(n_390)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_364),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_329),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_386),
.Y(n_396)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_380),
.C(n_378),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_381),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_358),
.C(n_350),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_342),
.B(n_313),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_339),
.B(n_332),
.CI(n_321),
.CON(n_382),
.SN(n_382)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_383),
.A2(n_354),
.B1(n_348),
.B2(n_357),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_353),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_385),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_353),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_311),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_379),
.A2(n_352),
.B1(n_360),
.B2(n_349),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_388),
.A2(n_400),
.B1(n_368),
.B2(n_344),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_387),
.A2(n_346),
.B(n_338),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_403),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_404),
.C(n_365),
.Y(n_412)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_371),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_379),
.A2(n_309),
.B(n_344),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_395),
.A2(n_367),
.B(n_370),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_383),
.A2(n_348),
.B1(n_327),
.B2(n_357),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_382),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_387),
.A2(n_349),
.B1(n_362),
.B2(n_324),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_359),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_335),
.C(n_312),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_407),
.B(n_410),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_419),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_404),
.B(n_366),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_411),
.B(n_412),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_416),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_382),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_414),
.B(n_417),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_388),
.A2(n_363),
.B1(n_372),
.B2(n_340),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_415),
.A2(n_402),
.B1(n_398),
.B2(n_390),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_393),
.A2(n_381),
.B1(n_373),
.B2(n_386),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_343),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_377),
.C(n_365),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_396),
.C(n_394),
.Y(n_426)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_398),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_331),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_396),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_410),
.A2(n_395),
.B(n_402),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_421),
.A2(n_323),
.B(n_310),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_407),
.A2(n_397),
.B1(n_392),
.B2(n_399),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_427),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_394),
.C(n_420),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_406),
.A2(n_389),
.B1(n_400),
.B2(n_373),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_429),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_343),
.B1(n_328),
.B2(n_317),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_416),
.A2(n_330),
.B1(n_326),
.B2(n_325),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_310),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_432),
.B(n_425),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_424),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_434),
.B(n_439),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_408),
.Y(n_436)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_436),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_422),
.A2(n_412),
.B(n_418),
.Y(n_437)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_437),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_440),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_441),
.B(n_444),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_310),
.C(n_258),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_442),
.B(n_443),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_252),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_439),
.A2(n_425),
.B(n_433),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_444),
.C(n_442),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_453),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_450),
.B(n_435),
.C(n_433),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_438),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_SL g458 ( 
.A(n_454),
.B(n_449),
.C(n_432),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

AOI31xp33_ASAP7_75t_L g457 ( 
.A1(n_455),
.A2(n_456),
.A3(n_449),
.B(n_447),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_429),
.B(n_423),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_457),
.B(n_458),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_459),
.B(n_206),
.Y(n_461)
);

AO21x1_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_206),
.B(n_208),
.Y(n_462)
);

OAI321xp33_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_460),
.A3(n_14),
.B1(n_2),
.B2(n_1),
.C(n_0),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_463),
.A2(n_1),
.B1(n_2),
.B2(n_344),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_464),
.B(n_2),
.Y(n_465)
);


endmodule