module fake_jpeg_30529_n_48 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_48);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_48;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_18),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_24),
.C(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_18),
.B1(n_17),
.B2(n_21),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_29),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_13),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_1),
.B(n_2),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_2),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_12),
.C(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_31),
.B(n_5),
.Y(n_42)
);

NOR2x1p5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_4),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_38),
.C(n_40),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B(n_43),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_42),
.B1(n_8),
.B2(n_9),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_7),
.C(n_8),
.Y(n_48)
);


endmodule