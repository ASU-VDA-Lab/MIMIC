module fake_jpeg_11063_n_454 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_454);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_454;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_11),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_3),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_59),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_61),
.Y(n_171)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_64),
.B(n_67),
.Y(n_142)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_65),
.Y(n_168)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_31),
.CON(n_66),
.SN(n_66)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_66),
.B(n_108),
.Y(n_166)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_69),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_71),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_72),
.B(n_80),
.Y(n_155)
);

INVx11_ASAP7_75t_SL g73 ( 
.A(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_76),
.B(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_25),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_81),
.Y(n_181)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_83),
.B(n_86),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_15),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_89),
.B(n_94),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_90),
.B(n_100),
.Y(n_148)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_98),
.B(n_104),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_23),
.B(n_0),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_23),
.B(n_1),
.Y(n_100)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_101),
.Y(n_164)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_35),
.B(n_52),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_107),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_35),
.B(n_1),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_17),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_111),
.B(n_112),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_17),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_38),
.B(n_1),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_113),
.B(n_97),
.Y(n_169)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_114),
.A2(n_101),
.B(n_65),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_47),
.B1(n_39),
.B2(n_24),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_66),
.A2(n_47),
.B1(n_39),
.B2(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_119),
.A2(n_140),
.B1(n_154),
.B2(n_158),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_27),
.B1(n_51),
.B2(n_49),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_120),
.A2(n_162),
.B1(n_185),
.B2(n_186),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_50),
.B1(n_29),
.B2(n_49),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_50),
.B1(n_52),
.B2(n_45),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_45),
.B1(n_42),
.B2(n_40),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_132),
.A2(n_149),
.B1(n_151),
.B2(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_42),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_58),
.B1(n_63),
.B2(n_77),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_40),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_38),
.B1(n_17),
.B2(n_3),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_82),
.A2(n_17),
.B1(n_2),
.B2(n_5),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_1),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_184),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_103),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_79),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_74),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_92),
.A2(n_12),
.B1(n_96),
.B2(n_106),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_178),
.B1(n_116),
.B2(n_174),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_60),
.A2(n_102),
.B1(n_88),
.B2(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_179),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_170),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_87),
.A2(n_91),
.B1(n_97),
.B2(n_56),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

OA22x2_ASAP7_75t_SL g174 ( 
.A1(n_69),
.A2(n_73),
.B1(n_68),
.B2(n_61),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_116),
.B(n_144),
.C(n_182),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_56),
.A2(n_70),
.B1(n_67),
.B2(n_115),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_69),
.B(n_61),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_100),
.B(n_90),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_58),
.A2(n_92),
.B1(n_77),
.B2(n_74),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_100),
.A2(n_90),
.B1(n_76),
.B2(n_66),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_190),
.B(n_194),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_192),
.B(n_229),
.Y(n_288)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_184),
.B(n_148),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_135),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_196),
.B(n_197),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_138),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_198),
.B(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

BUFx4f_ASAP7_75t_SL g201 ( 
.A(n_168),
.Y(n_201)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_202),
.B(n_205),
.Y(n_273)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_204),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_142),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_136),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_206),
.B(n_207),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_164),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_168),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_209),
.B(n_215),
.Y(n_285)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_211),
.B(n_212),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_168),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_213),
.A2(n_118),
.B1(n_124),
.B2(n_129),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_119),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_233),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_217),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_131),
.B(n_157),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_120),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_219),
.B(n_226),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_220),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_137),
.B(n_178),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_150),
.Y(n_226)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_131),
.B(n_157),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_150),
.Y(n_231)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_137),
.B(n_154),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_241),
.Y(n_269)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_245),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_161),
.B(n_133),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_236),
.Y(n_275)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_171),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_238),
.Y(n_280)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_128),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_128),
.B(n_183),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_160),
.B(n_158),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_129),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_242),
.Y(n_277)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_243),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_246),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_118),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_204),
.Y(n_279)
);

OR2x2_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_174),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_248),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_185),
.B1(n_175),
.B2(n_145),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_250),
.A2(n_272),
.B1(n_283),
.B2(n_199),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_255),
.A2(n_270),
.B1(n_271),
.B2(n_222),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_195),
.B(n_124),
.C(n_167),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_226),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_192),
.A2(n_139),
.B(n_145),
.C(n_156),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_267),
.A2(n_217),
.B(n_231),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_225),
.A2(n_156),
.B1(n_167),
.B2(n_139),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_232),
.A2(n_241),
.B1(n_219),
.B2(n_227),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_228),
.A2(n_189),
.B1(n_200),
.B2(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_228),
.A2(n_189),
.B1(n_200),
.B2(n_198),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_234),
.B(n_188),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_229),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_205),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_302),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_295),
.A2(n_297),
.B1(n_307),
.B2(n_265),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_187),
.B(n_191),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_298),
.B(n_265),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_208),
.B1(n_193),
.B2(n_210),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_301),
.B1(n_255),
.B2(n_300),
.Y(n_335)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_283),
.B1(n_250),
.B2(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_258),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_263),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_312),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_305),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_202),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_246),
.B1(n_243),
.B2(n_233),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_253),
.B(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_309),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_247),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_269),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_315),
.Y(n_338)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_311),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_253),
.B(n_201),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_220),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_313),
.A2(n_320),
.B(n_296),
.Y(n_342)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_260),
.B(n_224),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_221),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_259),
.C(n_274),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_270),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_223),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_323),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_249),
.B(n_203),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_319),
.B(n_278),
.Y(n_351)
);

A2O1A1O1Ixp25_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_201),
.B(n_236),
.C(n_238),
.D(n_244),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_280),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_249),
.B(n_288),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_284),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_294),
.B(n_284),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_278),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_325),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_326),
.B(n_342),
.Y(n_375)
);

BUFx12f_ASAP7_75t_SL g327 ( 
.A(n_306),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_345),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_287),
.B(n_265),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_297),
.C(n_319),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_348),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_335),
.A2(n_309),
.B1(n_298),
.B2(n_304),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_337),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_340),
.A2(n_299),
.B1(n_301),
.B2(n_313),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_295),
.A2(n_248),
.B1(n_267),
.B2(n_275),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_344),
.A2(n_352),
.B1(n_320),
.B2(n_308),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_323),
.A2(n_273),
.B(n_267),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_290),
.B(n_261),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_315),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_292),
.A2(n_266),
.B1(n_254),
.B2(n_257),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_317),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_368),
.C(n_373),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_357),
.A2(n_374),
.B1(n_376),
.B2(n_348),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_344),
.A2(n_313),
.B1(n_303),
.B2(n_312),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_363),
.B(n_364),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_359),
.B(n_305),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_334),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_360),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_324),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_369),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_332),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_362),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_331),
.A2(n_325),
.B1(n_293),
.B2(n_292),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_333),
.A2(n_318),
.B1(n_320),
.B2(n_316),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_332),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_365),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_350),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_372),
.A2(n_328),
.B1(n_326),
.B2(n_352),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_346),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_321),
.B1(n_314),
.B2(n_311),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_370),
.A2(n_342),
.B(n_337),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_330),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_389),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_346),
.C(n_329),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_388),
.C(n_359),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_356),
.A2(n_345),
.B(n_335),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_394),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_385),
.A2(n_387),
.B1(n_372),
.B2(n_394),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_357),
.A2(n_336),
.B1(n_353),
.B2(n_349),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_351),
.C(n_353),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_349),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_390),
.A2(n_358),
.B1(n_364),
.B2(n_375),
.Y(n_397)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_374),
.A2(n_347),
.B1(n_350),
.B2(n_343),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_363),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_397),
.A2(n_403),
.B1(n_385),
.B2(n_387),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_406),
.Y(n_414)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_400),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_302),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_402),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_386),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_383),
.Y(n_403)
);

OAI21x1_ASAP7_75t_SL g404 ( 
.A1(n_383),
.A2(n_361),
.B(n_368),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_404),
.A2(n_377),
.B(n_390),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_356),
.C(n_366),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_410),
.C(n_382),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_347),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_405),
.C(n_406),
.Y(n_428)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_381),
.C(n_388),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_418),
.Y(n_429)
);

BUFx24_ASAP7_75t_SL g417 ( 
.A(n_410),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_398),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_395),
.C(n_389),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_397),
.A2(n_379),
.B1(n_392),
.B2(n_386),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_419),
.B(n_420),
.Y(n_431)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_400),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_421),
.A2(n_405),
.B(n_408),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_422),
.A2(n_399),
.B(n_378),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_423),
.A2(n_426),
.B(n_430),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_425),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_422),
.A2(n_407),
.B1(n_399),
.B2(n_377),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_414),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_412),
.A2(n_384),
.B(n_392),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_415),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_433),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_367),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_429),
.B(n_411),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_437),
.B(n_371),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_423),
.A2(n_409),
.B1(n_384),
.B2(n_418),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_439),
.C(n_431),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_416),
.C(n_414),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_426),
.C(n_430),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_440),
.Y(n_449)
);

AO21x1_ASAP7_75t_L g447 ( 
.A1(n_441),
.A2(n_442),
.B(n_445),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_438),
.A2(n_384),
.B1(n_376),
.B2(n_391),
.Y(n_443)
);

AOI322xp5_ASAP7_75t_L g448 ( 
.A1(n_443),
.A2(n_256),
.A3(n_262),
.B1(n_281),
.B2(n_289),
.C1(n_276),
.C2(n_282),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_435),
.A2(n_391),
.B(n_341),
.Y(n_445)
);

AOI322xp5_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_436),
.A3(n_435),
.B1(n_343),
.B2(n_291),
.C1(n_281),
.C2(n_289),
.Y(n_446)
);

OAI321xp33_ASAP7_75t_L g450 ( 
.A1(n_446),
.A2(n_448),
.A3(n_256),
.B1(n_262),
.B2(n_281),
.C(n_261),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_450),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_449),
.B(n_440),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_451),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_447),
.Y(n_454)
);


endmodule