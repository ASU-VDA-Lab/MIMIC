module fake_jpeg_16403_n_293 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_36),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_23),
.B1(n_28),
.B2(n_15),
.Y(n_41)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_56),
.B1(n_29),
.B2(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_28),
.B1(n_15),
.B2(n_17),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_29),
.B1(n_39),
.B2(n_17),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_23),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_29),
.B1(n_17),
.B2(n_16),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_21),
.B(n_20),
.C(n_16),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_18),
.Y(n_84)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_67),
.B1(n_73),
.B2(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_21),
.B1(n_20),
.B2(n_16),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_39),
.B1(n_23),
.B2(n_21),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_33),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_75),
.B(n_79),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_45),
.B1(n_39),
.B2(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_48),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_33),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_53),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_97),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_100),
.B(n_18),
.Y(n_129)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_93),
.B(n_71),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_73),
.B1(n_93),
.B2(n_75),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_81),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_105),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_48),
.B1(n_45),
.B2(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_107),
.B1(n_78),
.B2(n_88),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_48),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_79),
.C(n_85),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_71),
.B(n_86),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_109),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_53),
.B1(n_35),
.B2(n_25),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_65),
.B1(n_83),
.B2(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_126),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_123),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_116),
.B(n_129),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_124),
.B1(n_90),
.B2(n_91),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_128),
.B1(n_95),
.B2(n_103),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_71),
.B(n_86),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_27),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_74),
.C(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_58),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_85),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_19),
.C(n_30),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_72),
.B1(n_35),
.B2(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_83),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_91),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_111),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_138),
.B(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_90),
.B1(n_108),
.B2(n_92),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_103),
.B1(n_96),
.B2(n_100),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_108),
.B(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_14),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_126),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_114),
.C(n_128),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_27),
.B(n_22),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_131),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_157),
.Y(n_173)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_123),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_133),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_163),
.C(n_167),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_125),
.B1(n_129),
.B2(n_119),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_161),
.A2(n_178),
.B1(n_181),
.B2(n_154),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_116),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_170),
.B(n_178),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_112),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_59),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_176),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_153),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_131),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_179),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_117),
.B1(n_118),
.B2(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_136),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_117),
.B1(n_83),
.B2(n_27),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_122),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_145),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_149),
.B1(n_139),
.B2(n_146),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_185),
.A2(n_188),
.B1(n_202),
.B2(n_203),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_199),
.C(n_175),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_158),
.B(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_144),
.B(n_159),
.Y(n_197)
);

OAI31xp33_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_168),
.A3(n_19),
.B(n_30),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_201),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_142),
.B(n_150),
.C(n_141),
.Y(n_200)
);

AOI21x1_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_193),
.B(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_156),
.B(n_142),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_140),
.B1(n_22),
.B2(n_49),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_181),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_30),
.C(n_19),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_182),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_0),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_217),
.B(n_203),
.C(n_188),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_160),
.C(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_214),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_170),
.C(n_172),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_184),
.C(n_166),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_52),
.C(n_58),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_219),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_52),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_52),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_26),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_191),
.B(n_200),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_200),
.B(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_207),
.B1(n_185),
.B2(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_210),
.B1(n_218),
.B2(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_19),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_243),
.C(n_59),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_30),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_209),
.B1(n_216),
.B2(n_214),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_22),
.Y(n_259)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_269)
);

AO221x1_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_243),
.B1(n_228),
.B2(n_241),
.C(n_229),
.Y(n_251)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_255),
.C(n_232),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_229),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_254),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_58),
.C(n_49),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_268),
.C(n_252),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_263),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_26),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_26),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_11),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_244),
.B(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_26),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_250),
.B(n_26),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_269),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_11),
.Y(n_268)
);

AOI31xp67_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_264),
.A3(n_259),
.B(n_265),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_278),
.C(n_268),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_245),
.A3(n_255),
.B1(n_49),
.B2(n_35),
.C1(n_59),
.C2(n_10),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_274),
.B(n_276),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_10),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_35),
.A3(n_11),
.B1(n_12),
.B2(n_6),
.C1(n_8),
.C2(n_13),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_18),
.C(n_8),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_4),
.B(n_5),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_263),
.C(n_260),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_284),
.B(n_4),
.Y(n_288)
);

OAI211xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_275),
.B(n_277),
.C(n_270),
.Y(n_284)
);

A2O1A1O1Ixp25_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_8),
.B(n_12),
.C(n_13),
.D(n_3),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_280),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_287),
.A2(n_288),
.B(n_5),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_290),
.C(n_18),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_5),
.B(n_285),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_5),
.Y(n_293)
);


endmodule