module fake_jpeg_13622_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_54),
.Y(n_156)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_61),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_63),
.B(n_73),
.Y(n_144)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_30),
.A2(n_45),
.B1(n_47),
.B2(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_102),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_25),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_105),
.Y(n_124)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_82),
.B(n_92),
.Y(n_167)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_100),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_98),
.B(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_43),
.B(n_17),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_46),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_103),
.B(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_48),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_15),
.Y(n_105)
);

BUFx4f_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_49),
.B(n_15),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_53),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_114),
.Y(n_175)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_87),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_54),
.B(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_138),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_79),
.A2(n_44),
.B1(n_39),
.B2(n_41),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_132),
.A2(n_44),
.B1(n_51),
.B2(n_29),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_55),
.B(n_48),
.Y(n_138)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_58),
.Y(n_143)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_35),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_58),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_150),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_89),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_89),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_155),
.B(n_160),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_62),
.A2(n_35),
.B(n_37),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_22),
.B(n_28),
.C(n_33),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_85),
.B(n_37),
.Y(n_170)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_65),
.B1(n_84),
.B2(n_95),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_174),
.A2(n_181),
.B1(n_184),
.B2(n_191),
.Y(n_245)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_177),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_179),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_101),
.B1(n_96),
.B2(n_93),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_91),
.B1(n_88),
.B2(n_76),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_185),
.B(n_214),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_173),
.Y(n_186)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_189),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_67),
.B1(n_74),
.B2(n_28),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_192),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_124),
.B(n_126),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_197),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_135),
.A2(n_44),
.B1(n_86),
.B2(n_40),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_195),
.A2(n_169),
.B1(n_123),
.B2(n_109),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_22),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_142),
.B(n_41),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_198),
.B(n_108),
.Y(n_260)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_199),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_200),
.A2(n_209),
.B1(n_224),
.B2(n_226),
.Y(n_264)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_132),
.A2(n_40),
.B1(n_29),
.B2(n_27),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_204),
.A2(n_134),
.B1(n_163),
.B2(n_172),
.Y(n_259)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_53),
.C(n_33),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_231),
.C(n_236),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_142),
.A2(n_51),
.B1(n_40),
.B2(n_27),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_157),
.B(n_12),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_144),
.B(n_50),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_217),
.B(n_225),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_112),
.Y(n_218)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_235),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_151),
.A2(n_51),
.B1(n_40),
.B2(n_27),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_117),
.B(n_50),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_151),
.A2(n_51),
.B1(n_29),
.B2(n_27),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_147),
.B(n_42),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_227),
.B(n_229),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_113),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_110),
.B(n_156),
.C(n_125),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_147),
.Y(n_232)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_147),
.B(n_42),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_110),
.B(n_38),
.C(n_51),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_190),
.A2(n_134),
.B(n_145),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_243),
.A2(n_258),
.B(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_180),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_249),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_175),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_198),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_250),
.B(n_256),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_251),
.A2(n_148),
.B1(n_163),
.B2(n_228),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_38),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_SL g258 ( 
.A(n_185),
.B(n_153),
.C(n_151),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_259),
.A2(n_271),
.B1(n_275),
.B2(n_212),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_260),
.B(n_216),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_206),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_265),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_187),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_202),
.B(n_136),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_207),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_200),
.A2(n_141),
.B1(n_109),
.B2(n_133),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_205),
.A2(n_141),
.B1(n_133),
.B2(n_172),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_188),
.B(n_136),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_201),
.B(n_158),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_220),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_286),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_194),
.B(n_233),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_282),
.B(n_283),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_194),
.B(n_140),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_125),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_221),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_228),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_SL g289 ( 
.A(n_224),
.B(n_123),
.C(n_115),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_269),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_291),
.B(n_304),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_238),
.A2(n_218),
.B1(n_196),
.B2(n_290),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_270),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_297),
.B(n_306),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_247),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_262),
.C(n_261),
.Y(n_341)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_299),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_238),
.A2(n_108),
.B1(n_131),
.B2(n_232),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_239),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_270),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_280),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_307),
.B(n_310),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_264),
.B1(n_289),
.B2(n_252),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_308),
.A2(n_328),
.B1(n_237),
.B2(n_267),
.Y(n_346)
);

INVx13_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx3_ASAP7_75t_SL g355 ( 
.A(n_309),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_242),
.Y(n_310)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_324),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_243),
.A2(n_207),
.B(n_219),
.C(n_111),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_314),
.A2(n_321),
.B(n_337),
.Y(n_379)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_327),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_317),
.B(n_319),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_250),
.A2(n_209),
.B(n_226),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_318),
.A2(n_245),
.B(n_215),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_260),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_248),
.B(n_195),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_320),
.B(n_322),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_247),
.A2(n_111),
.B(n_208),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_111),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_323),
.Y(n_351)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_325),
.A2(n_326),
.B1(n_245),
.B2(n_276),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_14),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_254),
.A2(n_216),
.B1(n_215),
.B2(n_233),
.Y(n_328)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_329),
.Y(n_378)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_333),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_259),
.A2(n_148),
.B1(n_189),
.B2(n_199),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_332),
.A2(n_334),
.B1(n_285),
.B2(n_276),
.Y(n_363)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_257),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_271),
.A2(n_210),
.B1(n_203),
.B2(n_183),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_275),
.Y(n_353)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_338),
.Y(n_342)
);

OR2x4_ASAP7_75t_L g337 ( 
.A(n_258),
.B(n_284),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_279),
.B(n_208),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_343),
.C(n_350),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_244),
.C(n_266),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_291),
.B(n_305),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_360),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_346),
.A2(n_348),
.B(n_362),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_272),
.B(n_287),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_284),
.C(n_240),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_320),
.A2(n_318),
.B1(n_312),
.B2(n_304),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_352),
.A2(n_354),
.B1(n_323),
.B2(n_300),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_353),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_312),
.A2(n_245),
.B1(n_253),
.B2(n_223),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_267),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_303),
.Y(n_388)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_245),
.Y(n_360)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_307),
.B(n_285),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_374),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_319),
.A2(n_208),
.B(n_215),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_369),
.A2(n_370),
.B(n_335),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_322),
.A2(n_162),
.B(n_52),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_241),
.B1(n_162),
.B2(n_12),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_373),
.A2(n_377),
.B1(n_306),
.B2(n_330),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_315),
.B(n_241),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_334),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_372),
.B(n_310),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_383),
.B(n_387),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_360),
.A2(n_325),
.B(n_332),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_SL g416 ( 
.A1(n_385),
.A2(n_362),
.B(n_353),
.C(n_351),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_293),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_400),
.C(n_407),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_365),
.B(n_295),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_388),
.B(n_342),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_314),
.B(n_295),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_389),
.A2(n_395),
.B(n_398),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_343),
.B(n_331),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_394),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_391),
.Y(n_421)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

INVx13_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_331),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_379),
.A2(n_323),
.B(n_335),
.Y(n_395)
);

BUFx12f_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_396),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_348),
.A2(n_323),
.B(n_337),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_341),
.B(n_299),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_340),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_410),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_323),
.Y(n_403)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

INVx13_ASAP7_75t_L g404 ( 
.A(n_355),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_404),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_405),
.A2(n_409),
.B1(n_397),
.B2(n_384),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_352),
.B(n_297),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_336),
.Y(n_408)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_354),
.A2(n_300),
.B1(n_327),
.B2(n_316),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_412),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_340),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_359),
.A2(n_302),
.B1(n_294),
.B2(n_296),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_413),
.A2(n_414),
.B(n_378),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_359),
.A2(n_333),
.B1(n_324),
.B2(n_311),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_342),
.B(n_309),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_415),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_416),
.A2(n_441),
.B(n_446),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_349),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_419),
.C(n_422),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_356),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_351),
.C(n_368),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_426),
.A2(n_428),
.B1(n_436),
.B2(n_385),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_382),
.A2(n_363),
.B1(n_346),
.B2(n_375),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_431),
.B(n_444),
.Y(n_450)
);

NOR2x1p5_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_382),
.A2(n_366),
.B1(n_347),
.B2(n_374),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_369),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_442),
.C(n_443),
.Y(n_461)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_386),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_402),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_406),
.A2(n_347),
.B(n_370),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_381),
.B(n_371),
.C(n_358),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_358),
.C(n_367),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_403),
.B(n_364),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_447),
.A2(n_454),
.B1(n_432),
.B2(n_416),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_396),
.Y(n_448)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_408),
.Y(n_453)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_428),
.A2(n_385),
.B1(n_397),
.B2(n_398),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_431),
.B(n_405),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_455),
.B(n_416),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_396),
.Y(n_457)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_457),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_419),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_459),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_389),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_423),
.A2(n_391),
.B1(n_392),
.B2(n_406),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_460),
.A2(n_425),
.B1(n_434),
.B2(n_329),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_464),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_420),
.A2(n_409),
.B1(n_413),
.B2(n_402),
.Y(n_463)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_423),
.A2(n_380),
.B(n_395),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_433),
.A2(n_446),
.B1(n_439),
.B2(n_441),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_465),
.A2(n_468),
.B1(n_469),
.B2(n_436),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_424),
.A2(n_414),
.B1(n_377),
.B2(n_410),
.Y(n_466)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_466),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_427),
.A2(n_364),
.B1(n_367),
.B2(n_376),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_432),
.A2(n_376),
.B1(n_355),
.B2(n_361),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_393),
.Y(n_470)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_470),
.Y(n_494)
);

XOR2x1_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_404),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_434),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_355),
.C(n_309),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_438),
.C(n_442),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_473),
.A2(n_486),
.B1(n_468),
.B2(n_456),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_476),
.A2(n_464),
.B1(n_461),
.B2(n_456),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_461),
.A2(n_421),
.B(n_443),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_478),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_481),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_469),
.A2(n_426),
.B1(n_416),
.B2(n_435),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_482),
.A2(n_490),
.B1(n_454),
.B2(n_447),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_484),
.B(n_485),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_451),
.B(n_0),
.C(n_2),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_2),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_449),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_0),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_450),
.Y(n_511)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_480),
.Y(n_495)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_497),
.B1(n_506),
.B2(n_508),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_498),
.B(n_501),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_SL g499 ( 
.A(n_475),
.B(n_479),
.C(n_451),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_505),
.Y(n_520)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_503),
.B(n_504),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_483),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_472),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g506 ( 
.A(n_484),
.B(n_455),
.CI(n_450),
.CON(n_506),
.SN(n_506)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_509),
.Y(n_514)
);

INVx13_ASAP7_75t_L g508 ( 
.A(n_487),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_478),
.A2(n_453),
.B(n_459),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_471),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_511),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_493),
.C(n_491),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_516),
.C(n_518),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_505),
.C(n_497),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_511),
.A2(n_473),
.B1(n_487),
.B2(n_467),
.Y(n_517)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_517),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_507),
.B(n_476),
.C(n_482),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_510),
.B(n_485),
.C(n_492),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_7),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_488),
.B1(n_490),
.B2(n_6),
.Y(n_521)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_521),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_506),
.A2(n_502),
.B1(n_5),
.B2(n_6),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_512),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_502),
.C(n_506),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_534),
.Y(n_540)
);

MAJx2_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_4),
.C(n_5),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_528),
.C(n_519),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_4),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_6),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_530),
.A2(n_533),
.B(n_8),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_532),
.B(n_523),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_7),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_537),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_526),
.A2(n_515),
.B(n_518),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_538),
.B(n_539),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_531),
.B(n_514),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_541),
.B(n_529),
.Y(n_544)
);

AOI21xp33_ASAP7_75t_L g546 ( 
.A1(n_544),
.A2(n_530),
.B(n_527),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_543),
.A2(n_540),
.B(n_535),
.Y(n_545)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_545),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_547),
.Y(n_548)
);

AOI322xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_542),
.A3(n_546),
.B1(n_514),
.B2(n_528),
.C1(n_525),
.C2(n_10),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_525),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_8),
.Y(n_552)
);


endmodule