module real_jpeg_25895_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx6_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_0),
.Y(n_146)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_0),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_0),
.B(n_2),
.Y(n_191)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_2),
.B(n_45),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_2),
.B(n_43),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_2),
.B(n_32),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_37),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_2),
.B(n_26),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_51),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_2),
.B(n_73),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_5),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_5),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_5),
.B(n_37),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_5),
.B(n_32),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_5),
.B(n_45),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_5),
.B(n_43),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_5),
.B(n_26),
.Y(n_316)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_7),
.B(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_7),
.B(n_26),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_32),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_8),
.B(n_45),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_37),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_8),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_8),
.B(n_43),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_8),
.B(n_26),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_8),
.B(n_51),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_8),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_9),
.B(n_37),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_32),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_155),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_9),
.B(n_45),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_9),
.B(n_43),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_9),
.B(n_26),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_9),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_9),
.B(n_98),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_10),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_10),
.B(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_10),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_10),
.B(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_10),
.B(n_202),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_10),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_10),
.B(n_32),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_12),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_12),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_12),
.B(n_51),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_12),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_12),
.B(n_37),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_13),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_13),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_13),
.B(n_37),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_13),
.B(n_32),
.Y(n_269)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_16),
.B(n_43),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_16),
.B(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_16),
.B(n_45),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_16),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_16),
.B(n_37),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_16),
.B(n_51),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_17),
.B(n_37),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_17),
.B(n_32),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_17),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_86),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_21),
.A2(n_22),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_62),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_23),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.C(n_47),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_24),
.B(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_SL g85 ( 
.A(n_25),
.B(n_31),
.C(n_34),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_30),
.A2(n_31),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_SL g93 ( 
.A(n_31),
.B(n_78),
.C(n_81),
.Y(n_93)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_32),
.Y(n_188)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_65),
.C(n_68),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_34),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_36),
.B(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_40),
.B(n_47),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_330),
.SN(n_330)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_43),
.Y(n_296)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_47),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_49),
.C(n_50),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_53),
.A2(n_62),
.B1(n_63),
.B2(n_367),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_53),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_58),
.C(n_61),
.Y(n_91)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_56),
.B(n_187),
.Y(n_246)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_56),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_71),
.C(n_74),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_64),
.B(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_65),
.A2(n_66),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_65),
.B(n_307),
.C(n_308),
.Y(n_329)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_68),
.B(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_70),
.B(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_340),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_74),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_74),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_74),
.B(n_336),
.C(n_339),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_75),
.B(n_86),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.C(n_85),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_76),
.A2(n_77),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_79),
.B(n_82),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_83),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_101),
.C(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_82),
.B(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_84),
.B(n_85),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.C(n_94),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_107),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_90),
.CI(n_91),
.CON(n_88),
.SN(n_88)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_101),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_368),
.C(n_369),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_356),
.C(n_357),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_344),
.C(n_345),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_320),
.C(n_321),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_287),
.C(n_288),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_252),
.C(n_253),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_222),
.C(n_223),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_196),
.C(n_197),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_158),
.C(n_169),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_141),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_129),
.B(n_136),
.C(n_141),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_131),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_137),
.B(n_139),
.C(n_140),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_142),
.B(n_150),
.C(n_151),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_145),
.Y(n_284)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_153),
.B(n_157),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_168),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_192),
.C(n_193),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.C(n_184),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.C(n_189),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_211),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_212),
.C(n_221),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_206),
.C(n_207),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_201),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_205),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_207),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.CI(n_210),
.CON(n_207),
.SN(n_207)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_209),
.C(n_210),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_219),
.B2(n_220),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_218),
.C(n_220),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_238),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.C(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_234),
.C(n_237),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_229),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.CI(n_232),
.CON(n_229),
.SN(n_229)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_231),
.C(n_232),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_245),
.C(n_250),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_245),
.B1(n_250),
.B2(n_251),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_241),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_244),
.B(n_277),
.C(n_278),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_273),
.B2(n_286),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_274),
.C(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_258),
.C(n_266),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_262),
.C(n_265),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_270),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_282),
.C(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_318),
.B2(n_319),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_289),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_309),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_309),
.C(n_318),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_300),
.C(n_301),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_295),
.C(n_297),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_304),
.B1(n_305),
.B2(n_308),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_302),
.Y(n_308)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_324),
.C(n_343),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_331),
.B2(n_343),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_329),
.C(n_330),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g376 ( 
.A(n_330),
.Y(n_376)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_331),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_342),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_339),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_355),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_349),
.C(n_355),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_352),
.C(n_353),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_360),
.C(n_365),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_364),
.B2(n_365),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_370),
.Y(n_371)
);


endmodule