module fake_jpeg_25572_n_200 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_9),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_20),
.B1(n_12),
.B2(n_17),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_10),
.B1(n_21),
.B2(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_25),
.B(n_24),
.C(n_22),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_35),
.B(n_22),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_30),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_47),
.B(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_28),
.B1(n_29),
.B2(n_20),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_52),
.B1(n_44),
.B2(n_47),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_53),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_11),
.B1(n_18),
.B2(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_21),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_66),
.Y(n_88)
);

NOR2x1p5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_47),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_43),
.B1(n_38),
.B2(n_53),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_40),
.B1(n_32),
.B2(n_45),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_66),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_25),
.B(n_26),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_68),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_43),
.C(n_24),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_90),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_43),
.A3(n_41),
.B1(n_35),
.B2(n_34),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_43),
.A3(n_65),
.B1(n_32),
.B2(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_11),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_63),
.B(n_64),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_103),
.B(n_107),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_102),
.B1(n_81),
.B2(n_34),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_90),
.B1(n_88),
.B2(n_78),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_34),
.B1(n_31),
.B2(n_14),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_105),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_71),
.B1(n_35),
.B2(n_41),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_65),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_75),
.B(n_85),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_67),
.B(n_18),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_116),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_31),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_122),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_136),
.B1(n_137),
.B2(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_106),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_104),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_113),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_103),
.B1(n_112),
.B2(n_14),
.Y(n_150)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_134),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_114),
.Y(n_142)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_31),
.B1(n_11),
.B2(n_18),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_111),
.B1(n_116),
.B2(n_103),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_144),
.B1(n_129),
.B2(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_147),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_93),
.B1(n_97),
.B2(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_149),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_108),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_97),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_150),
.A2(n_135),
.B1(n_117),
.B2(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_117),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_163),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_150),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_133),
.C(n_125),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_160),
.C(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_124),
.C(n_122),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_132),
.C(n_139),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_119),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_145),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_162),
.B1(n_159),
.B2(n_158),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_148),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_152),
.B(n_1),
.C(n_2),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_SL g176 ( 
.A(n_170),
.B(n_0),
.C(n_1),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_9),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_0),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_166),
.C(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_1),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_1),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_161),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_8),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_8),
.B1(n_14),
.B2(n_3),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_158),
.B1(n_173),
.B2(n_3),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_174),
.Y(n_190)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_177),
.Y(n_188)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_179),
.C(n_4),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_190),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_181),
.C(n_4),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_187),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_194),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_195),
.B(n_190),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_6),
.Y(n_200)
);


endmodule