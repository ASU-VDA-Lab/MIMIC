module real_jpeg_18801_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

NAND2x1_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_0),
.B(n_57),
.Y(n_123)
);

NAND2x1_ASAP7_75t_SL g124 ( 
.A(n_0),
.B(n_125),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_4),
.B(n_63),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_4),
.B(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_6),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_6),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_6),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_6),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_6),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_6),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_6),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_7),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_7),
.B(n_239),
.Y(n_238)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_223),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_147),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_127),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_16),
.B(n_127),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_17),
.B(n_83),
.C(n_115),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_52),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_40),
.B2(n_41),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_20),
.B(n_40),
.C(n_52),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_21),
.B(n_33),
.C(n_39),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.C(n_26),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_22),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_22),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_22),
.B(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_118),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_22),
.A2(n_77),
.B(n_78),
.C(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_22),
.A2(n_50),
.B1(n_78),
.B2(n_176),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_22),
.B(n_47),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_24),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

O2A1O1Ixp5_ASAP7_75t_L g70 ( 
.A1(n_26),
.A2(n_71),
.B(n_76),
.C(n_77),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_26),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_26),
.A2(n_76),
.B1(n_118),
.B2(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OR2x4_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_28),
.Y(n_239)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_31),
.A2(n_39),
.B1(n_43),
.B2(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_31),
.B(n_132),
.C(n_157),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_32),
.B(n_90),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_33),
.A2(n_34),
.B1(n_124),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_34),
.B(n_122),
.C(n_124),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_38),
.Y(n_141)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_43),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_43),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_43),
.A2(n_58),
.B1(n_60),
.B2(n_157),
.Y(n_259)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_46),
.B(n_50),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_49),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_65),
.C(n_69),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_53),
.B(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_55),
.A2(n_56),
.B1(n_171),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_55),
.A2(n_56),
.B1(n_67),
.B2(n_165),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_58),
.C(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_57),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_61),
.B(n_140),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_67),
.A2(n_160),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_67),
.A2(n_122),
.B(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_71),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_71),
.A2(n_132),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_78),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_78),
.A2(n_170),
.B(n_177),
.Y(n_212)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_115),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_98),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_84),
.B(n_100),
.C(n_102),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_86),
.B(n_89),
.C(n_93),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_89),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_97),
.B1(n_123),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_97),
.A2(n_159),
.B(n_160),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_140),
.C(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_104),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_126),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_126),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_118),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_118),
.B(n_197),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_122),
.B(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_124),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.C(n_145),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_128),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_145),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.C(n_138),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_131),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22x1_ASAP7_75t_SL g236 ( 
.A1(n_140),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_140),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_142),
.Y(n_183)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_222),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_217),
.B(n_221),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_205),
.B(n_216),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_186),
.B(n_204),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_167),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_167),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.C(n_163),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_163),
.B1(n_164),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_178),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_179),
.C(n_185),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_196),
.B(n_198),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_185),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_183),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_194),
.B(n_203),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_191),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_200),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_199),
.B(n_202),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_207),
.Y(n_216)
);

XOR2x2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_261),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_260),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_260),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_243),
.B2(n_244),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_257),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);


endmodule