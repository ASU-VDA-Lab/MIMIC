module fake_jpeg_18376_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_32),
.C(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_15),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_25),
.B1(n_23),
.B2(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_43),
.B1(n_50),
.B2(n_27),
.Y(n_67)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_42),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_18),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_32),
.C(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_31),
.B1(n_28),
.B2(n_20),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_18),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_75),
.Y(n_92)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_51),
.B1(n_24),
.B2(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_72),
.B1(n_0),
.B2(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_69),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_31),
.B1(n_20),
.B2(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_21),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_30),
.C(n_22),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_30),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_32),
.B(n_29),
.C(n_26),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_12),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_9),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_88),
.B(n_93),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_42),
.B1(n_53),
.B2(n_44),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_95),
.B1(n_97),
.B2(n_105),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_101),
.B(n_81),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_32),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_59),
.B1(n_78),
.B2(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_85),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_55),
.B1(n_24),
.B2(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_102),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_79),
.B(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_55),
.B1(n_24),
.B2(n_19),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_83),
.C(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_22),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_10),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_22),
.B1(n_30),
.B2(n_26),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_14),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_73),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_82),
.B1(n_60),
.B2(n_63),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_62),
.B(n_61),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_129),
.B(n_92),
.Y(n_147)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_91),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_71),
.C(n_77),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_70),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_139),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_167)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_93),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_82),
.B1(n_81),
.B2(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_105),
.B1(n_109),
.B2(n_112),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_70),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_140),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_82),
.B1(n_77),
.B2(n_86),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_88),
.B1(n_93),
.B2(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_103),
.B(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_150),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_115),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_92),
.B(n_113),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_129),
.B(n_126),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_124),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_162),
.B1(n_169),
.B2(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_161),
.C(n_122),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_127),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_90),
.C(n_87),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_90),
.B1(n_6),
.B2(n_9),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_26),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_167),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_9),
.B1(n_11),
.B2(n_10),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_192),
.C(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_175),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_170),
.A2(n_121),
.B1(n_118),
.B2(n_116),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_170),
.B1(n_151),
.B2(n_171),
.Y(n_203)
);

XOR2x1_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_117),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_163),
.B(n_155),
.C(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_171),
.B1(n_133),
.B2(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_165),
.B1(n_163),
.B2(n_166),
.Y(n_213)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_183),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_124),
.B(n_130),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_196),
.C(n_169),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_187),
.A2(n_150),
.B1(n_5),
.B2(n_11),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_136),
.C(n_140),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_5),
.C(n_11),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_149),
.C(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_144),
.B(n_5),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_178),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_159),
.C(n_160),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_206),
.C(n_212),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_203),
.Y(n_228)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_188),
.B1(n_168),
.B2(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_161),
.C(n_156),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_192),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_213),
.B1(n_215),
.B2(n_191),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_156),
.C(n_143),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_177),
.B(n_173),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_216),
.B(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_227),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_207),
.A2(n_187),
.B1(n_177),
.B2(n_179),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_193),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_225),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_195),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_174),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_190),
.Y(n_227)
);

AO22x1_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_188),
.B1(n_194),
.B2(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_214),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_213),
.B1(n_211),
.B2(n_215),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_202),
.B1(n_212),
.B2(n_198),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_236),
.B1(n_224),
.B2(n_218),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_210),
.B(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_221),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_198),
.B1(n_204),
.B2(n_4),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_229),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_244),
.B(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_241),
.B(n_242),
.Y(n_259)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_249),
.B(n_250),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_222),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_224),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_219),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_243),
.C(n_241),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_223),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_230),
.C(n_14),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_240),
.C(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_260),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_240),
.C(n_246),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_253),
.CI(n_255),
.CON(n_266),
.SN(n_266)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_266),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_247),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_269),
.B(n_2),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_2),
.C(n_3),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_256),
.A3(n_262),
.B1(n_230),
.B2(n_260),
.C1(n_2),
.C2(n_3),
.Y(n_271)
);

OAI21x1_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_272),
.B(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_266),
.C(n_3),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_270),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_3),
.Y(n_278)
);


endmodule