module real_jpeg_17574_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_2),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_3),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_3),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_4),
.B(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_6),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_6),
.Y(n_117)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_7),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_8),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_8),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_8),
.B(n_151),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_10),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_10),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_10),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_10),
.B(n_54),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_25),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_123),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_121),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_101),
.Y(n_15)
);

NOR2xp67_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_56),
.B2(n_57),
.Y(n_16)
);

INVxp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_38),
.B2(n_39),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

XNOR2x1_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_24),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_22),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_22),
.A2(n_156),
.B1(n_157),
.B2(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_23),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_27)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJx2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.C(n_47),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g137 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_53),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XOR2x1_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_74),
.Y(n_57)
);

XOR2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_66),
.A2(n_73),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_66),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_87),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.C(n_96),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_96),
.B1(n_97),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.C(n_118),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_118),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.C(n_114),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_110),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2x2_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21x1_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_141),
.B(n_182),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_139),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_139),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.C(n_137),
.Y(n_126)
);

XOR2x1_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_130),
.B1(n_137),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_134),
.Y(n_146)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_167),
.Y(n_166)
);

AOI21x1_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_175),
.B(n_181),
.Y(n_141)
);

OAI21x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_158),
.B(n_174),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_155),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_155),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_149),
.C(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_166),
.B(n_173),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);


endmodule