module fake_jpeg_30905_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_34),
.Y(n_45)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_12),
.B(n_3),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_38),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_49),
.B1(n_37),
.B2(n_32),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_46),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_23),
.B1(n_14),
.B2(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_21),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_34),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_71),
.Y(n_87)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_75),
.B1(n_28),
.B2(n_22),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_58),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_25),
.B(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_29),
.B1(n_36),
.B2(n_33),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_0),
.B(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_33),
.C(n_28),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_14),
.B(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_20),
.B1(n_2),
.B2(n_9),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_25),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_86),
.B1(n_73),
.B2(n_69),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_48),
.B1(n_47),
.B2(n_31),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_57),
.B(n_60),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_96),
.B(n_97),
.C(n_98),
.D(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_64),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_63),
.B1(n_68),
.B2(n_20),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_68),
.B(n_20),
.C(n_2),
.D(n_7),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_11),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_101),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_80),
.C(n_78),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

OAI321xp33_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_94),
.A3(n_93),
.B1(n_100),
.B2(n_76),
.C(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_94),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_110),
.C(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_98),
.B1(n_90),
.B2(n_89),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_114),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_118),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_111),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_79),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_123),
.B1(n_119),
.B2(n_77),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_127),
.C(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_128),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_130),
.Y(n_136)
);


endmodule