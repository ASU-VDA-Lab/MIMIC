module fake_jpeg_31420_n_183 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_183);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_30),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_12),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_81),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_24),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_86),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_65),
.B1(n_68),
.B2(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_59),
.B1(n_68),
.B2(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_77),
.B1(n_59),
.B2(n_65),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_77),
.B1(n_53),
.B2(n_74),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_66),
.B1(n_54),
.B2(n_72),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_100),
.B1(n_75),
.B2(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_52),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_72),
.B1(n_75),
.B2(n_70),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_112),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_64),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_69),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_87),
.A3(n_58),
.B1(n_57),
.B2(n_69),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_4),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_26),
.B1(n_51),
.B2(n_46),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_137),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_143),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_145),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_69),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_122),
.A2(n_21),
.B1(n_43),
.B2(n_42),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_7),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_45),
.B1(n_20),
.B2(n_23),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_16),
.B1(n_41),
.B2(n_39),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_1),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_3),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_149),
.B1(n_28),
.B2(n_32),
.Y(n_169)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_161),
.B(n_135),
.C(n_137),
.D(n_34),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_152),
.B1(n_130),
.B2(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_9),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_155),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_9),
.C(n_10),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_158),
.C(n_142),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_13),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_15),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_159),
.Y(n_163)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_33),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_15),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_27),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_133),
.B(n_134),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_167),
.B(n_169),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_166),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_148),
.C(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_160),
.C(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_164),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_162),
.C(n_170),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_163),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_152),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_158),
.B(n_130),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_182),
.B(n_36),
.CI(n_37),
.CON(n_183),
.SN(n_183)
);


endmodule