module real_jpeg_5039_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_1),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_194),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_1),
.A2(n_26),
.B1(n_170),
.B2(n_270),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_92),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_2),
.A2(n_92),
.B1(n_167),
.B2(n_170),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_2),
.A2(n_81),
.B1(n_92),
.B2(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_3),
.Y(n_169)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_5),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_5),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_5),
.B(n_9),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_6),
.A2(n_85),
.B1(n_122),
.B2(n_127),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_6),
.A2(n_45),
.B1(n_85),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_6),
.A2(n_85),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_9),
.A2(n_23),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_9),
.A2(n_52),
.B1(n_160),
.B2(n_164),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_9),
.A2(n_52),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_9),
.A2(n_52),
.B1(n_181),
.B2(n_226),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_9),
.A2(n_136),
.B(n_262),
.C(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_9),
.B(n_57),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_9),
.B(n_296),
.C(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_9),
.B(n_120),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_9),
.B(n_115),
.C(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_9),
.B(n_28),
.Y(n_333)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_11),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_12),
.Y(n_421)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_13),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_415),
.B(n_418),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_409),
.Y(n_15)
);

AO21x2_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_143),
.B(n_408),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_18),
.B(n_140),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_129),
.C(n_138),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_19),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_54),
.C(n_87),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_20),
.A2(n_191),
.B1(n_202),
.B2(n_203),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_20),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_20),
.B(n_150),
.C(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_20),
.B(n_241),
.C(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_20),
.A2(n_202),
.B1(n_241),
.B2(n_334),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_20),
.A2(n_202),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_50),
.B2(n_53),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_21),
.A2(n_27),
.B1(n_50),
.B2(n_53),
.Y(n_228)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_24),
.Y(n_134)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_25),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_27),
.B(n_50),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_27),
.A2(n_53),
.B1(n_130),
.B2(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_27),
.A2(n_50),
.B(n_53),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_27),
.B(n_53),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_40),
.Y(n_27)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_30),
.Y(n_194)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_31),
.Y(n_262)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_33),
.Y(n_264)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_36),
.Y(n_128)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_52),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_53),
.A2(n_130),
.B(n_137),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_54),
.A2(n_87),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_54),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_54),
.B(n_228),
.C(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_54),
.A2(n_383),
.B1(n_385),
.B2(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_83),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_69),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_56),
.A2(n_69),
.B1(n_154),
.B2(n_159),
.Y(n_153)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_56),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_56),
.A2(n_69),
.B1(n_154),
.B2(n_159),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_56),
.A2(n_69),
.B(n_159),
.Y(n_345)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_59),
.Y(n_171)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_59),
.Y(n_175)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_69),
.B(n_159),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_69),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_76),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_83),
.A2(n_207),
.B1(n_209),
.B2(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_86),
.Y(n_208)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_87),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B1(n_120),
.B2(n_121),
.Y(n_87)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_88),
.Y(n_386)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_94),
.Y(n_266)
);

AO22x2_ASAP7_75t_L g191 ( 
.A1(n_95),
.A2(n_120),
.B1(n_192),
.B2(n_197),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_95),
.B(n_192),
.Y(n_387)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_97),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_96),
.A2(n_97),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_112),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_97),
.A2(n_386),
.B(n_387),
.Y(n_385)
);

AOI22x1_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_105),
.B2(n_108),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_114),
.Y(n_316)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_129),
.B(n_138),
.Y(n_405)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_139),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_140),
.B(n_411),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_140),
.B(n_411),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_141),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_403),
.B(n_407),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_374),
.B(n_400),
.Y(n_144)
);

OAI211xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_273),
.B(n_369),
.C(n_373),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_248),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_147),
.A2(n_248),
.B(n_370),
.C(n_372),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_229),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_148),
.B(n_229),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_204),
.C(n_216),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_149),
.B(n_204),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_190),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_165),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_151),
.A2(n_165),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_151),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_151),
.A2(n_258),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_152),
.A2(n_153),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_165),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_172),
.B1(n_179),
.B2(n_186),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_166),
.A2(n_221),
.B(n_224),
.Y(n_220)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_169),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_169),
.Y(n_299)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_172),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_173),
.B(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_173),
.A2(n_225),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_173),
.A2(n_225),
.B1(n_269),
.B2(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_178),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_191),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_191),
.A2(n_203),
.B1(n_218),
.B2(n_219),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_191),
.B(n_218),
.C(n_313),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_191),
.A2(n_203),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_191),
.B(n_254),
.C(n_345),
.Y(n_363)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx6_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_211),
.B2(n_215),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_211),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_209),
.B(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_215),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_211),
.A2(n_235),
.B(n_236),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_212),
.B(n_225),
.Y(n_319)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.C(n_228),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_218),
.A2(n_219),
.B1(n_292),
.B2(n_300),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_218),
.B(n_300),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_228),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_228),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_228),
.A2(n_254),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_228),
.A2(n_254),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_228),
.A2(n_254),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_228),
.B(n_379),
.C(n_384),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_246),
.B2(n_247),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_237),
.B1(n_238),
.B2(n_245),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_237),
.B(n_245),
.C(n_247),
.Y(n_399)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_241),
.B(n_244),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_241),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_241),
.A2(n_330),
.B1(n_331),
.B2(n_334),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_244),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_244),
.A2(n_389),
.B1(n_393),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_249),
.B(n_251),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.C(n_259),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_252),
.B(n_256),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_268),
.C(n_306),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_258),
.B(n_326),
.C(n_328),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_259),
.B(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_260),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_261),
.A2(n_267),
.B1(n_268),
.B2(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_261),
.Y(n_351)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_267),
.A2(n_268),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_287),
.Y(n_288)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_353),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_338),
.B(n_352),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_323),
.B(n_337),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_310),
.B(n_322),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_302),
.B(n_309),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_289),
.B(n_301),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_286),
.B(n_288),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_284),
.A2(n_290),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_290),
.B(n_332),
.C(n_334),
.Y(n_348)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_312),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_321),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_319),
.B2(n_320),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_320),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_336),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_336),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_328),
.B1(n_329),
.B2(n_335),
.Y(n_324)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_340),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_346),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_348),
.C(n_349),
.Y(n_365)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_356),
.B(n_364),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_356),
.C(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.C(n_362),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_360),
.A2(n_362),
.B1(n_363),
.B2(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_360),
.Y(n_368)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_366),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_395),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_375),
.A2(n_401),
.B(n_402),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_388),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_388),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_384),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_385),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_393),
.C(n_394),
.Y(n_388)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_389),
.Y(n_398)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_397),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_399),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_399),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_404),
.B(n_406),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_414),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx13_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_417),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

BUFx12f_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);


endmodule