module fake_jpeg_11410_n_163 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_35),
.Y(n_91)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_37),
.B(n_44),
.Y(n_77)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2x1p5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_3),
.B(n_33),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_12),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_45),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_48),
.Y(n_87)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_17),
.A2(n_19),
.B(n_31),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_25),
.Y(n_53)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_20),
.B(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_26),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_73),
.A3(n_78),
.B1(n_84),
.B2(n_91),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_31),
.B(n_26),
.C(n_22),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_13),
.B1(n_14),
.B2(n_22),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_68),
.B1(n_85),
.B2(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_19),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_61),
.B1(n_57),
.B2(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_92),
.Y(n_102)
);

OAI22x1_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_51),
.B1(n_47),
.B2(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_36),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_34),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_35),
.B(n_30),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_35),
.B(n_3),
.Y(n_86)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_73),
.CON(n_111),
.SN(n_111)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_38),
.A2(n_3),
.B1(n_39),
.B2(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_33),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_78),
.B1(n_79),
.B2(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_103),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_76),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_85),
.C(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_91),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_72),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_85),
.B(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_65),
.B1(n_74),
.B2(n_86),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_112),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_111),
.CON(n_121),
.SN(n_121)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_74),
.B1(n_67),
.B2(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_67),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_97),
.C(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_125),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_70),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_93),
.B(n_102),
.C(n_104),
.D(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_103),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_110),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_134),
.B(n_135),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_104),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_101),
.B1(n_116),
.B2(n_120),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_93),
.B(n_124),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_142),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_128),
.B1(n_136),
.B2(n_135),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_116),
.C(n_127),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_121),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_134),
.B(n_117),
.C(n_120),
.D(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_147),
.Y(n_151)
);

FAx1_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_122),
.CI(n_127),
.CON(n_149),
.SN(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_141),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_144),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_141),
.C(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_146),
.B1(n_123),
.B2(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_146),
.A3(n_102),
.B1(n_95),
.B2(n_100),
.C1(n_113),
.C2(n_88),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_151),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_156),
.C(n_105),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_159),
.C(n_88),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_160),
.Y(n_163)
);


endmodule