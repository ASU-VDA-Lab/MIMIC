module fake_jpeg_25089_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_38),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_29),
.B1(n_23),
.B2(n_25),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_47),
.B1(n_32),
.B2(n_26),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_29),
.B1(n_25),
.B2(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_35),
.B1(n_31),
.B2(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_30),
.B1(n_16),
.B2(n_22),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_38),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_30),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_76),
.B1(n_31),
.B2(n_35),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_75),
.B1(n_17),
.B2(n_20),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_39),
.B1(n_35),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_44),
.B1(n_38),
.B2(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_71),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_39),
.B1(n_33),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_44),
.B1(n_34),
.B2(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_33),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_80),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_27),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_18),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_16),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_82),
.B(n_98),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_52),
.B(n_38),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_85),
.B1(n_73),
.B2(n_59),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_44),
.B1(n_15),
.B2(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_51),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_99),
.B1(n_76),
.B2(n_79),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_20),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_63),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_18),
.A3(n_19),
.B1(n_22),
.B2(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_30),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_106),
.Y(n_140)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_108),
.B1(n_120),
.B2(n_110),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_68),
.B1(n_66),
.B2(n_60),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_118),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_70),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_54),
.B1(n_56),
.B2(n_72),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_76),
.C(n_58),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_37),
.C(n_34),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_72),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_82),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_87),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_61),
.B1(n_57),
.B2(n_55),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_128),
.B1(n_37),
.B2(n_34),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_15),
.B1(n_17),
.B2(n_51),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_122),
.A2(n_85),
.B1(n_83),
.B2(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_51),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_125),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_12),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_19),
.B1(n_22),
.B2(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_143),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_0),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_137),
.B1(n_153),
.B2(n_65),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_86),
.B1(n_94),
.B2(n_103),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_103),
.B(n_2),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_145),
.B(n_37),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_141),
.C(n_123),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_114),
.C(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_37),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_89),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_150),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_92),
.B1(n_65),
.B2(n_19),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_149),
.A2(n_34),
.B1(n_2),
.B2(n_4),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_0),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_156),
.C(n_161),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_128),
.C(n_105),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_145),
.B(n_148),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_164),
.B1(n_130),
.B2(n_136),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_34),
.C(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_0),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

BUFx12f_ASAP7_75t_SL g163 ( 
.A(n_145),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_129),
.B1(n_138),
.B2(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_11),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_2),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_132),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_170),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_137),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_5),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_11),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_134),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_150),
.C(n_139),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_149),
.B1(n_157),
.B2(n_145),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_163),
.B(n_148),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_167),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_156),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_155),
.Y(n_195)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_188),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_191),
.A2(n_193),
.B(n_194),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_176),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_144),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_171),
.B(n_158),
.Y(n_198)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_201),
.B1(n_183),
.B2(n_184),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_164),
.B1(n_161),
.B2(n_133),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_190),
.B1(n_201),
.B2(n_194),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_174),
.C(n_178),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_206),
.C(n_207),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_178),
.C(n_175),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_175),
.C(n_186),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_166),
.C(n_173),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_146),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_199),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_190),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_198),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_210),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_204),
.C(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_222),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_159),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_217),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_220),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_224),
.A3(n_159),
.B1(n_209),
.B2(n_219),
.C1(n_207),
.C2(n_5),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_228),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_230),
.A2(n_6),
.B(n_7),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_SL g233 ( 
.A(n_231),
.B(n_7),
.C(n_8),
.Y(n_233)
);

AOI31xp33_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_233),
.A3(n_9),
.B(n_10),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_229),
.C(n_9),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_10),
.Y(n_236)
);


endmodule