module fake_ibex_1472_n_1202 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1202);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1202;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_1148;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_1196;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_1182;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_972;
wire n_947;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_1199;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1152;
wire n_1034;
wire n_371;
wire n_1036;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_457;
wire n_412;
wire n_357;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1044;
wire n_1106;
wire n_1018;
wire n_1129;
wire n_449;
wire n_1138;
wire n_547;
wire n_1131;
wire n_727;
wire n_1134;
wire n_1077;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_1174;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_1189;
wire n_531;
wire n_647;
wire n_1187;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_375;
wire n_280;
wire n_340;
wire n_317;
wire n_698;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1166;
wire n_1181;
wire n_1140;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_1193;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1172;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_1169;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_1201;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1177;
wire n_1068;
wire n_1057;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_1184;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_1195;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1136;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_1075;
wire n_574;
wire n_1168;
wire n_1197;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_1179;
wire n_1192;
wire n_933;
wire n_1081;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1191;
wire n_1101;
wire n_518;
wire n_367;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_1178;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_1082;
wire n_1137;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1200;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_968;
wire n_625;
wire n_1180;
wire n_953;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_1171;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_1183;
wire n_253;
wire n_234;
wire n_300;
wire n_1151;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1038;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_472;
wire n_229;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1173;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1126;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_1170;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_1158;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_1176;
wire n_940;
wire n_444;
wire n_562;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_1160;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_1198;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_1167;
wire n_653;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_1190;
wire n_517;
wire n_744;
wire n_817;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_285;
wire n_247;
wire n_379;
wire n_288;
wire n_1128;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_820;
wire n_805;
wire n_670;
wire n_728;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_1175;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1102;
wire n_1005;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_1150;
wire n_462;
wire n_1194;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_1185;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_890;
wire n_921;
wire n_874;
wire n_912;
wire n_1058;
wire n_1105;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_1000;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_1186;
wire n_657;
wire n_764;
wire n_1156;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_58),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_141),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_155),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_71),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_41),
.Y(n_228)
);

INVx4_ASAP7_75t_R g229 ( 
.A(n_82),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_75),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_196),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_1),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_107),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_21),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_148),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_109),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_90),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_116),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_L g245 ( 
.A(n_3),
.B(n_168),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

CKINVDCx6p67_ASAP7_75t_R g247 ( 
.A(n_158),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_137),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_67),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_103),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_134),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_39),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_145),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_14),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_132),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_133),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_15),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_12),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_26),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_156),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_125),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_30),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_19),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_197),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_184),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g273 ( 
.A(n_33),
.B(n_13),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_152),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_73),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_106),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_150),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_147),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_95),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_0),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_58),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_18),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_42),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_92),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_13),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_179),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_64),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_138),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_77),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_93),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_101),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_52),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_10),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_127),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_33),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_129),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_38),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_70),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_182),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_102),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_175),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_164),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_188),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_185),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_68),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_17),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_60),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_57),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_208),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_169),
.Y(n_312)
);

BUFx8_ASAP7_75t_SL g313 ( 
.A(n_217),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_130),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_211),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_209),
.B(n_65),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_23),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_59),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_195),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_49),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_104),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_83),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_146),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_118),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_22),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_28),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_157),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_149),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_105),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_84),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_113),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_94),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_100),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_1),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_215),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_44),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_39),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_37),
.B(n_36),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_57),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_216),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_203),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_79),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_210),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_51),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_97),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_22),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_32),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_122),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_207),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_212),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_80),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_165),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_167),
.Y(n_354)
);

BUFx2_ASAP7_75t_SL g355 ( 
.A(n_47),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_206),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_191),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_112),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_142),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_24),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_151),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_74),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_99),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_205),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_50),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_201),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_63),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_10),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_87),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_143),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_32),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_144),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_91),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_110),
.Y(n_374)
);

BUFx8_ASAP7_75t_SL g375 ( 
.A(n_257),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_234),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_253),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_253),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_238),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_243),
.A2(n_66),
.B(n_62),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_234),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_283),
.B(n_2),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_253),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_283),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_253),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_236),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_253),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_310),
.B(n_2),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_253),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_253),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_223),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_270),
.B(n_3),
.Y(n_394)
);

OAI22x1_ASAP7_75t_R g395 ( 
.A1(n_257),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_270),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_281),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_281),
.Y(n_398)
);

BUFx8_ASAP7_75t_SL g399 ( 
.A(n_265),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_265),
.B(n_294),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_313),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_243),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_340),
.B(n_244),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_267),
.Y(n_405)
);

INVx6_ASAP7_75t_L g406 ( 
.A(n_234),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_237),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_294),
.B(n_5),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_237),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_244),
.B(n_6),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_269),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_237),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_271),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_338),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_256),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_225),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_255),
.B(n_7),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_267),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_228),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_230),
.Y(n_422)
);

BUFx8_ASAP7_75t_SL g423 ( 
.A(n_360),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_235),
.B(n_9),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_315),
.A2(n_328),
.B(n_322),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_254),
.B(n_12),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_315),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_262),
.B(n_14),
.Y(n_428)
);

AOI22x1_ASAP7_75t_SL g429 ( 
.A1(n_360),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_328),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_332),
.B(n_16),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_228),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_352),
.A2(n_119),
.B(n_220),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_352),
.A2(n_366),
.B(n_232),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_286),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_231),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_228),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_228),
.Y(n_438)
);

INVx6_ASAP7_75t_L g439 ( 
.A(n_237),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_374),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_256),
.Y(n_441)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_333),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_366),
.A2(n_120),
.B(n_219),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_255),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_246),
.A2(n_117),
.B(n_218),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_282),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_249),
.A2(n_121),
.B(n_213),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_333),
.Y(n_448)
);

OAI22x1_ASAP7_75t_R g449 ( 
.A1(n_260),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_449)
);

BUFx12f_ASAP7_75t_L g450 ( 
.A(n_286),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_333),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_332),
.B(n_27),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_250),
.B(n_28),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_251),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_252),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_333),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_296),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_296),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_457),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_412),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_457),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_410),
.B(n_355),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_457),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_417),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_419),
.B(n_304),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_419),
.B(n_259),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_382),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_387),
.B(n_241),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_383),
.A2(n_284),
.B1(n_295),
.B2(n_287),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_401),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_387),
.B(n_264),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_419),
.B(n_261),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_458),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_401),
.B(n_346),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_378),
.B(n_273),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_419),
.B(n_263),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_418),
.B(n_266),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_412),
.B(n_224),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_425),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_378),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g492 ( 
.A(n_431),
.B(n_260),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_403),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_378),
.B(n_389),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_418),
.B(n_275),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

NOR2x1p5_ASAP7_75t_L g497 ( 
.A(n_450),
.B(n_247),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_425),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_404),
.B(n_286),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_422),
.B(n_276),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_431),
.A2(n_308),
.B1(n_309),
.B2(n_299),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_377),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_389),
.B(n_319),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_377),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_404),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_379),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_389),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_379),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_384),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_384),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_452),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_386),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_422),
.B(n_326),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_441),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_388),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_436),
.B(n_335),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_436),
.B(n_279),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_375),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_391),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_444),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_391),
.Y(n_528)
);

INVx8_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_454),
.B(n_289),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_454),
.B(n_455),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_392),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_392),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_427),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_444),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_399),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_435),
.B(n_373),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_434),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_455),
.B(n_290),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_415),
.B(n_291),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_434),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_411),
.B(n_300),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_411),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_406),
.Y(n_547)
);

AND3x2_ASAP7_75t_L g548 ( 
.A(n_402),
.B(n_305),
.C(n_318),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_SL g549 ( 
.A(n_390),
.B(n_277),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_393),
.B(n_307),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_380),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_396),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_413),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_390),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_411),
.B(n_311),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_396),
.B(n_227),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_400),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_376),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_411),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_397),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_397),
.Y(n_562)
);

AND2x2_ASAP7_75t_SL g563 ( 
.A(n_381),
.B(n_312),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_398),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_406),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_411),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_398),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_423),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_433),
.B(n_323),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_408),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_408),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_424),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_426),
.B(n_324),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_421),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_381),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_453),
.B(n_325),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_428),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_381),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_421),
.B(n_330),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_421),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_421),
.B(n_233),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_432),
.Y(n_582)
);

NOR2x1p5_ASAP7_75t_L g583 ( 
.A(n_400),
.B(n_409),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_SL g584 ( 
.A(n_440),
.B(n_278),
.C(n_277),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_432),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_446),
.A2(n_342),
.B(n_341),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_577),
.B(n_381),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_529),
.B(n_416),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_553),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_513),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_460),
.B(n_443),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_554),
.B(n_327),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_517),
.B(n_443),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_570),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_529),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_443),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_473),
.B(n_443),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_473),
.B(n_343),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_513),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_490),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_570),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_475),
.B(n_344),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_461),
.B(n_356),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_479),
.B(n_239),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_476),
.A2(n_440),
.B1(n_292),
.B2(n_278),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_468),
.A2(n_345),
.B1(n_347),
.B2(n_365),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_498),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_478),
.B(n_240),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_466),
.B(n_359),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_468),
.A2(n_337),
.B1(n_368),
.B2(n_371),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_536),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_508),
.A2(n_292),
.B1(n_374),
.B2(n_320),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_468),
.A2(n_348),
.B1(n_320),
.B2(n_327),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_551),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_529),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_477),
.B(n_242),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_467),
.B(n_361),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_584),
.B(n_437),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_536),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_500),
.B(n_248),
.Y(n_620)
);

BUFx5_ASAP7_75t_L g621 ( 
.A(n_468),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_469),
.B(n_362),
.Y(n_623)
);

INVx8_ASAP7_75t_L g624 ( 
.A(n_463),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_472),
.B(n_268),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_539),
.B(n_272),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_463),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_463),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_519),
.B(n_523),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_554),
.B(n_409),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_490),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_482),
.B(n_274),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_487),
.B(n_280),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_586),
.A2(n_327),
.B1(n_364),
.B2(n_370),
.Y(n_635)
);

O2A1O1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_531),
.A2(n_258),
.B(n_297),
.C(n_369),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_483),
.B(n_285),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_492),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_531),
.B(n_573),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_508),
.B(n_288),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

OAI221xp5_ASAP7_75t_L g642 ( 
.A1(n_504),
.A2(n_339),
.B1(n_245),
.B2(n_293),
.C(n_298),
.Y(n_642)
);

BUFx6f_ASAP7_75t_SL g643 ( 
.A(n_483),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_562),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_540),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_483),
.B(n_301),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_558),
.A2(n_395),
.B1(n_429),
.B2(n_449),
.Y(n_647)
);

OAI221xp5_ASAP7_75t_L g648 ( 
.A1(n_550),
.A2(n_357),
.B1(n_302),
.B2(n_303),
.C(n_306),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_489),
.A2(n_438),
.B(n_437),
.C(n_367),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_494),
.B(n_445),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_535),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_543),
.B(n_445),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_497),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_548),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_496),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_506),
.B(n_226),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_492),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_545),
.Y(n_659)
);

BUFx6f_ASAP7_75t_SL g660 ( 
.A(n_568),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_564),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_465),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_567),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_470),
.B(n_447),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_549),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_491),
.B(n_317),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_470),
.B(n_447),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_480),
.B(n_447),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_574),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_571),
.A2(n_449),
.B1(n_395),
.B2(n_314),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_510),
.B(n_316),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_542),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_480),
.B(n_329),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_489),
.A2(n_429),
.B1(n_331),
.B2(n_334),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_493),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_503),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_511),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_514),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_485),
.B(n_336),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_521),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_556),
.B(n_349),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_485),
.B(n_350),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_496),
.B(n_353),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_532),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_486),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_586),
.A2(n_438),
.B1(n_437),
.B2(n_358),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_581),
.B(n_354),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_576),
.B(n_363),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_538),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_499),
.B(n_372),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_501),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_520),
.B(n_438),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_501),
.Y(n_693)
);

O2A1O1Ixp5_ASAP7_75t_L g694 ( 
.A1(n_569),
.A2(n_229),
.B(n_439),
.C(n_442),
.Y(n_694)
);

NOR3xp33_ASAP7_75t_L g695 ( 
.A(n_525),
.B(n_29),
.C(n_30),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_545),
.B(n_495),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_537),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_495),
.B(n_439),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_502),
.B(n_439),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_524),
.A2(n_442),
.B1(n_439),
.B2(n_448),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_547),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_530),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_530),
.B(n_442),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_547),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_541),
.B(n_407),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_558),
.B(n_72),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_563),
.B(n_407),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_579),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_505),
.B(n_507),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_563),
.A2(n_456),
.B1(n_451),
.B2(n_448),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_579),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_507),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_509),
.B(n_407),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_509),
.B(n_31),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_544),
.B(n_76),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_575),
.A2(n_526),
.B(n_512),
.C(n_534),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_589),
.B(n_515),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_691),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_587),
.A2(n_555),
.B(n_516),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_629),
.B(n_515),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_672),
.B(n_555),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_595),
.B(n_518),
.Y(n_723)
);

AO32x2_ASAP7_75t_L g724 ( 
.A1(n_670),
.A2(n_605),
.A3(n_659),
.B1(n_702),
.B2(n_685),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_664),
.A2(n_668),
.B(n_667),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_612),
.B(n_522),
.Y(n_726)
);

NAND2x2_ASAP7_75t_L g727 ( 
.A(n_628),
.B(n_546),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_693),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_596),
.A2(n_533),
.B(n_528),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_600),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_676),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_645),
.A2(n_585),
.B1(n_582),
.B2(n_580),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_613),
.A2(n_560),
.B1(n_566),
.B2(n_462),
.Y(n_733)
);

OA21x2_ASAP7_75t_L g734 ( 
.A1(n_652),
.A2(n_462),
.B(n_459),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_639),
.B(n_676),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_639),
.B(n_560),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_662),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_624),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_606),
.A2(n_481),
.B1(n_488),
.B2(n_484),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_615),
.B(n_557),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_621),
.B(n_464),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_630),
.B(n_31),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_674),
.B(n_34),
.Y(n_743)
);

BUFx4f_ASAP7_75t_L g744 ( 
.A(n_624),
.Y(n_744)
);

OAI21xp33_ASAP7_75t_L g745 ( 
.A1(n_592),
.A2(n_474),
.B(n_565),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_611),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_650),
.A2(n_696),
.B(n_707),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_627),
.B(n_35),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_635),
.B(n_414),
.C(n_448),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_619),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_624),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_600),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_605),
.B(n_35),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_640),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_614),
.B(n_40),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_634),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_638),
.A2(n_665),
.B1(n_588),
.B2(n_715),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_675),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_683),
.A2(n_690),
.B(n_593),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_641),
.B(n_40),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_644),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_661),
.B(n_41),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_590),
.Y(n_763)
);

OR2x4_ASAP7_75t_L g764 ( 
.A(n_706),
.B(n_43),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_663),
.B(n_43),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_610),
.A2(n_414),
.B1(n_448),
.B2(n_451),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_692),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_R g768 ( 
.A(n_697),
.B(n_45),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_591),
.A2(n_414),
.B(n_451),
.C(n_448),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_677),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_667),
.A2(n_668),
.B(n_717),
.Y(n_771)
);

CKINVDCx8_ASAP7_75t_R g772 ( 
.A(n_588),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_SL g773 ( 
.A(n_621),
.B(n_559),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_709),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_588),
.A2(n_456),
.B1(n_47),
.B2(n_48),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_656),
.B(n_46),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_678),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_680),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_653),
.B(n_52),
.Y(n_779)
);

CKINVDCx6p67_ASAP7_75t_R g780 ( 
.A(n_660),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_654),
.B(n_53),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_689),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_620),
.B(n_53),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_594),
.Y(n_784)
);

NOR2x1p5_ASAP7_75t_SL g785 ( 
.A(n_621),
.B(n_78),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_684),
.B(n_604),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_713),
.B(n_54),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_686),
.B(n_471),
.C(n_56),
.Y(n_788)
);

AO21x1_ASAP7_75t_L g789 ( 
.A1(n_649),
.A2(n_55),
.B(n_56),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_L g790 ( 
.A(n_712),
.B(n_55),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_637),
.B(n_60),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_601),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_616),
.B(n_61),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_633),
.B(n_222),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_647),
.B(n_81),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_631),
.Y(n_796)
);

OAI21xp33_ASAP7_75t_L g797 ( 
.A1(n_598),
.A2(n_85),
.B(n_86),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_599),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_598),
.A2(n_88),
.B(n_89),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_710),
.A2(n_96),
.B(n_98),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_694),
.A2(n_108),
.B(n_111),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_646),
.B(n_114),
.Y(n_802)
);

OR2x6_ASAP7_75t_SL g803 ( 
.A(n_660),
.B(n_123),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_643),
.B(n_126),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_636),
.A2(n_128),
.B(n_131),
.C(n_135),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_602),
.A2(n_136),
.B(n_139),
.C(n_140),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_643),
.B(n_154),
.Y(n_807)
);

AOI21x1_ASAP7_75t_L g808 ( 
.A1(n_705),
.A2(n_159),
.B(n_160),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_603),
.A2(n_161),
.B(n_162),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_648),
.B(n_163),
.Y(n_810)
);

CKINVDCx10_ASAP7_75t_R g811 ( 
.A(n_695),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_609),
.A2(n_166),
.B(n_170),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_642),
.B(n_172),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_607),
.Y(n_814)
);

AOI21x1_ASAP7_75t_L g815 ( 
.A1(n_705),
.A2(n_173),
.B(n_174),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_SL g816 ( 
.A1(n_714),
.A2(n_180),
.B(n_186),
.C(n_187),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_617),
.A2(n_189),
.B(n_193),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_623),
.A2(n_198),
.B(n_199),
.C(n_202),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_655),
.A2(n_679),
.B(n_673),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_626),
.B(n_688),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_744),
.B(n_651),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_759),
.A2(n_625),
.B(n_632),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_737),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_774),
.B(n_618),
.Y(n_824)
);

AND2x6_ASAP7_75t_L g825 ( 
.A(n_774),
.B(n_708),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_721),
.B(n_666),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_813),
.B(n_622),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_747),
.A2(n_681),
.B(n_687),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_757),
.A2(n_711),
.B1(n_666),
.B2(n_682),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_735),
.A2(n_657),
.B1(n_669),
.B2(n_671),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_718),
.B(n_753),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_726),
.B(n_608),
.Y(n_832)
);

AO21x1_ASAP7_75t_L g833 ( 
.A1(n_817),
.A2(n_716),
.B(n_703),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_771),
.A2(n_699),
.B(n_698),
.Y(n_834)
);

NOR2x1_ASAP7_75t_L g835 ( 
.A(n_788),
.B(n_701),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_772),
.B(n_704),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_748),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_744),
.B(n_700),
.Y(n_838)
);

BUFx4f_ASAP7_75t_SL g839 ( 
.A(n_780),
.Y(n_839)
);

AO32x2_ASAP7_75t_L g840 ( 
.A1(n_775),
.A2(n_733),
.A3(n_739),
.B1(n_766),
.B2(n_767),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_754),
.B(n_742),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_751),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_756),
.B(n_761),
.Y(n_843)
);

AO31x2_ASAP7_75t_L g844 ( 
.A1(n_769),
.A2(n_789),
.A3(n_805),
.B(n_806),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_782),
.B(n_820),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_748),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_719),
.A2(n_728),
.B1(n_787),
.B2(n_777),
.Y(n_847)
);

NOR2x1_ASAP7_75t_SL g848 ( 
.A(n_802),
.B(n_731),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_736),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_729),
.A2(n_819),
.B(n_720),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_768),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_724),
.B(n_803),
.Y(n_852)
);

AO22x2_ASAP7_75t_L g853 ( 
.A1(n_724),
.A2(n_795),
.B1(n_788),
.B2(n_776),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_802),
.B(n_743),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_R g855 ( 
.A(n_811),
.B(n_804),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_R g856 ( 
.A(n_807),
.B(n_722),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_781),
.B(n_758),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_770),
.B(n_778),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_793),
.B(n_783),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_784),
.B(n_792),
.Y(n_860)
);

OAI22x1_ASAP7_75t_L g861 ( 
.A1(n_791),
.A2(n_810),
.B1(n_764),
.B2(n_802),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_790),
.B(n_779),
.Y(n_862)
);

AOI221x1_ASAP7_75t_L g863 ( 
.A1(n_801),
.A2(n_797),
.B1(n_800),
.B2(n_817),
.C(n_749),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_755),
.A2(n_760),
.B(n_762),
.C(n_765),
.Y(n_864)
);

NAND2x1_ASAP7_75t_L g865 ( 
.A(n_746),
.B(n_750),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_764),
.Y(n_866)
);

AOI21xp33_ASAP7_75t_L g867 ( 
.A1(n_745),
.A2(n_794),
.B(n_732),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_800),
.A2(n_818),
.B(n_809),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_814),
.B(n_763),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_763),
.B(n_798),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_723),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_798),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_734),
.A2(n_815),
.B(n_808),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_785),
.A2(n_799),
.B(n_773),
.C(n_812),
.Y(n_874)
);

HAxp5_ASAP7_75t_L g875 ( 
.A(n_727),
.B(n_740),
.CON(n_875),
.SN(n_875)
);

AO31x2_ASAP7_75t_L g876 ( 
.A1(n_741),
.A2(n_816),
.A3(n_752),
.B(n_796),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_796),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_774),
.B(n_738),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_737),
.B(n_630),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_774),
.B(n_460),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_774),
.B(n_460),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_718),
.B(n_554),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_774),
.B(n_460),
.Y(n_885)
);

AOI21xp33_ASAP7_75t_L g886 ( 
.A1(n_754),
.A2(n_672),
.B(n_508),
.Y(n_886)
);

AO31x2_ASAP7_75t_L g887 ( 
.A1(n_769),
.A2(n_759),
.A3(n_717),
.B(n_789),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_759),
.A2(n_725),
.B(n_747),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_780),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_774),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_780),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_774),
.B(n_460),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_744),
.B(n_751),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_774),
.A2(n_549),
.B1(n_492),
.B2(n_441),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_774),
.Y(n_897)
);

NOR2xp67_ASAP7_75t_L g898 ( 
.A(n_721),
.B(n_813),
.Y(n_898)
);

AOI221x1_ASAP7_75t_L g899 ( 
.A1(n_788),
.A2(n_759),
.B1(n_769),
.B2(n_801),
.C(n_797),
.Y(n_899)
);

OA22x2_ASAP7_75t_L g900 ( 
.A1(n_737),
.A2(n_400),
.B1(n_612),
.B2(n_647),
.Y(n_900)
);

AOI221x1_ASAP7_75t_L g901 ( 
.A1(n_788),
.A2(n_759),
.B1(n_769),
.B2(n_801),
.C(n_797),
.Y(n_901)
);

AO32x2_ASAP7_75t_L g902 ( 
.A1(n_775),
.A2(n_578),
.A3(n_733),
.B1(n_739),
.B2(n_766),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_774),
.B(n_460),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_718),
.B(n_554),
.Y(n_904)
);

AND3x4_ASAP7_75t_L g905 ( 
.A(n_743),
.B(n_695),
.C(n_628),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_737),
.B(n_630),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_730),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_737),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_774),
.A2(n_721),
.B1(n_529),
.B2(n_517),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_774),
.B(n_460),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_774),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_L g912 ( 
.A(n_805),
.B(n_788),
.C(n_754),
.Y(n_912)
);

OAI21x1_ASAP7_75t_SL g913 ( 
.A1(n_817),
.A2(n_800),
.B(n_735),
.Y(n_913)
);

AO31x2_ASAP7_75t_L g914 ( 
.A1(n_769),
.A2(n_759),
.A3(n_717),
.B(n_789),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_737),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_817),
.A2(n_759),
.B(n_800),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_737),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_730),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_774),
.B(n_460),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_774),
.B(n_460),
.Y(n_920)
);

INVx5_ASAP7_75t_L g921 ( 
.A(n_751),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_774),
.Y(n_922)
);

OAI21xp33_ASAP7_75t_L g923 ( 
.A1(n_786),
.A2(n_672),
.B(n_554),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_924)
);

AO31x2_ASAP7_75t_L g925 ( 
.A1(n_769),
.A2(n_759),
.A3(n_717),
.B(n_789),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_774),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_718),
.B(n_554),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_805),
.B(n_788),
.C(n_754),
.Y(n_929)
);

BUFx6f_ASAP7_75t_SL g930 ( 
.A(n_748),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_718),
.B(n_554),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_759),
.A2(n_597),
.B(n_587),
.Y(n_933)
);

AOI221xp5_ASAP7_75t_SL g934 ( 
.A1(n_754),
.A2(n_642),
.B1(n_636),
.B2(n_635),
.C(n_658),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_780),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_880),
.B(n_906),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_908),
.B(n_915),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_917),
.B(n_823),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_892),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_831),
.B(n_884),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_849),
.B(n_898),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_843),
.Y(n_942)
);

INVx8_ASAP7_75t_L g943 ( 
.A(n_921),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_930),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_904),
.B(n_927),
.Y(n_945)
);

OA21x2_ASAP7_75t_L g946 ( 
.A1(n_899),
.A2(n_901),
.B(n_873),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_932),
.B(n_841),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_900),
.A2(n_852),
.B1(n_854),
.B2(n_861),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_839),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_835),
.A2(n_916),
.B(n_868),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_921),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_921),
.B(n_878),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_886),
.B(n_923),
.Y(n_954)
);

CKINVDCx16_ASAP7_75t_R g955 ( 
.A(n_851),
.Y(n_955)
);

NAND3xp33_ASAP7_75t_SL g956 ( 
.A(n_905),
.B(n_856),
.C(n_895),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_894),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_890),
.Y(n_958)
);

OAI22xp33_ASAP7_75t_L g959 ( 
.A1(n_854),
.A2(n_846),
.B1(n_881),
.B2(n_910),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_821),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_845),
.B(n_922),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_926),
.B(n_848),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_879),
.A2(n_888),
.B(n_928),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_833),
.A2(n_863),
.A3(n_874),
.B(n_850),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_926),
.A2(n_919),
.B1(n_882),
.B2(n_903),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_SL g966 ( 
.A1(n_837),
.A2(n_909),
.B(n_866),
.Y(n_966)
);

CKINVDCx14_ASAP7_75t_R g967 ( 
.A(n_935),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_858),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_838),
.B(n_857),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_869),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_883),
.A2(n_896),
.B(n_924),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_931),
.A2(n_933),
.B(n_889),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_842),
.B(n_885),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_930),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_893),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_827),
.A2(n_934),
.B1(n_826),
.B2(n_859),
.Y(n_976)
);

AO21x2_ASAP7_75t_L g977 ( 
.A1(n_912),
.A2(n_929),
.B(n_864),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_834),
.A2(n_822),
.B(n_835),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_872),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_920),
.A2(n_832),
.B1(n_829),
.B2(n_853),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_824),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_853),
.A2(n_847),
.B1(n_867),
.B2(n_870),
.Y(n_982)
);

AOI221xp5_ASAP7_75t_L g983 ( 
.A1(n_836),
.A2(n_830),
.B1(n_828),
.B2(n_855),
.C(n_871),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_825),
.B(n_925),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_862),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_865),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_887),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_887),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_887),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_877),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_875),
.B(n_907),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_914),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_907),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_918),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_914),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_925),
.B(n_840),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_902),
.A2(n_876),
.B(n_840),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_918),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_925),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_844),
.Y(n_1000)
);

NAND2x1p5_ASAP7_75t_L g1001 ( 
.A(n_891),
.B(n_744),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_SL g1002 ( 
.A1(n_898),
.A2(n_852),
.B(n_817),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_839),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_908),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_891),
.B(n_744),
.Y(n_1005)
);

BUFx12f_ASAP7_75t_L g1006 ( 
.A(n_890),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_839),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_R g1008 ( 
.A(n_890),
.B(n_568),
.Y(n_1008)
);

NAND2x1p5_ASAP7_75t_L g1009 ( 
.A(n_891),
.B(n_744),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_831),
.B(n_884),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_854),
.A2(n_849),
.B1(n_911),
.B2(n_897),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_923),
.B(n_670),
.C(n_647),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_891),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_SL g1014 ( 
.A1(n_848),
.A2(n_817),
.B(n_913),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_908),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_892),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_839),
.Y(n_1017)
);

INVxp33_ASAP7_75t_SL g1018 ( 
.A(n_890),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_899),
.A2(n_901),
.B(n_873),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_1012),
.A2(n_956),
.B1(n_954),
.B2(n_969),
.Y(n_1020)
);

AO21x2_ASAP7_75t_L g1021 ( 
.A1(n_963),
.A2(n_971),
.B(n_978),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_996),
.B(n_987),
.Y(n_1022)
);

INVxp33_ASAP7_75t_L g1023 ( 
.A(n_1008),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_988),
.B(n_989),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_992),
.B(n_995),
.Y(n_1025)
);

CKINVDCx14_ASAP7_75t_R g1026 ( 
.A(n_1016),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_943),
.Y(n_1027)
);

AO21x2_ASAP7_75t_L g1028 ( 
.A1(n_978),
.A2(n_972),
.B(n_951),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_993),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_941),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_998),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_998),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_961),
.B(n_942),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_998),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_969),
.A2(n_1011),
.B1(n_947),
.B2(n_949),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_977),
.B(n_948),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_994),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_940),
.B(n_1010),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_972),
.A2(n_1014),
.B(n_1019),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_SL g1040 ( 
.A(n_1011),
.B(n_965),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_959),
.A2(n_936),
.B1(n_983),
.B2(n_985),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_965),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_997),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_980),
.B(n_1000),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_980),
.B(n_999),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_968),
.Y(n_1046)
);

INVx5_ASAP7_75t_SL g1047 ( 
.A(n_962),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_943),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_984),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_986),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_970),
.B(n_975),
.Y(n_1051)
);

OAI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_976),
.A2(n_966),
.B1(n_945),
.B2(n_973),
.C(n_1004),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1024),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1022),
.B(n_964),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1022),
.B(n_964),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1043),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_1042),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1022),
.B(n_964),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1025),
.B(n_946),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1025),
.B(n_982),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1031),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1025),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1036),
.B(n_1002),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_1042),
.B(n_937),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1033),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_1049),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1045),
.B(n_938),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1036),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1021),
.B(n_981),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1045),
.B(n_1013),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1050),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_1049),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_1026),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_1029),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1054),
.B(n_1044),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1053),
.B(n_1045),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1054),
.B(n_1028),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1074),
.B(n_1023),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1059),
.B(n_1039),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1070),
.A2(n_1052),
.B1(n_1020),
.B2(n_1035),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1055),
.B(n_1028),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_1065),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1056),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1061),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_1064),
.B(n_1028),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_1073),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_1072),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1071),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1055),
.B(n_1028),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1071),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1055),
.B(n_1040),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1072),
.Y(n_1092)
);

AOI222xp33_ASAP7_75t_L g1093 ( 
.A1(n_1060),
.A2(n_1041),
.B1(n_1038),
.B2(n_1052),
.C1(n_1046),
.C2(n_1030),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1062),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1077),
.B(n_1058),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1082),
.B(n_1058),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1094),
.B(n_1058),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1077),
.B(n_1063),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1094),
.B(n_1069),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_1085),
.B(n_1068),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1093),
.A2(n_1061),
.B(n_1038),
.Y(n_1101)
);

NAND2x1_ASAP7_75t_L g1102 ( 
.A(n_1087),
.B(n_1066),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1083),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_1084),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1088),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1088),
.Y(n_1106)
);

AO22x1_ASAP7_75t_L g1107 ( 
.A1(n_1087),
.A2(n_1066),
.B1(n_1057),
.B2(n_1027),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_1092),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1081),
.B(n_1063),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1081),
.B(n_1063),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1105),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1105),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1095),
.B(n_1089),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1106),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1103),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1106),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1096),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1100),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1098),
.B(n_1079),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1101),
.A2(n_1080),
.B1(n_1102),
.B2(n_1108),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1104),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1100),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1097),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1103),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_1104),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1102),
.A2(n_1092),
.B1(n_1047),
.B2(n_1067),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1117),
.B(n_1123),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1115),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1119),
.B(n_1098),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1112),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1118),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1113),
.B(n_1109),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1120),
.A2(n_1086),
.B(n_1078),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1122),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1121),
.A2(n_1093),
.B(n_1048),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1125),
.B(n_1109),
.Y(n_1136)
);

AOI32xp33_ASAP7_75t_L g1137 ( 
.A1(n_1119),
.A2(n_1108),
.A3(n_1110),
.B1(n_1095),
.B2(n_1091),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1112),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1126),
.A2(n_1091),
.B1(n_1110),
.B2(n_1089),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1114),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1114),
.Y(n_1141)
);

OAI211xp5_ASAP7_75t_L g1142 ( 
.A1(n_1116),
.A2(n_1029),
.B(n_1037),
.C(n_943),
.Y(n_1142)
);

AOI32xp33_ASAP7_75t_L g1143 ( 
.A1(n_1129),
.A2(n_1108),
.A3(n_1037),
.B1(n_1027),
.B2(n_1060),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1129),
.B(n_1079),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1138),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1133),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1128),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1128),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1135),
.A2(n_1107),
.B(n_1040),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1127),
.B(n_939),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1131),
.B(n_1134),
.Y(n_1151)
);

OAI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1146),
.A2(n_1137),
.B1(n_1142),
.B2(n_1139),
.C(n_1136),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1150),
.B(n_1008),
.C(n_955),
.Y(n_1153)
);

AOI222xp33_ASAP7_75t_L g1154 ( 
.A1(n_1151),
.A2(n_1130),
.B1(n_1140),
.B2(n_1141),
.C1(n_1111),
.C2(n_1116),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1151),
.B(n_1132),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1145),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1147),
.B(n_1132),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1143),
.B(n_1130),
.Y(n_1158)
);

OAI221xp5_ASAP7_75t_L g1159 ( 
.A1(n_1149),
.A2(n_1076),
.B1(n_966),
.B2(n_944),
.C(n_1067),
.Y(n_1159)
);

OAI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1144),
.A2(n_1099),
.B1(n_1076),
.B2(n_1085),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1148),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1154),
.B(n_1115),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_1153),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_1158),
.Y(n_1164)
);

AOI211xp5_ASAP7_75t_L g1165 ( 
.A1(n_1152),
.A2(n_1017),
.B(n_1007),
.C(n_1003),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1155),
.B(n_1124),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1156),
.B(n_1124),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1159),
.B(n_991),
.C(n_974),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1160),
.B(n_1090),
.Y(n_1169)
);

NOR4xp25_ASAP7_75t_L g1170 ( 
.A(n_1163),
.B(n_1161),
.C(n_1157),
.D(n_979),
.Y(n_1170)
);

NOR2x1_ASAP7_75t_L g1171 ( 
.A(n_1168),
.B(n_1027),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_L g1172 ( 
.A(n_1165),
.B(n_1164),
.C(n_1162),
.Y(n_1172)
);

AND4x1_ASAP7_75t_L g1173 ( 
.A(n_1169),
.B(n_1018),
.C(n_967),
.D(n_1006),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_L g1174 ( 
.A(n_1167),
.B(n_950),
.C(n_958),
.Y(n_1174)
);

NAND4xp75_ASAP7_75t_L g1175 ( 
.A(n_1166),
.B(n_1048),
.C(n_1032),
.D(n_1034),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_SL g1176 ( 
.A(n_1165),
.B(n_1027),
.C(n_952),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_L g1177 ( 
.A(n_1176),
.B(n_952),
.C(n_1015),
.Y(n_1177)
);

INVxp33_ASAP7_75t_SL g1178 ( 
.A(n_1174),
.Y(n_1178)
);

NOR2x1_ASAP7_75t_L g1179 ( 
.A(n_1171),
.B(n_957),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1173),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_L g1181 ( 
.A(n_1172),
.B(n_960),
.C(n_1048),
.Y(n_1181)
);

NAND3x2_ASAP7_75t_L g1182 ( 
.A(n_1170),
.B(n_1064),
.C(n_1033),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_SL g1183 ( 
.A(n_1175),
.B(n_1031),
.Y(n_1183)
);

NAND3x1_ASAP7_75t_SL g1184 ( 
.A(n_1171),
.B(n_1051),
.C(n_1070),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1179),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1180),
.B(n_1075),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1181),
.B(n_990),
.C(n_1031),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1185),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1186),
.Y(n_1189)
);

AOI211xp5_ASAP7_75t_L g1190 ( 
.A1(n_1187),
.A2(n_1177),
.B(n_1183),
.C(n_1178),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1188),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1189),
.Y(n_1192)
);

XNOR2x1_ASAP7_75t_L g1193 ( 
.A(n_1191),
.B(n_1182),
.Y(n_1193)
);

AOI32xp33_ASAP7_75t_L g1194 ( 
.A1(n_1192),
.A2(n_1190),
.A3(n_1184),
.B1(n_960),
.B2(n_1034),
.Y(n_1194)
);

AO22x2_ASAP7_75t_L g1195 ( 
.A1(n_1191),
.A2(n_1032),
.B1(n_1034),
.B2(n_1046),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1193),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1195),
.Y(n_1197)
);

XOR2xp5_ASAP7_75t_L g1198 ( 
.A(n_1194),
.B(n_1001),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1196),
.A2(n_1032),
.B1(n_953),
.B2(n_1009),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1199),
.A2(n_1197),
.B(n_1198),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1200),
.B(n_953),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1201),
.A2(n_1001),
.B1(n_1009),
.B2(n_1005),
.Y(n_1202)
);


endmodule