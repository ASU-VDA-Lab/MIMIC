module fake_netlist_6_2130_n_72 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_10, n_72);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_72;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_18;
wire n_24;
wire n_21;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_17;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_64;
wire n_30;
wire n_43;
wire n_48;
wire n_47;
wire n_19;
wire n_29;
wire n_65;
wire n_31;
wire n_62;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

AND2x4_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_2),
.Y(n_21)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_18),
.B(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_20),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_25),
.B(n_23),
.C(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx2_ASAP7_75t_SL g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_40),
.B1(n_41),
.B2(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_48),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_21),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_30),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_23),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_47),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_50),
.B(n_43),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_43),
.B(n_44),
.C(n_25),
.Y(n_60)
);

NOR3x1_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_54),
.C(n_19),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_56),
.C(n_55),
.Y(n_62)
);

AOI221xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_57),
.B1(n_42),
.B2(n_44),
.C(n_27),
.Y(n_63)
);

OAI211xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_44),
.B(n_17),
.C(n_19),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_50),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_24),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_7),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_69),
.B(n_27),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_10),
.B(n_11),
.Y(n_72)
);


endmodule