module fake_jpeg_2740_n_132 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_43),
.Y(n_61)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_15),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_48),
.B1(n_41),
.B2(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_9),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_16),
.B(n_12),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_30),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_59),
.B1(n_73),
.B2(n_70),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_70),
.Y(n_88)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_89),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_42),
.B1(n_60),
.B2(n_71),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_93),
.Y(n_100)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_63),
.C(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_88),
.B(n_91),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_92),
.B1(n_93),
.B2(n_82),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_99),
.B1(n_101),
.B2(n_100),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_81),
.C(n_80),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.C(n_100),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_82),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_112),
.C(n_113),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_106),
.C(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_123),
.B(n_96),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.B(n_124),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_117),
.B(n_119),
.Y(n_126)
);

AOI311xp33_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_128),
.A3(n_103),
.B(n_111),
.C(n_102),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_118),
.CI(n_114),
.CON(n_128),
.SN(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_97),
.B(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_97),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_79),
.Y(n_132)
);


endmodule