module fake_jpeg_21027_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_29),
.B1(n_31),
.B2(n_30),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_44),
.B1(n_40),
.B2(n_18),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_29),
.B1(n_31),
.B2(n_30),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_37),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_52),
.Y(n_98)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_44),
.B1(n_35),
.B2(n_45),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_84),
.B1(n_23),
.B2(n_58),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_73),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_86),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_39),
.B1(n_41),
.B2(n_40),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_85),
.B1(n_89),
.B2(n_48),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_53),
.B1(n_25),
.B2(n_23),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_58),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_28),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_63),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_94),
.B(n_96),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_101),
.B1(n_67),
.B2(n_81),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_57),
.B1(n_54),
.B2(n_48),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_104),
.B1(n_110),
.B2(n_112),
.Y(n_128)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_42),
.B1(n_38),
.B2(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_25),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_42),
.B1(n_38),
.B2(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_28),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_88),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_43),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_66),
.C(n_91),
.Y(n_139)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_27),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_66),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_32),
.B1(n_21),
.B2(n_34),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_122),
.B1(n_89),
.B2(n_85),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_32),
.B1(n_34),
.B2(n_33),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_123),
.B(n_95),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_68),
.B(n_71),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_133),
.B(n_108),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_71),
.B1(n_86),
.B2(n_83),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_132),
.B1(n_143),
.B2(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_134),
.B1(n_147),
.B2(n_149),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_94),
.B(n_84),
.C(n_68),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_78),
.B1(n_69),
.B2(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_145),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_120),
.C(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_105),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_92),
.B1(n_69),
.B2(n_93),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_92),
.B1(n_82),
.B2(n_76),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_32),
.B1(n_34),
.B2(n_33),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_112),
.B1(n_98),
.B2(n_116),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_95),
.B(n_105),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

AOI22x1_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_117),
.B1(n_98),
.B2(n_104),
.Y(n_152)
);

AOI22x1_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_139),
.B1(n_135),
.B2(n_124),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_156),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_137),
.C(n_150),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_169),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_98),
.B1(n_113),
.B2(n_99),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_172),
.B1(n_176),
.B2(n_134),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_175),
.B(n_152),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_97),
.B1(n_106),
.B2(n_115),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_174),
.B1(n_178),
.B2(n_148),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_106),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_173),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_97),
.B1(n_118),
.B2(n_15),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_97),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_22),
.B(n_19),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_32),
.B1(n_27),
.B2(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_124),
.B(n_28),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_178),
.B1(n_159),
.B2(n_158),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_189),
.C(n_195),
.Y(n_225)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_206),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_150),
.C(n_145),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_125),
.B1(n_14),
.B2(n_2),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_125),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_200),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_79),
.C(n_70),
.Y(n_195)
);

XNOR2x2_ASAP7_75t_SL g219 ( 
.A(n_196),
.B(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_79),
.C(n_70),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_199),
.C(n_209),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_22),
.C(n_19),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_20),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_202),
.A2(n_176),
.B1(n_172),
.B2(n_167),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_20),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_20),
.C(n_4),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_3),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_169),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_185),
.B1(n_153),
.B2(n_160),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_216),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_215),
.A2(n_236),
.B(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_182),
.B1(n_210),
.B2(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_229),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_162),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_160),
.Y(n_237)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_205),
.C(n_184),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_242),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_193),
.B(n_155),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_247),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_243),
.A2(n_212),
.B1(n_232),
.B2(n_214),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_200),
.C(n_199),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_233),
.C(n_225),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_155),
.C(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_209),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_258),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_226),
.B(n_211),
.CI(n_173),
.CON(n_256),
.SN(n_256)
);

XOR2x2_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_3),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_162),
.B(n_5),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_220),
.Y(n_267)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_251),
.C(n_254),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_233),
.C(n_226),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_223),
.C(n_215),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_275),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_213),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_274),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_217),
.C(n_212),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_264),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_271),
.A2(n_252),
.B1(n_257),
.B2(n_248),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_285),
.B1(n_5),
.B2(n_6),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_250),
.B1(n_252),
.B2(n_241),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_269),
.B1(n_262),
.B2(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_255),
.B(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_243),
.B1(n_244),
.B2(n_239),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_246),
.B(n_256),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_299),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_3),
.Y(n_296)
);

OAI221xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_279),
.B1(n_281),
.B2(n_285),
.C(n_282),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_13),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_7),
.C(n_8),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_303),
.C(n_291),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_13),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_9),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_7),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_280),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_7),
.C(n_8),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_310),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_290),
.B(n_10),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_298),
.B(n_301),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_9),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_9),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_308),
.A2(n_293),
.B(n_297),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_316),
.A2(n_307),
.B(n_300),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_312),
.B(n_12),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_306),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_303),
.B(n_307),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_315),
.B1(n_317),
.B2(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_315),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_327),
.C(n_12),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_11),
.B(n_13),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_11),
.Y(n_332)
);


endmodule